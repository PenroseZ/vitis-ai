/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
aB5EHAkrB6NT/NTMoBINikqg8EwKYDaK54FjPax2CptnClXJaFSk1P6Y/9u3FWJjIsff+dSOe3bi
iAx0iPp0pZj8xWoo7D2kuRg+plJgYo3eEH77LyOgJ8X7XStkvgjstpA8MmqOdtjObA2+nWfOXV+w
qbssx3RmnSBBdhARD6rqOFwTf7/3cDuK7QTo3GD8GmkOY+DCob0TXNl7kc1BlYaNbdaJok+U9OEg
YjjGCk5uikHjY6JmbT5Bd71P+OPQhQWHoUBkHUIrhbxZIfDop7LhnylOAsOUmH6p7xY7O9pS50TQ
NpvG9Wsvg8pUSyb0Hyecew+1A6TcJyANzCU7xg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="MxahWTeDMTwz2fyFkxR0OEw6OdcfpBcLNutRaEfsJI4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 816)
`pragma protect data_block
hbfFuBI0Xp74waLCAt9YsPf3nERZBjJfb54Ehp+xys54vuJEGqb3T8TDEJ3ZCjXaS1Cg5lzQVdZS
EDhU0fwqHdgFS26Jn1m6lphap7MMvwhlvzqgRFjXpZcaTDRZKR9IXd/eY+AHWHtTC9r86WZTcjXs
hbsXBt8t0UnRgSe/SLrfp4fkVjan+HocoTVb4J8WEFKxdW5dalibFwU6BpZg3/5YIi950u0gXDB8
uo7lS1qi6R+C+LWiava4RRJvCoT8ucBEVX9Tq1buCti8Sn4vKZSd8sVT/SCdW/EwMG6Dl37Ooj7I
4HElcKv32//HXzS4yN5CT4CjA254aUj23U+xh2T5qbyGdjoCORK/zFHMU55u77SWlaR04t92Jkzk
xACB6OkLCo1ApDykhsCAIyrHDlUibW1TOD41vlNtpYkvHyb7gWWYdHV+qzlWDkWwRocwRDQqaA8H
vzEnvFqxWGwSLACu0BKiPQbMhCioKccNpWYVdmmfJsXPXZelwXO7nIiy3C//kuQ9Ojq0oqZNaFP6
S9tvrjelI1acaly2jxWazjuBU4gMqCFiQkiT5gMs6l5osVxR/w1zQulCUTHhiK48mc7CVzz2Lkby
CmbrhZMm8JqmCJ4niCw6lobXnmcYvmhFL3/8au5H5gBh865SAIAs00thO66a8uA1xVbbx8FXnFo7
dZERMvY+zMDE3q7KJl8DoJhIIv9QhYI3CUivINTO0r5YIaoDYl3xVVbkx3JH6Ik9+/3HxQi8QkeM
ZwrUYF7zUhLwqokI6mXSBjLRxQhHHc6RL8FxQl4oGtSLlX39bz4BUS79uIBv+/YGuqiO/ZkTAdUi
GD6KYaLBnWUlMR+OWUtxHDs+85Qb/6ciWJmUEfzQMe0PlilkAe3G1wd2P+lwKJzSQSBtd9HokvMh
QBQ/lYZnZ0N9z804pEHAIghT4PmrsYzqX20mRGUF57/b3gD/pt2vSgaXaNI1R+ib1LjigPQvpLGj
BVvxiuq/q61KL1gYJycje9Cf7Pyg/iKSSO9Yc3l3dAtVBPvnms1FjjsaKRDOU/yGENE41D8kInvh
Av+IUL2RJxlwhwX2ECb82QCt
`pragma protect end_protected

