/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
aB5EHAkrB6NT/NTMoBINikqg8EwKYDaK54FjPax2CptnClXJaFSk1P6Y/9u3FWJjIsff+dSOe3bi
iAx0iPp0pZj8xWoo7D2kuRg+plJgYo3eEH77LyOgJ8X7XStkvgjstpA8MmqOdtjObA2+nWfOXV+w
qbssx3RmnSBBdhARD6rqOFwTf7/3cDuK7QTo3GD8GmkOY+DCob0TXNl7kc1BlYaNbdaJok+U9OEg
YjjGCk5uikHjY6JmbT5Bd71P+OPQhQWHoUBkHUIrhbxZIfDop7LhnylOAsOUmH6p7xY7O9pS50TQ
NpvG9Wsvg8pUSyb0Hyecew+1A6TcJyANzCU7xg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="MxahWTeDMTwz2fyFkxR0OEw6OdcfpBcLNutRaEfsJI4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2944)
`pragma protect data_block
hbfFuBI0Xp74waLCAt9YsNdA/S3kOfwALoULO4ZwP3AT7V/OmymIQg1C99IeI0py/GDW7aKroOIY
6xJcSalsJuCT0P+fRgokVPl9rlQ+3zk0HqbVhBBQNIBNcRf+lM38nyWka3bXFBZkKn7PAQx7n2Dv
dyeHyRa2BB8xh4rWslRdye9dhQjHKEWIog03Ryoo82wrpsacnm4SnSwoLbxgKctf05RdeDS+hFxP
8PYaLIithUUKYipG6eLon5OgTAtM8AZCkmf12ZLVlJ2kNbsq7SU+uClpMpb/oiI0DtXgvA2sjFrB
nSR8lzzN+IM0Kmm7OtTM2VOHRpYGRg6JLlz5M10Riw051a2Vks4keqdLA4FRIKrGxx6tAHitgFl1
8k2L08S5f7q/LfZxiceZobbqdMLmEIRTpJ5Dop9wNiQ1Cr0dDC0XYKizTmB46sgyCFvKTANMlydA
r+NStKNBhqCX/IZV66v3ZuP8dE6vhHS2sH1g2xRXjYj27ds0Yo5SsTeJ6blrFQSgmHA8pOxckKY6
d5OdLCZ14nCGrZcE4fIVyhRvvyU2tALGRITUhIb57OEhN3iTlvy300t3gbZzV/iFRdBM9PjGw3nT
BK04Sxgf2HrBceYoz1qxmKWQ7T8eU67pLrkrHpy40Kb8OyOuCOzuLWt2Nm9W/G1ppkP0dAlqKXTb
af+GhnGbqlRk5iHP78SDt4Jpl+UuRgSqaeCN5VnLHuHEyGgOIFGVLD9u/cEFk58p5ekLS+RU9sEw
fnHlz0qciOliftfEYTFBOeROy1IDA3gbnEhnrW37f6yF72QXuaecoGqzIjq9rkTPNxIzRgHtZfT3
42WiDSaoRPK9uRoT8ZDcmigh4RBbVFAEp5NDldgUmFePxi9HSS0OS7YtmmIo7SsvS5M4Z7axeXd2
JnRfKbmqplIPoLdBqt40DrM1vjxjDcSl+Y2U2nHAImWvMhxNcdoPE3maalna0h2oatoTS5HCdy3d
OTVEXiMcJ1vsmhhLuBaVrTMpRbqZb1b/tAJ9UiBARV+alsQbKWyBEmUZob3MVtOFo9BFvitjW+hw
NawreY8Eb1Uwi+L/m4+sZQ0p7dRgmzped6pa9T3yO9sJE+lqZf7CjonDYszor9P8ENHQ5ZuTFwos
t6qjUadWYMFQ0gKzNFdSpDL5aBSK5n3LVVLujEtBoI/O2VYc4fbTD2oejS/ksxQkcPPxdEeyBURA
6tNTo9pSUiaAt/szF+WxDHt36+lLn3Ll89MaatHAJ710PgJJIMX6mqsiJbGXU1lvIjaH99hCSIJw
8sGHG6CZuNdnOak5IhoZunZpSxsCvqJt71Y0Ru+nziGc3VWNrQXzvZ2JQ0oMNT7aWdJOZwaggQ5B
tE7XbUvoxCeasUKuwitQ/e2D0Cd4r1n8KWGxmNPZS7FWrwqb98o3jy1qnz0cAvliE3q9Qg2gQATy
tCyjtrVjiPjwvRYB7ItWk0B1zldAt+4mgHjzAdKcKEWezH/9STM31Hb0+UX4JNXlvcZEf8QtR/4E
kzZJYScMFdF3ribuioFt4NkdQY0gRFLXFGu3Mo5uGidiB7/i093e++3SnTff/51p09TKOEWBtq41
8kJrQaDNDIwBAaCX7ZK/iLuWQgrFcQew/VQAAYBbS/lMKifyEPdKoY4IvNM+lpimvUZCeCVkdtQ2
7pywqF+lDwT0kNTN/Wo0bLY4/ETDnYS5M1sjpAKS6+A+zuvw8quTZYUS24A6pt7xocCrbzmeODxA
4fi0od+Xnzfl4Avlh8rxK02TTZS0DKeIMrTbgRE3HWVU4AM3vLVRK8O5xIbrvJZYwEDynKrNQILH
ODLhJ/4FdjqmzpA+ERBkI0vBEUSmg+WidG/bVfgfbJTbCVkkVlYIu2TM4EfCAB5sn9SA1gpjNGaD
g0ym5YGWl4GOTHyNp691aPkCCHop8Prl3aOx50CLq/b7TFTi3vxHcPXHUX5B+lhvVkj/MPMOibA3
HSC9ogKmyrV4LzmCjZLnMYQm6azq1yQyptrBzS0oPBG1HPWzQs+b0WFNL2So6wm+dvJbrQAqn9aU
MKGvfPZmKgXlgBn3YboDTQrEKxvC8kueUAcLy2X01f5wQ/FkDaH7Xat6dTx27TBuXqejG9n/lGBO
vedujzGIOGaNdI8cIfR4nlo7G0ShGqce+d9Z3Z/mYUzrV5WknPsdF2GpfhTYkNAyRFuSeLIlmSp/
E9uI4Vc9F0onr2fmy4rA+jReiDVUHRcAfqy5b2vm0X/cz74JaA7IVaFep5VTFs/Vg54onbqoF4CB
0SSu8uIfkdL+c6MLgr1urAQKOp2aedl+SyWGK2B3hglQZrZ5Jddc0/Ng3pdazLQ9KJChPosW5cO5
6viKQ563vepQ1dMFCHbQQf+gN+OAks9NYUzl2AIIErg2yEw/okP/5e9Ms9myBfwSa4aU5uQ16u1a
bX8zXgDvm2akcll3DS1+l/zs/M6NP+MiOU6wYQs8YwrUwHSR5abdTM4sBA6g1eV2WDrDt1hhur3d
3ixEvEK4WkMVcliQG/irCFjJVX8+gATFqWvriJdKIAm6ZA8ZBm4hLP3tWpTnJ9Lmw8/Jl3IGVyHU
Kc3ssfjeFceh6xg+cfU8XMvByMuQ2/q1VlCpPU92ajnHbOheX8u6ZS+pobFXYnHA3K72BaGbSjrs
u/jwDSgK8RXwAAEdHJ8GQXqHJ2bgUIlgD8ZtQDqxnDYztk+9SGk4o5+cXkdir1EzClVMjf3DKk++
P33wjCP0/Xl7FIhXd+p7iwKwn6p5iyzlHz5MeB9yB6fvETmrdgQvHgSNuwW0HTiSemeEpugivVBb
q18hO1bgnOOZNjy0gNd8lzkXtfKuXDz8H1d3x94sdFuXueI4WTFjXKIWuEoxLHcrw7YfHrehnSxM
vcMwcrUoS+67h1Joe1rL/VA5Bx/jtZAoY+nsCHRZYSprHb2GrcQ48NfOfU2sybwksXsgDRCxAwcA
XT3kn5+4OX7KuuvdYnNAEtad6XuwNqqzi9xgfWTG41FLYs0yEzsNvwMDX6CkNvAtgIXzxKLWV9U5
NAehh55A8zLABycoFl7ctEiLbA4rCVt9lnKu+9clfoKVoDMrnuvju39OoQUm0dlm9AlFf03miLCf
WjpNu/ZC/rhRUg6BPesfikbtX4l20408fT0khBRu75cx09nlx3JUj90nS21aAGWs78rPfgZTQWkF
ZQBD6pk86tGHRSUECt9WV3E7/fMdDEIYopjqTNAC083sf7GJMe6IruG9FSPBaBNqTxaarFN74wyu
INU3KPjeZDHSTvNodNvue9rh5FwH08M3XrG0E7tg8qzEKdSKuZ7TREBdAxWXdVJDDqL4T4uuImcD
kPXyylP5yclnfu3IocEmZAoluXrg/J//4Mr5goAl+w83S1vPwbnyhNhHP8W5kHMFXY1ru3tYAPKX
Ire67N/pH5jfilnx+TV1CK1FpoZjQq1Eacunav4LuOKdaqBIQhGHRiYwMbSkNQfoBviBcY+Q8349
Q5/w4HePfwDpoNfUYGftha6NZ2VDGoCqRxB2SRTaO6vgRQXSN8Tz3vzCu75O6bFaT6s0+aVOTHLT
Xc7v6QFJlj6fI0hffy006SwkiZWWjjQKvm4lZOxtv3HZthUolWN5B6rsfhq5CSoVXdEC4ASXRuyR
xPVg+PjcAsYW30EUEZg5Gsn3rk5bqnRp9tpW++kW70y4HPruNv4X0ZTbaXaMytDmDNw0vTo2FSzB
qLY1PcuQd8jzdb0ZdRxHB/NNHfG3fmUFur+g9wmiXQQwXg4QIx76kgNIMWnLi4hmqyYJKIRO4HOL
2LgiMmFcvZJkXWegS2/oRgj9/auej9UCXJRobfhXCHnrSu3wDBoOiSWQLAuLXACkc+ij3H/b2Yqt
CzXLH+2gP65aH2YcSdJqryZngqjRVha2jrhVcixAKWDjGi0ZJw==
`pragma protect end_protected

