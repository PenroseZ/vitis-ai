/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
aB5EHAkrB6NT/NTMoBINikqg8EwKYDaK54FjPax2CptnClXJaFSk1P6Y/9u3FWJjIsff+dSOe3bi
iAx0iPp0pZj8xWoo7D2kuRg+plJgYo3eEH77LyOgJ8X7XStkvgjstpA8MmqOdtjObA2+nWfOXV+w
qbssx3RmnSBBdhARD6rqOFwTf7/3cDuK7QTo3GD8GmkOY+DCob0TXNl7kc1BlYaNbdaJok+U9OEg
YjjGCk5uikHjY6JmbT5Bd71P+OPQhQWHoUBkHUIrhbxZIfDop7LhnylOAsOUmH6p7xY7O9pS50TQ
NpvG9Wsvg8pUSyb0Hyecew+1A6TcJyANzCU7xg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="MxahWTeDMTwz2fyFkxR0OEw6OdcfpBcLNutRaEfsJI4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 992)
`pragma protect data_block
hbfFuBI0Xp74waLCAt9YsL6W9TzzqoCCYhCVj0l3sInszhvzPi/e1dgpDs9c9O7szLYHfN+1Z6fZ
U2YwKJptzcH8DkbiHOdcg8Wfp//D7YG8gQJMGfcCaeO6oFbHUC9Pv036OqbLWpaV76oqQw1k+Yzb
aExdWG+PrjAwl6+zkfEksCK7MZxXEoiVUupDE+BKF6OtOcUjATpvZnk2M+F7KsTx8yFqXXok+6oD
2RD31Q141pf7kQlL43uyHszWwjcHEBZ+hfLc6N961u2Fiyu2K54ABn7GK3NEQaGCzI7DB4U3309C
uRfCjiBTT2dimYCWv/kV5XFtkYtjiL/Q0Ph6vZtxJgi3xLDkfXM11gYxXp+0JXi9JDlRcgHl4r1W
qViYMqlwCD9s0zieZBih1QRDWj4maimIwQJ8I8KOG2lPhrbgJQEYoGf7vSI9hOMOEA9mOpLtLu72
9gBc4Bld1/dCzKmf5qGAmrsYJH1JVXyzhrEaMPFUf5oNbHBVO4he09+vWp7Z+Sfm9FjHHL7wtwYN
9//nz743g9sA+vZn1USeazMjBLtO7M9bx7pUmcIi0P/1SUox074AvOeAnDDHNXfmdiQK8hrt7pe+
9OhalTQY/Qze3BClL+GQaoSe5KErxzQMxuPw//tadrrIXXB0zMN+9aE3mnyFOVdOqvDvyZneI4xj
Qw+ZK+ospwBq5RRxYAhadqaHfoK6+k+ZNdnv+fXc5bXeQ09vJRChVIYZpMdukOWtBgfQjHm/079A
P5qasV7Gm8freA/O1qsk8kZgUwt7y2WymLA7un89QD8Ifd+IVStHsdJ9Z4lLZ6HxY95ZNHeLqKdW
RYAgg1q4g86sa5UWU8BInGSRudUNisnEOqK2v2hz6OzVIBR4z1YCu+AqkEJNqIvC6jIC492Bj0QR
QH2HVoJ154QkkNRjRxpb+PbSs1fmb5+cnBlC7m5sgIOfYB7cgcGDZ79UMlczOoA6OzlIcjYNUeEd
9Feb/Tc9IpB/pMj4RjqoBg8y5uj2qYoHC/p2xd5ZtfbyTlvkZYnJ5Eg9UmILhV+eBj4UQRbHXWWB
DpN/y4nwYcc1qh+MUmeuzDrY3qbR4EyfX9BsBDjfPKp+PCOrnrWCmKR31gFsqZYK2X+mpOEIWTOY
deLZsNhrRWxFsflEt8fjpk5FE5GI18lVzohs49vX7xe/xKuxUE+PL6kTVqFy5fwYWRA+XGFjd6nR
A2UXxMtWJC4I1fhOZMIpzzssqmezK/Q/t832hVqpb1Gu65mbgbnjMvfnS4VfKcI3JrwJLaCMvUPM
k5p/rUvCZ71smuYJ2qKTn6/B1rxoWY8=
`pragma protect end_protected

