/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
aB5EHAkrB6NT/NTMoBINikqg8EwKYDaK54FjPax2CptnClXJaFSk1P6Y/9u3FWJjIsff+dSOe3bi
iAx0iPp0pZj8xWoo7D2kuRg+plJgYo3eEH77LyOgJ8X7XStkvgjstpA8MmqOdtjObA2+nWfOXV+w
qbssx3RmnSBBdhARD6rqOFwTf7/3cDuK7QTo3GD8GmkOY+DCob0TXNl7kc1BlYaNbdaJok+U9OEg
YjjGCk5uikHjY6JmbT5Bd71P+OPQhQWHoUBkHUIrhbxZIfDop7LhnylOAsOUmH6p7xY7O9pS50TQ
NpvG9Wsvg8pUSyb0Hyecew+1A6TcJyANzCU7xg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="MxahWTeDMTwz2fyFkxR0OEw6OdcfpBcLNutRaEfsJI4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56960)
`pragma protect data_block
hbfFuBI0Xp74waLCAt9YsGebtb27RHl0kutnm4sG/ZLLvdv/HQsfRJA16IablFZqkMOyh7LeWFal
PfULlo3GDfxegAAVLGbOzJ/XbIumvLfsfSWOvKyRkob4G+ukRtdFKJgzVXym2S9kxDVbLYmLIpdO
tGm5nq2wnKDBfb/yPOrp9l8uYU6zERHy4M5RVhayxbcaagj/LVN5ldnemc6X6hKUWVLFM049Eobd
vusT51tWDDEJWpUH8WuzR6KVA+fOPX7/aNTCQB1d8UF/Qf3ArCGp8neajyDjKlxFrqTWwgcewAu1
fmismWg+/w4a7QmSfrOWBY7d3ThXQQYdOXAzfKmmqoBGHZ6H1fo5dBLyQU1e4U5badAx11c6i8M2
ryVoc/3LfPCO/lF6ad+gAl7hhT3pladvGHairYVdTQAULyANfRhQ+Yu8qgAxYFBDKUcE7GWbnM/u
4V3G75r1nB9lT0zNlwJoJ+WbKRLdF8Q3jUaNDYfZDVoI0zvd74XdRl9kFqXYU3FsTpLcmsjgwLMV
7gbQ4JwLx1DslOGijga/TxUZ1cvX+66lE6ruyvnQAHluC4AANomP8oSliw0NNcwKwP8dAPuIdOeK
KUbmqU/+u8yJEDxYIAgTnTBdJf6wxMO5BjYF0ibIDZFYV5TzOsQYV6ouJWaiCpQBBrckH7rsuPeW
ZxjTq9XWtq3KA9IHNGcwGhhiHafKQueBvc5Cvw42eskMXmTpN9Tz88vTeyF/bGVvwFrTDP3knviF
NVJ3VSJEsFaZdX85e6QKE8xasQM3wqwzoAJnp8kWJSHsixwB3aXMpqZNL7OH2tzndl12PyZ8THdc
2Po+g+oeMKeW7/x+N/wyHniGQAmz2Q37RYE1M5YeT4hyrceAhF4l/GWVjkMyG3qMh/8Vci7wGijg
UITwvTStACKlFtnpS77hIucn6blNcvKs2uGADuylFrJ1gVVP7ECMZM6f0UMWXkfeOG8Krbi3WNbQ
uIiJXh1nQVi825eR8RSpsUW35ZCDB1zix3Kblq9Jy7sJihRIWt9nRjidVrRR+aJQbAdUsEXqZHdV
L/EFiD4axII+dXOkHX0tgrSMRyEkyEUvKo9ahJmxPCW3m95jsgcFwdfxVBu7AeSCnuXnLiC5h2xU
ZVjuN5Fv0jgnVpwZCT09XaS3l3323WYcGEZ3+UcZzaw551FIYX+Zjn3/rh6mqVJ2gJEZrcr5vOTV
2oDS3ev2WH66ORCcYSIelNygnc/8srZnUPnDh8pOHsj6PEE7Dw+piYUfpxzETADWgybHn0aksa4r
yDb22RvoRVhFwBCflX5g/T9CEyzF+d56f80/8jXHBg8d9s0hzkqUiFzGZWPBaH+BpXC9OhDB4VKv
Q+WYSnBAF5PNCx7DcP93TlO1x91FPD+5t1iTN8CnUVaA1opb/D1yLWuZ4VA3DGW5DLs2Sij5e99u
6vSuiQgfjGabFgcKVt9WohvyOpr79hB3c1R5NpIJzKpCu3AAXyZRk6oTJpZ947PnGP5yXQaNfk/U
uQDEaNTZ/fJQ4N0KqVnSblq4hlhc9Nv4L53plfKf1vcovhMQWRvRB3HuPPzk0gle3A8Z2vgIuqvG
m+5btNbdBy6Z6iR/t0FgUwbKopDBqphL/dMTS7OmqCRo8eGTqddG7g7LCm+7G6Uko5J+Isempd8w
eg/H363dRNHpeIEC7pz4gv41lDpLVGGfNYA5aImpcTjEhjj+raQ7LTRb64uPoCgAR7nrAMw28m1T
WwesH+PMO0QvZbjfl98aa6x4+Jf5XtL2ecLtDzkgQ9YCmYsBkiPjMiRm5rq1Qy6ntDd1VkUkTVO+
GdW8XmJWg+lwOu66W51RmwwC1QdJLdMNI+YGV8XGQghGBeG+RtM/ZFWAQpQVd6rEsSk+A5c3aVWq
09INvc7VEEhpCQImHGSVCrDHGPXlN4OadS1HcM0N/CDJxW2obYthFJjr9t2fx9ENz7Hdwh/3Em4k
Vns+FNaw7wkyo383D0wiB7fNhnHXNbJpIvSO2/Nnyw2dMJqx2zlioPEngKT9s1JW79BuISfVnHRe
3ZdufPUPnhDUJ6dbFQaKTjw8yWS6UoitNA77MF3LVjpFqRat7N2r2FgSU0RweOtgKVSshSyn8aDy
g8ne0x8FBmbWmRVPnZqBzj5pAeTaK+xJk6Zj2OtqwCr9Tqp1AgQr84krd11YQS6Z901V5xKITo3V
FJwat37o7mo/qDemrsjNr07Yq7oMk2s8c+pcUi1J1s+DS44MlidqKneExGljoChlyD9BqcD70wHi
NFjzUqaqs7KpOLiGPB+RQmCfvGMuqFmPwltWEh5wU3q7G6BxLLWXR+Ygx/0YcTO4xDsaG0FRp94E
LO8z/YZHe1VZik5cQzxllywtOfb4VMHWtJjf0vFn54pVhFJ3PufWg6r4KkLxodzRfPsTHBGNgxQy
katGzNKWn1Rpmg1NRosj8pDaBWF3eUGdx7MOmbPsE/zvxqFlBk8bkZWma/bS7Byyr23gX1VJKndu
j2G/wiWvK3GouS220eIJiwSdDP2PUDe8s11+afmyp0UGf++e0WjUKrZhCx10CH9/47hx0HFX/e7l
TToEuN69mZ1ofbIPxwi3U+JbF3NIVWU5dWXW8RcI0NQZKGgX9VFk1T6o5lSujxYlnuU5o+nYDnSZ
qQ36thXGuuVo2e2pr3KS522p6o0N/tei9/y0O4ui+HguYuibFTpOtEDUPeKt709BYWC/uNkrRoV8
W+dvEM5c+cxdobjGTR3e2wDGs3y6ivlfzO4BlVTtsWj98ioUG/VarQm1kR29brXgN1GBwCjedlEz
qiR8ihlEUs2RWjRMG73mC1sc6JfZ6LTp6BQEs+PuaH28IM/+iQ2TpDFm9DYRwfQjsY472wrJOwWj
miolN/13vGy/JLrLx1woLESytksm80S8y5tbROeJKmEXNtcsZh25+emOU3mFoABzwOOkQrcS1Xug
W0E9RRLhPC6TxsIXzT4QMuvHXAOqbgriNWLgEZXZGsn0IuI56SHI5qVs0J0Enaq+0FLMQHDn31wJ
bNZzRWAeTcS2/O3n6CzbLkACmEjS83xGYp/4pG21R6L6wWaQSR2lMGdcYsN7zycWOKbPCv6z5Gq1
Eq7faTZ05czkkYYJ9Lsb6Ft5y2ypuMMg70I8fiIADscUxE3q4Spds1yGaWC51vOEmJnYNV13G8ID
63YssCkUFzieIhN70d7bbatpj8KtuEgkuVdGcwcySL+xh8TuSq6+gI8bF39+PlzpyCuhZRjjLPrB
sKHejzkJHflXMOjCQlcwwnGIyOFJXWmXPRpQoynuzBiDexVSelB9n1u9s6kyI+5hqa1YTaseIBvO
QX71o6B1mwrE6T71hGrLT3kfDHT/5fVaFjylmt6UGiR4WT/NsUkJXvldSbUQKKxV2sYMRBflA1/R
6JEpqIuR1H1CmtF4Yjbw9wvYxqKT7UK4ZtHPRWt6cTWmEfhhVrBaegjy0MojlaVXvHkGSHwsRg+l
kQCeUmyeVujvjxuTxnvQ5xkQ1xp85S9d6B9OuxdC6F+tVo/EovSxpyhlCSiwl7hO4NvcgT40xgnU
AivnHWJe18E+kQ8BpzO/mCCNjZSVRmvqgrTVyskXwr1htyNZOxfLzJbMGnvbfD3+qIsd6KklOHzy
/Vqptxy3mrmY+pRno0HTDeIvpo8hjXxpZjF9iIDtjOEibWFKGLJ25Z1E7ngDHoMFdlCw/101m0yP
eXbgfn/9124KBpIe3g90nnzQgmALHvLt+VXF8wXFPFqvc8zwDc8gW1JqOvYZC/LHBYaJLvtIS8nV
Og20nX56rZbNzjDxaitiOYQClqn9PlTbOptiuNLJSPMTch6sIZkhkaTudoWZrMFLgzvCTzfE74QY
Lp1h9a0Fx5Pl0RNbS/neGYfHGmStBl+JZvf8afhpEI862341yM8AYyJ/9E36ueCi8j5mV1r4n/BX
cxU3ze3dj0vJyUJyT7Z9FdSoFg9k7cZUkqedkQYCK3J5a9YcbT2i583nkoqI9Orh341K2TCr6Kpc
EyIz7fJhJTx57tyT/w3A7niUva6EJjU1lBvGC2u2tR38Y+irG/R3+VVG3uDspy3+lTg17tyEdfgg
QjGEolmT5/HLSzcOVzLKZAFBvLPh0f88dUoFh/jpPQeq/kg4WsvQPjt+081JdIdECPZbEIOm7wRg
ntMJBUIRLtnDKfv0+HueErLZBKp+UzDsONL5Juaa1z5BivxFJiCjgD+0hftUrwE1ah8PLYsCBgRI
Hk5CZmYmP+m0nIVXkYsSjkHEpeCc8dv/6BV7OKpVl2lIm0qqnFtKNbiqL91MS4Yw1AF6nXeb8EL7
4C2qBIBlZ/F0PLaIpp0RqegXhfbTOkLVOU0WNzTavhZGVi1qNcBQxcueE2Xy3sVezMqPP0V/KLkY
AS1uQvwUkvzQZgxRyP25qkIoWH/hMyn1o1pKnhmp/PTvl4HBB8MmMoS18XvZUQkgLqFvPPHPnuxy
Vv3mi1rtkcNoFOWJrVfX/reoSCkJU0etZ5dRn62iESZU9Jh9jUJc9tRx066VEOJVYZj9o0a6MODq
q/YXnueygbXkcE51Dd6Yy1rqXqQ93jYzLkNR6Vr0YgkLCu9csElbWvhOsxBCLV/NyXh71vreGpyD
km7ePlbJKNoZlnONj5SlX15Kf63yKRopAbujeEZjYa8Nfv5VAEBqxz1VhH8rjpkAav1YmV+b/FSS
G1EpXFsJ9/wATlpWqRisrZ+RQ9z9mTxlpYMZv+LZvuMZ1ymZlFQinRYECT6zdrNWPjuU0amemLBN
jP2Z40KZRTwm/Hl0YdM5lB7eWxsP7swA3swTFY7yG+Xpu/yqkgMMU+UEbHroOayJYLsn9IWR9C0t
r6sGdxrwEwGEQBHNeQnFwcOXao5MQneziiZbBKsArE0/eALGfQ6CR2903UXp7tN6Eui8ykuJxu5b
SzXrOw9Fkm1EXXdIMRoFe5YZO3Cux0SQOayuwc0utj2d4TjsOVAmAeV1YKNju70fR9DfcZWFitso
lOhZRp4cJQYwar/kKpvHi8AZQRwjnYMFgLv42J+pOXZO8wC1C8aTVJNK//5PLDYdl0BUU5GRzTQx
xko+BCfkx/uvF0nP0JrN/sHjqlN5WWfbuvTW0eX0/++eS9mS4IdmcIGKR8fmgaHBLU0EQBgpNppu
hFr/5GyIAV8FjXEUKWHLmMnhOPTxIJbPfLoepEjH8b4dX28enEaPEeaJ+mGBGnGUg2pmJO3WhTvz
EQorJcyRrf5IbXGeFoskBn3pYJFPpsEcBt/UfRNdc7PxQozpskzw3hfHb8itxjpbwFnNthSZiMe7
I1RC8gF3tJ0X9l5sjDHrB8uUvTHK3FQavk5W6ThrSoL9TqGtfEvj0ufNyoQJjGRzSnyuRxVH53tg
3ANbbskWSpsrzEHkDhNuVIeaEvyzJzC7+brsyK/rUQSvqmEmvEyIW7j95lvNVgHi4XRrn22Wavvo
XZQjmPXq4IME07iY8X74mrtGuvIDuPEx//oFbvnnB2ibko47kUT38P4c/e3W/awj0JMgE844q7iZ
hReOPmXvMKVEuhwhSTH3xBB2NPb2JFOB5cznSfo/WCAByfL8UzbMVJBzqTwss1t/A/M93ickm9Lu
jG3WtrSNFTYZFepw9Q23t+FTIr0Jmon9rdB4k26s5reYvuzBY2HRAXrmfFMhhsPGIcqaWFlBCOyY
VndKONrYnTr182rTX8sb4KzDtHL9beCOZUTjDT+/poWtb1mzxs4vgcCYxsb0iwGLOo1rNRgAe8xb
iPWv0F39EQvcccI52eoqTXSzk7jrZ7pAdiGVziS+BnXc41WB41FskyDWLAZp9Fdq1vyja8ycxZDT
mH3bGprg0LvobmNyi5aRvEvXZ4O27IbNQZvfW0arQqxTiJK6VpZ2sd9dy9HSr+4cK3pcUjpQkhIJ
g8dfIjT9EInm5m2DgcFOPoVTJ93s/te+cuW4dIH3Ql3Ux9e3UDYVen7kDvf5AVrglde8lgT1LXJ5
/c5kW6/vvrNDxO/z7hFcAXwXTJ/tVgsU0gb7AfwTKf3EJkf6zQYLPsj5yM7OebvsRkuuejf/yU4z
2ZCLeNxOtj2djlEh4A1gMrpPDat6Psv5ZVkBzyh21iR/7DNezXXyCeDWfMwMzPEXC2cgfVy+EL9s
GqK/Gpt+gjVSkeSfW549cBz8fOEp6Gzy6qhgdbZ0FE+NE5P6v6PpYNtWjfk4x/1WU6HVu10STiNk
x0XnLV0DfqNjXHcw14AD30Ig/7eJdJllZDSNJfTmPne0c78kdJ2JK0NAB7RESGgqyhB5iCRuPYt/
r3AfZUequgg3neis1djSyiWUv+OMegMm4d/ikJNHnDJEBiVht9bAMCkpWLA4FksUp3X11/HnPO3R
3/dehvPAQF47eK0Qw5DoWmrVnpSm5oQWBaG3MpWqud7hOJJ3NqR6Yk4hVUFsxrybaiOHCJrwzPer
6ytUW+c7rOIzxLLOBtdepeRjYpog/6KydXjvclZFm8k9JwuQYKlKoh+n4ZJsntcs2dCYcLvjuZor
83q1NkVkuFc8Yzk7y5itMo98MXxOJpDdAvNL6VkOIggTixb8Dd4ZmUDGzVAQelfSHV3Co/ksGW/e
eN1njcN07c8QwQfS1glMQsYhqsoMFZNIj8c/E9sd3Ned83nqFpPCBA0E3+ARzHbcspWdXJ16ZfV6
rjLB2wIjJmFRTfGi7elgtpIWpcc922UhvK2tyVAgz3gPFdf9DjjZzwzCNUrzScGRv+/SJzxk5ndE
nLEkBzslGZZzrZDQK/dTGc28VE46x6CY+WY0Hs6UkOk9fRnn/RyLeIHGfioUqmSQPm8c0nxAjrfS
Ncp864HCur4z554slFCv0d7fsKSu/vedaORoT1zi6o9VB/rxqmQ5t9Om8PIUBn527ceIuSZOmakY
uMZBDEe+NNoi1uYQP+i5f1ekqdNWRNzOKuShytpNX8Tt2LveKU5D7wfkmaITdLlzw8zngg+Lp0H0
6ZUDHMm0Jz7ezN/9tn2+7qZOK4PWuKF5LjuOpj/3Bpea1KBx71ckIh8GI8h9/lbQIRKNVmSGQCyv
3VfRgHInbZjC9FPi4085sVTip69Lvg+89N5I1ODnzmSTWyskTqo6T6fQkGtSDRuQ6IKlOF8jtMx9
tKDt5sjVLl5KnBAiRP5gRwihBaJRjc0o8ybzQ9av+XZE2x35QoCMWtsWtOwEJE6rTbrLPVendZNY
TaPgHjjQ/UFL4ZLUM0oYhMLQmQ3cOlnx47sT5ul/wVQujL2UO3AuYaCHLyS86dRR7eQVx21dUAB0
5Z0eXigcVMKI9gyjhvKzRjELVTdWqBXRYEOBY8UH+EcVUd4Ex0OcUqWNQbvVoC9GpLBaWfht0icA
k+4FPNZ57fLuQeV6K3xcDT0vkfl9D+bYdSDPIwqG8ZBOOacwqjGErk63a5EmuSJtvHNvfFtgxb2x
6LGN3y8QSDE0b6HRlkKTRuRoCVm1DQ/UdKijMaBC76pypy4KCBk/booxsz+y/P4NLp7kMeuI1/kh
P9mhAinedFeZixHyxmRAY7Ue46z6nclAHkZs/AtJ+xuD952TbTBdYUsP4Cdf8tRZyGWjLt9iEuxv
8TeYufl+KpjNQHFf4UbmMDr8XL+smOgds601CHfKiVcb2G+lpN4wkXEv50fmu57273nr8ryj+YjA
q+OwT8OXljGNIoRBpZvO9K0UCzUYsLeaNN6Vh1p8G9j2KhUIefV+gUYlzF7BuJZA4QJ29X+JF9y2
gEt/thtCp/dmA6JmX+Nc8C+WPPekdgFPSOHuAiGEqSBodoSDguVO2VEm1rUOlukZ9rTBl4fVlC7h
U6nwaasY6/wqRdsWDfO+ad9P6tSJ3HBlpXbfELKBvmaxvBneALmoVyISU7zIxYITAPBAEnSH9k8N
qkv8QQY8qU15rRq5PbdHB1CbVa5uRMon74tLz+x7bZRW+mvyzG4qg25azlZcz6DYtmK+FWqYeeIg
Mnl0QYx0Z9InkKd+L0VLDuOMxvGO4gGpHUM5L3iD8f/shIOf+eiF7aHSib4lg9QHbLF7akTJpM8w
eZF6CXhH6ikmeKoLoBCf2AwvL7Quir3ytx0xi29GEILO8LjZwijg6206zGCQ7t/TiwsfY6ZzZ3eo
Qhlq2mvmPqhkh3r10GZX9X8u1P5CbREsGY3H67AQFgG0ulKuoSGilstyoA8RHb7Hg6ecOhnDDfYn
RJMGdsIz7c+97ciy7AL17JJyHDqEsvG9CFElY4K51AXRc4erP1qPuc8LCddK2wtLzc+YIkibjhyU
tVRNe70e5aNB5xuj1ZpeYCCP7M14GBvwPll8wYKQTaqekfT9STwZJh3MjAZZFfUyG5IUbxGoK9J/
3nD+YGWR+Y/di8v2tOx99Yt5TQo+/gGnblTPcu5kp5cr1q5GLerBHZGYYkoMFEKWO4xfr6bwq/U+
tLRbE6lSk8EDsEdJtJJZNggO99gFeXViMYhQrSIwvH4MD5zOGvsv5VaJbFNgXabEwJf6EUBKkPh6
KVe1Hc1AOIxjcOv4W+CopbcxLLlPebp3RHe/UYAvFYHo4abZF7owgv2mUm5q9pqjAHM1b+UchOYI
OjzIUFj0//RRQbRLzv+HZh0Zoh6UpBMkd5RVeH7+6JCLOGdqxkHNtolDvaAZ7Py2g1+B0uxR1L+p
7ReslgyKDi3hACzTY+d2cdKnP0ef7b1M4pXd3DSg8aUyIRtmliXHEw37Wh/8ZXxPDIsUTqTqQlzP
92ARZQOcNRk4cLjZJepBfikis96DQKv2ivOZmnKoQdLVwDIeroNyVAsfvWi9ROAJI+pDpzu5mZxJ
1NN8tBHg0os9IbQo3OuoXpxKJGH/B271MZCQY5SnNOCRCR7gT3ahTYOdn1cZYQXvXuwKj+3XeVvX
vDeW4f1N811BomaxLISrrE+87xh3vPisv7SOhGnb9nDJJrZWsc4KGbp/r/Rfy2+pKe3+cZLqYx9h
khzK6OKUYcLFYmK4/Lfjw5X4MASa4XrOtzQbqzFLTjZfD771UYG8Qq8/vzsmh2sSsVBTJhijbjng
TDglRRiIVLi9V9GOKOJlYezkrskuCkP/VH8p/yEiuiKXpnReB7lkFIOezhZlZCo10LcOkIH9sJZr
ep40vtKvQOgs6T5ggaeb9tGgttejRPfwiVBEWiyNcl3hXQHMyxALDrkVwjEXt5+Duc3+Mj9tlht6
WikZPgo7/q5EkGEhmYRdgb82CABJMj4p3FunZic0FDVHKJIDzHrV+7nMH/bgXZAaxl87t9D7yEwD
TsFqt25OaQWe5UPZPBKSO6+ts2/tlOk4uNdfSiJFlmUdXUgMvJj0oM342KOdD1WwU3L/dq/ZXn/o
oJxG7AheQIA8ncNTQOMXexsoQaEJ8YODZFmKKqRoC6bQ8Gje2bORJ9QIXQkOf5ZyAMLoBakEugXK
gB8KaZ6ZVTjSXfc1IvGuQrF7SqxNlZ5Y0Gferi1sRL/3hs3v2E81swcY+NasjsO2tiF+bQPHkJoQ
WnfCX7Ot4t2I5uwpo1k88BTG65By2QLIo/cDpRR7nO7G7/1E6HSweVZRxU6cgwN4x2qpPRmHJD6X
WMGYe9/kju4t2k3c4VZVia8pnoG0wcKC4+US0rfbO1sEF53lGnToU7p++yvogzAoUB4+KAaLPpbO
zzGW5QDRBUqOP40cs3t4sBxasj2B5RoFYMrPlRKK1lOMKNURIo3NacaI1w4NsmyN1dKB+xKtq6aF
AD2u/W39y5C47o45/p5aCV95lbkztDzXRE7P6DpVhKuEspNOHd3auLKydVm5k3a2Xr8ELcr1cKDD
8CdPb+XJ6eXz7f6Ri0yQgZqCFRZ9RLN5w+zFnSCyfpREXVBs4HLPexBDihji07E+/TA5PoAjvN2k
KS69HRrOLXU62RNmc+xRvdwyF3GdgRKui+BrFlH2hajKjQTV6fcWKxFESSmtUy1knwiN8Q8PTElG
Alm/75P4aZpdD83lzTy/XsbRsZAXUiBScKd0KV9kvHe88n082reijjw2HdfZ54YdW6O/aQkuxv+Z
7iHpYjdiIDUz4B4Fr+v1hhw4GyJ2GqyIowJRkBW5Y8SM934QQpTsN66Ni4VaZ0ZYIuBBJIgXYq/n
Yl6W0KyopRRV+m0vTJq4N0psoZzDx0VOYyl0KJUuf86aOQt4VYwVUJZxWxbnCnhYUn56IFYG0m58
jQnk1Zlc/GzsXFGzHoxvxagvkXlVzn6vmHuPpmHXIt/DFQu+w2LmSQEdJCiY39lgSCHDkf1WFnwQ
j7U3B4H1ofVwXo+6xBLPSs8cMN3qR/29VGFbUrmZrQ6YXIw5PxA572tUnFbm5F6vO1wstyxNgvFz
4pZZdrAZMeH98z1SNUJsBxUhXlya3FoySIViLPTC9DVQNoB8Ky/3k7Hr6/29S+DglA2m+KpKo0K4
UGUGpKeOklkOqmYzKc1+hFUmYmAbiaMRbRPlqQmTwO1pLyYxPZZ58iHNexInDH9rrkPLz36H1X6R
dLkZgyE7OyY0yM5fiYoB9l6yeR+AH0aydGDaDx2ImJOiTfwOAiTvOAHaJWnrveXy0Jsb2iBmIC/I
zUIj5qRHd81majwImwTf6NILEnNU3L8+V3OHnAZpRDB0b5NhSEi1+4u3qInM+M/USYJc83U0vYcG
wXATIhIvt7BRJkjQuwQmCbauPvEwuvv827GwwS2k0RlGCPg6CVCtHVxA+VRLhOqqK50zA08qUr7O
dhh3FwLXGtVl/eIhAmk0t09eVoofBWLWBCCA9CwPh1llg5X4arbmnRI/Sl86x/QtShEUYutjzxA6
756U+cVG9mPG/DPm/By5FeEffEvbcxubdr9rv9yLHaJ6yJ6+PyxfNVLN/UKNNVu17mzPRLtjqgLZ
C19st/jkozfEYNqbwXwr3EKKqk/8R8cN1oMMJ0w/pasrMnFLx3IlMFVhaS5q1OpuE733RNSqxthM
hkh2M2PBeuYAdbJbpYyzQy5lL6KWhOQ8HVXCliZToVSOg89WMP29efz7Cd0mJEUIao10cosRCQaZ
0ZgVCoh8ePujovVb2f4LkU8Zsdf0meUSDujCUKeG9TVSbp8ms28yLi+1r4eTB8E+Vro/y0p6JgcI
OoI2RvitmVlWbrgljSdLa0BG6iKFGvo1eMUU40ynVEmegf5VMA/pfz6vqWRF3BB4Z/OZ5ZPMrdjb
MtHZzYSRSSSQG4gap7szs+sybFOhjh35DYj6h6XEkH1Ku5Vd/AmUKv2N9BiYOznxIB0Rcl6maBga
sb1A0WEgf+G2kQS6UJTuNWcNtg1Fi+7rhlgKdzYNkoBMhsIiBUrl1GpNZCq1V84L603hhqQI/9HF
jHUa1FcZCb8dCDBF80sR0YlLmEITvESE9j6kAzOuYlOvwTtqDiRaicdQ1sV6U7TgT0sxnMRuWZNW
2rWinK1LZZjIHoRNjDL9TeHsSejjPatIgR20DxMiwkitlPgjpDSpon5jwjFILcMo6obDkafLDlve
Ze1rG0Ikmzy2opb7/Q1Ry6VBcftVUcy/BdL5whsMnGjY662nDCowedNUM4TgRfXX3bXYvOB2VacM
9l5oLGbcL//QTc+EakGKmQKgAdbZV7yg79pS011Ma8bVUlgOAYKK2zqVcsES9mtxrwke4R7bKjOY
5ihU+IppG33G7G+NJTyI5/NSrng9KTqY8BcWHTzVtdoS9Hy4IZyC15UTuNSykTKHuJMCVaLvutnI
Sq5Z4tnhrsKexO+TIEyUBWTOXafZNDg2CwKp3JoWOdC0+ktO9MSaaWGd0Xr/srUKnYCBELMWp+wk
3FnbxHgHisBkX9DtWshL92K8F4q1zXZK0hcH+lSCNvNucScgdOrMieJR995HGGHpbR6l+Cf35Fot
axQdl9KBt+RP8eRtbiJ3hmPq5yk1/LEuhF+bmJmJ7GJXtRqkq5/LtcQHdXVv43sqWT75xNVdiSI3
esm+S1bfpIAKd+T2v077rY+zVlFgRCBXVMYBpQuRrGCTNl+3YsRWHSGXSrH/BTHlWzfr2J0kMr/m
3+GLgRQ7clTd5AGxfi4NaoDS0SFqSxng/UvP2AWAW0xtEHlu9VWp87pdDjsC6cveGAd451IoCO98
Eibtu/A+gX6gPWJL8FIIoD5JEPo8PvQcShp7pEpwrSLr/q4lfBIKvrgne++LuINu34cefFgefql0
xJssFYmeM3mC/dt598wjN6H5QuVeQreLjsMOPJV+Wx/pkQdrBVihpNM5B2KxgHh34Z0YvoYDwgzY
Z9LbpDXa4egLL+cEyAtUXij07zMQGMCd4fbHoPAtVNxKzxMiRVjyphc3NLNqxTPjqcI5mxBPGh95
oEY16d942YcZAtbD5xfD1agK82HUV7SGd7mKFaR1S0mK27OmY5IeQcoXU07NRr6x9sAeIYSD/frs
Km2F7jreDOsZUcTuGBGVLLaKMQkyXoksRmaR99Am/NtCBX9QfFuv0rkQcKm5wPP06OwTxam54j2l
8jt4Kc2nIzdwqSYXK8IFNPCdhi0qeF9ZhB/s3pap6xbcZL/SmJGxJqVmsnk13mtGJcHbi7J2UubL
At+/C36mhnqNuwYDqHPiEjrTpqzmjPAS7iUbeB6TVfLD1fRD2PxV7RtcjxiD+BOZ8fp4/ks8eZyN
5FT6QQSSnCEWS/xdufr6wsdEMIJ6g49OUCfevBe5jpKbvLj43Reub9Edhrx2hSARgbDymH8aerP4
0lSwUIXyOBRZ6z8V7I23BXh3/7w2Yq5D+E2UrHkb35l5WEmsmlJO4Pivw+lchGkhH/AKcw/7p1zK
nt51E+5vq0Ishvo/hq3vpKz9+F/PiPSblljHVuwCl3HS92PEexrd4lUJ3L6RgJDU4OOAdjo9euXd
AqMBEW+Xf7OhOLKq2n1uc+qstl1hUfYQ+ukvkjVL10DhvTumDFg39wmMjO/ghSh4qGyrRVWC2YVG
rZqcS++IkEX4L+WpCGiTVgwFBDFF+1oxFrbhgWeAiaXPMcSWj5FUG+h2/teL2bX7g63+bCcoE23E
R3NhZyXDZNCrDZLZ9YFA0pj6vad8rl+r5dgEDq+YKQKBjKMv1uuwVwRu3X+3sz/yiQ+rIBJsmTAp
39ARTrfqcLxbLVeHzfixv3MPlqwTzrbEppnme1UiiuRgOzavwK3ZsyxEGKjiark0z7p9P5i8nWyI
FcxIQxA5c06J4ZtGJqqMGvs3zSrZoaPNfJi/+V4xI+MWS06YStQD051LX8budz1HiTocSnGibnaT
cg+FwkOEZXNqOO/UO4hVnFXCf3iqyfuGol8YoelLtEy4+K8UeuxJwoW6UvMKMBGgTi5Q1s6Rp2dW
Bm8lpLH6bzyBb7h7SMX2mV8uJbyrFbML9oeO4uPoxCIIpNe38HzEX+4i/BHu4oSKdm3avdTtXJms
AybaXbsEo9Yx2roUlCkGAI3yyz0+X/GtSjCPIubAZ6/RnWNrAoK9Srx2lN4AJSkOhcicSVGakH0G
ZLATdOXAFio2YvGDZjo4Vq+eWwZ3Be2pGbCj5dyCYHoEBkkGN0w9t2Ty6mHNprzwciQJyBybAyBh
367gLXxNc0A9qQljyE71ZjsZ6mwkWBluLZeLGwcRlA2bPPHCg7+uAPT2YbTkZ6etUe+JOBdWCzi0
TRQhftE8uvwTV2ON89O+B6OLP+2/uAenasbOJe3/Xue4Q+Xq/hABpkYdy8Y6r6eYOoFz7WYfh7OZ
TsVbgjTTJiJDcDpRjUF08F4biJqeBPoSfcOWcNcSGrNWBSL+Jn/cjJOW6IygjZAlApIeq0TFJbUI
/MQ58rxsU87dL9WWKKk3HXJUVM8KjnOGdKl5uS6PEKYU5zoyQUFgj3jCdfb0WzwCMtrJxPDqBorN
WL2/mNY0CR7npiX3sRMghbpsTkVJjTiu6vKdHHPxcgB9gwb1nOCEMvGPL5RX8MNoctAzbM9m9lP8
qlShBZnOINpRU7vXZDDyWWJuod1V10pHvoxdyvPE94ElQpTG040sBDrA/sPi/MJ+qru/UQjdcUxY
4lieT1VDD6wVCcKQiVHGA/1J4mo/l1kLXnau1DoxLgzk1YfUy4gK8KczTpmDr5MKbkT+gtUn9ey/
kOeOY3dJRA7BSxS4eEVzlClT2YKNlI5AiedSegTByFIZHjECGEqYEI1MCYRP4ittgSGIJjnH8sRs
+VdryWzjSFRkny74spm5kp+72SvokmMUSycaKlRkLvLf9q0crICvsGJYmsyBSgjGbbI2XW7YHof+
/gvcRHd54ypXJw67EtWc+BLCqwYOMhi6+ZdD2zGaAIkEYeg0tyvB1MwlXa6BIOtGAVp9EMwb25Uh
gceFQISjYyvhnsEedvWFXCyHGmM37lpwgmynyRksJvGHw5+CgDsSxFcshnCRi4yq6vwCKppbvMsP
1H6PLRW9XYxm+jQ3bSNq4nIf7yPWSebu5fBlKuIlezlNdKsbncZSkmu1B+U99PqGCr8tzfPpywpa
tiGTr1uyKxlQQcMaf82SUdBHYVVHS01LlQsYlzbX1vj30t84MDJSUBvPgMxKIRYj8ulIbPApXoa5
R1LEp+LfkJ/Ca5tiZO7WMQ3CKR7Vdtg2IygQpZiJeU3TgTgveNrgHLYD//6O7hWVXm9TACqc8yeQ
6HJA5L4ypSoWTuhtXbKmrDkn1Qzc5Nl3pk+SPxT9CE/Y2wI+bljWu5hILnjywAP1ArKBv8P06nwf
UhllAlgBI4J4mKj/JDo2kjox86oWtAzhwDXjK9yKjkh8u3oOg2DfqxHM+fowPLWyUyhWkTHWSOXR
RcN00zOrtMUFlZiZNC4nNCFfTj/sMvHu8JVFAqz0G9R953SiSxGiCEl9x67eFCSAbRm/QrVuUXGg
YZh4ZwCHYxmDlybliVe1tq3msiJt2Bjk6+KI5DKchQD0ZTJzVPSP2nhSZHMLUxmiS2f0O5egU6kn
Ve9Y7luLtsNykIOFnQSn72qRsMXcI7ICouhY5MTUS3kc97pO2p811ITaojrHam4MjH75uDfNqthg
oTYArmAYMV/fQjDjkz5HZ4erPa4dPdven0XjPNnP9MZki9AbWMHxl2AELRXfAg3ABYHgp2WjA5A0
rwcYNf2LH/BAAi8sBvj0ZlCjor/agHm8nKpIyRBmc3HJJS7eoPg952QmjXiGmzrTMHOF7YdsCIQY
4kN5XFF9bO1n6Fq4TY1hFYI/Xduok+32aWg9vCSlLGUMqtKRg5/4BU0aV4bgZYzRJtS1DJCMB5yU
a0GLNzuxY3xn2o+TJCqFqdbZ9BGGK8F5uD6in2rbIwEEkpQfRQO4DLDLiEOBYTOYUfJENPMjZI3w
bBzU9WCWKjI8vsQBVDG5IBof3+giBNoWjaLEYVhr6BeWmrEXSXihRIVb6KwzRLoL/LutSr1xAmqK
UlvOVp70kwFnGIX/8b8bGbmPFByjlXaitG8y/FuZQYyrDyB2gNyrmZwYG81yybh9wAp++dwvhMVq
vHUksbsTfAFEGUsjXZKzzUFVQQoYXaVZ8WcMHc4bgis1qG8sdNGCVWIwbau2c2WweyRbzx2zXr7O
pIQLhCAiX4sNA7p/uC3R0wcdmstDNIh+V61JA28q5o+LsPmYpm7/soLz6uYjXmEh3SdAlo0vu9Fe
ALQg9X7aGLokxEBfCE3ODPPasFgkzpfrsB/+oUK2GgWt3QZCXX9G+JvY6AZM091jDryVN8HgT8je
6VZKanm/iW4w3aazaIb8xnCBfeO9XvpDFtpZvFEcbYQ7DpjINhKAS9NyninmTUYkDs/1ENQvMWDi
ehGtYoWHKWJ6qpuDAt92sOnkesMBZdiznI5kBJXeLNJ1oCj4cTAsoNNhnz/AsXDH9SZ25DpV6Uow
LC34rxQYTVzI9l8ugpas0x1eE4MOId8eZ+lF1KcvtpZxVO0SbYgAANOegmO46j5nqG+ZSA1/BJNc
xn/UL+gzEFO66KC77PSZqEd1dJ1LmNNgX5zJz1JM81ZF50nrJZsH127z3yqKqfLncX1+O/T/ionp
Lm6vhXrRViUW5uXqT/l/ZgX9sEJpNcMZq8t5L/igu/y35ud7B24MzMKHvEnHtf9lq01K4ZAFAPHl
d/wQM48+ZB0fGER4UuIA9JpYyMfSeV3A9Vn1LCV6PAuKtzTNVly3Cj0opPrlIiF6ggoNe2LOFeWn
6ClNVZfVw3yYUmtQNnV71F8oD66k7B+wUQFvq1HCoC7sbETCsrcuNY+te3lmLPG2Zv4vVy9O33O7
YtMNVUCd0GXzKvfBh2hIZwz5yExD+rG7oj8VNouifAndI2VUd3c2qC+pOfwOOSIa0JJarEYD0dzE
SofulA44ow0ElsGWNm5lMGcIe0UeAScYWo7qLiTa1+yBTwkmxJSr9U3yHl5gMw76s+oE+YZdRpNn
pqmDEdbkhGYeKjQbFwpVRfLS3bQFoYwyNPLZKgb2X5zKRcgANuisWDV7FfvzW4gt091jrTFnMxZO
kVaAP3zpWBOncKUIbxWaN4Yu4dKGQx2rWw6LrqoREAKkBL49glW4qttiei5aM5gpB7uWcIGxvPRg
Wk3mjgEqRPF4A5s8INszwBsvGweAdRd37PTYcLIeJJpdTAoPHUAXyrb6qLgUvXMW5N3Ya31A4NeG
dQN8xVw7DTN/dgU7DUmIH0QEHQ0gxctrMmzxSnt+I9pJdK/NrI1d9ASvDRI7M6sr6h7BRL1H3GBp
/ciAcvLboXI151wk8o4aXIULoR8RVEKZGw9sW4wJAwhumLQIVhvJFe1Wpf9dL+9A02MKWx7xlmNg
i9o97VDL6R0Xv1guGJIKeSopp2KSlEJ0GSmOD2HgtqyPhdwsy6TKhUKLMQZfUHKYnMmAiSuh2wRc
R7w7jN64Krx65o3OXuiiDP0gFgYbK0WLCKzm4LudSMMv2XXf1DdKeRIFwghjLFTBvuA7jPuPlmlb
su6397ESuvPBG6XspAKo74eeNh5fxBOgyyTHLZqiy5flsSFiongwN+6DFjSu7oBEq3+iCRivdqJG
u5sTe124Dtwk0R+vqxCl4O2OVy8MAYwWuy3i8DhB0+1euXAL1jH7Nn3hXa+iv74mwmDNyY0lkQyn
67ypnWgRBedEjvugXAoN+UaB4B1GpFXgyK1Jn/1Uh7DAaw7WT9BqjoCNnKysshwUlU1/MvoLu2Ud
ZXhP+TH16DHFzt+iCgr5XllzkUtdqH72D2l1UdmdLsmiRg+YO5euitUb5Zncd7RDqg98fQzHnAvw
LKu6p0bYgBitupIX4qyEobuQRxs7V/9j3ltVj4JpBN52is89pWHJk/yEzEl1Dk/snyDoIwbc3fsC
Bp9uUpEE9JzdqC5E38HFw5iBZrC2xwgMBNm7ML9+UeiezlDxPTrCLUD4tgekQF8F2bEkAyQkxCDg
GbMJ0JLsFMiiyjPzvy4vQ7xqzwU8gExzerTSqfWhb/m/HXjWUNfMnZlqmYdZEIPZNLARYRjwmCJI
QwX407tq6jW9e7MA+SO7tN6JUNFMC27ZOWw2arP2bkfjDLNAicHq4IpMuYO39YK/gCZtJXLe2Ibm
YM6PcD8C8wcSB7qeb6nYqNhJ7PC8h1WmfBKF6jloWr3pNm4evJW/c4uqvWhDUMeefI8mvc/z3F8A
EhK3RMBPankqHarHhPvBK/vBC1mWpvKKG5Fn17Gr5xQO6ooKEe484Q45x5QzC8k3y0EReDVfjBJJ
9MEp+GN+MNkzNEEXCSbiT7F29kvksZXa43UmiETWwJ0SEGzCSzKsi+BRAG1v6XsPi6cwUJsYFX0I
h29VCptIwevivLaSbhfQliwXcmn5yl2I8wZsGnLx2AJJ2KxDn7iKuuif+Fv4v7qlrm9cxaVO2Z7p
WUZkMhceN4O0Eac7lEKb4slt4NVusj77H0XH7cjVFsx5yWiWJqvWdGk8YW9a7w4w44eDPNAcKzOQ
c+NRceLlnnPpMTLwAUJkXUViqG5JSRyicVJJpNaDB2bGRk6FVMYwFDg6ouHOdcQZXlCLIFf7e1xb
T5hDhqUZE637AMTGdIEc/OvPWcRboHupEDLvgmIciBEtAWtUDA2B5TJb57XSuHYYtdZzeMmuFTnV
qslvBGuRLT76MVMl5v25rhGtyxiu2RWX7RcTSGUnNjAkJrbg80NPg1EppbKqm4yns9j0Qmh5iumf
jVpO9J/f8eZgn7PZvXquidXrdDH6hgpnDc+nfw7VA6vptr6nTagrDGJxklwXsBw/+EMZYOLNc6D8
W9BeWgE7c1NfqraRDeZt/D/asdkLU7V9LNqZZX0tBaOXz1dhY4aRufYfO2k9TsT5U4Cm808gYtVa
nKSA8fEWdc7FQCMCiCCJh1bpC1orJKrF1RKb1yAh6M59eKVYBkeYYksFAdSOD0WUUKYhxxvKrS2v
UE7lzs66n8TXTt7bmu4e0hxKc8qnDE0CF8s8ywaZMb4hE/5iUBHF6AELcrog2kPsiX8DZyqvpFNf
3Eaum7ciulDUHLyXRhZiIHu4ohL31J3hBmlGxx18PfmtvtU43Jer2jQdzdWhcDkg3mLY9F47KkmJ
97VM3GV+i3KCC10LEG9niHRxCJFMhNTYzrMghrQcPA98voB3OLxQuESJzHsXMiDiM0+qJbBYRcZs
6aKDACervM5XoQBRlaGoc5R8veV93o8jRPc9pamY6DmF8RJ6svBq3ZTnvedIPyqCZ3odlN1cZV15
Sg81OdAHug8PqEtTmeSCvWxVEx6vETVE4DqRCsa5K4XqSuoPjJ2pOKo+Qy77lP3q7saN1nXh4ovW
G0uohAT/bTpoxMyAoZWHf6xSleRtplX5iGbAhGSgMkcm0BcZa/rhrJd04aF6lEL3I0sO1ZKQsrQm
WfOCnijozCMKTM7BGFRYPpTsMwTc5uuJFTJik/DzuNIIti0ag2WAADpQ6/4RcSXgwnV+2eEzwtNI
LSTgrB2gSJaSoHPZgqJCQL6so8yibThssJQQqd/2G3AiAA4163UPUh1DCaReYegKC0FAYEWFGQkw
8g/x5jaccUGcoNTHzSoUdb0+jHTCKRpb8jOAJ3M9VhH0PWXjmEOuocYW6eRuIYL4OlMTGsfRRZm8
6Wn5yVkKj/zD6l5NcP9Ifw24NZi/Wf31AoQdYMPrJkd6fXaQPIDtIzys86t69MrStE+Zj9r+xUPy
p83HhHuqWJz4zE8WRmh6sNupFiIakrXlEKTuOy79trv54i1sPYBTHJ+IteymsH2jsKiRrK/NZLmn
miJin0EIK98qj+B8p8IW/qqX6akjQlO0vt4JY4ONKf0E2UCz5455eBbs0DWVi8sjLYvk2ZRt4/pW
3lR45wv459II4uV6/Tqm8vhLscAI/+Ezr89MmQGT19lpLzYIgBsm6UFRq9T9/nGOxDd65B3nUE3d
SNvj+gKNkhLrOh7HK+QdVDCN+HIWw9uA5xMPNW8pPrYqMPC0NMPMUzkBMhopMwWejXPWhmSanNOV
7KUQzv6y23F0VAoNB3v6RUSS0Bx9dxGV0TKlyb1zzX3twkOaBPAU3RlIv0mGNlwalndGMjGc9D55
5RTZLsv0uo3guLjlw27rRMf3zElfMh0SaIM7iu4OqXif7SMKL/rXDspAh4P011Io5+HIufYM2r0E
uRYjtCpJnViTaS3RwZGPZOOrQnLDa5RX10e7q8JyHGFuCxmI4RSFQRqaC4HPYfNJHZrUgkoqBjY+
PaUlOJBmdED5YH6U9qs5fbMmt28M7QIfBGNgDEMARz/E+sffFRSLhwiopqgwj0mDtVlSdiztNNyq
OnzlHCjr5Vyq40ddkIGURztA1FDohUChU+NkGBvh2Ybd7cwFtpz/d1pQ0LMiXSWb3VTxfaVbO1Y7
BtMG3ODuWO9k3YbKPCOD+bbVFXNtOF6+hKL5gMJeGUPEVRZq3kmny0sfNixpUVvVPe7vXk1uKcWZ
vTd8d5aqZEPy+R6+3GFRlHMaXB8wJR+iYI67PT/VHFS6pO1r2xgtfKo3dJMn3vb8JbJZEqYHXdVV
fpkpPmEQJMl45H+Q+ivugxgkyK5HLy1dCChRIXPz6cA1RayXNinvDG+5OxGMDjaUKkUsrOKNloei
OwkaqXZ9p7jSAtMnn1HjflWr5MxeJ4myQkuPivc/ocJ/ejqK4uX5Q58cPfAeI/QuvYq97WG384aI
9JV9lkKtq3S6d6ezpi6Si60j5DuJJ6Q+lBi3UKxIyfV1CyNDYGCTkJdlComwofS/mz27XVa/k4vi
6pi85orUQOuo90IqYCYWTAitfFHuWc/FaIUe02nFzZ5gHw/lR0FGPqu9wTXGHQC+P7lw2zFLybx7
7kFovvnIyXRR+yQVnSwKAAvX2xPJJTfDQ16eONCaZpTvuTooHheCC+ey68u9MmP6e0O1NsuNQIUf
mVYvebkz680UUk0RiCxdjAjGZZApkFXw8n5OE/y24FP9IyDwosXxsyXgDkDUvnp2Zxa7NRMo+rK0
6HSxmzhLpiM2CTD6j7MDbvytF0X/ZOr8vlScmaKAA2BeTfkkitmTbuSM9PBWdKeiQJyiov8Y7CK+
Y3bD4KXqw/hdTRGoNcfYqZfd5n2movUqLoe//6GfmKKxWtUA6KbCAn1vGgxKW9YIvx6eDhdM8G67
pcNtRgQT62D5gSjbSrIBFNbXuTTE9jS3un//mL/e0uol1gGll8+ohTtk4tUE/iqL5r4/OevGMifw
d32oJ/xxAGISH6nMjTPmeS+f7YQXYBK3/0oLQt+Lc83/D/p/GuWM66gIgQN6Hv4r22P6iVvhfc6b
Q5EvtlxWzmdB23zFCYOlUTdzGERYfv9MF1T7OdI0A8mamFkQISSD1B4oYbhW9ALYBgxWCm8wySL2
MW5Sx2xUahuOVQQieS4WiSoJ/KP99kGZ69XEVhtLNoAtmCPmBLcaNZT5bqNjGcSgJVWJNQkdqgG2
QE8gIRe3Lql5M75Yeb3bUPuYDnnAmLj69BQbf9bRjaup6C7C+9zXJh8H4gBZ1jzbGZPRoBQc7x8m
14N+9w6/9Vy0qfF2/jo+Bj32ow1a4EjgLvyrOA/lSd7ZFz7Gu2vpt8P6wnd6DpRbPMZyj2N/+Kos
RAT3uLIuG2MFMoxY3BBBsN4Fp0VoOuo/VYGmDls36qJlxX/pFAxPLQHdgy9Tg/hMEvGllejQ0fJf
cs8vMev7n8OQUxvg2kd/qQOLHCeuGHWhg2ci6WRJr+ru1E9E+PYEFuPFMaMaaKJO7neB8JlJpLKE
rlSYAC4pZUPAGlkP28TAxuVCP2hWfpp829MkCIJL7wKyxQMZgVf4UupNvbd4nUR1IRGwfN66k+BW
AgoLWp3uaCZfuUTxC2GIdrOF85HVmqDqpBcmtnToahwbyCsDJOf+50CQEYUq7jS/AvfjMwlqcdux
cZhBzvxY3EEKEc9IG0P301L7KsuP1JAHmCIaxTmez5AEHVGEf4tMoEhckkB5tgMjtHXqdnkOrhzk
WbQvKOByu/A3UgvpDC2UswQ7hpdfBS1OVUKEj6aNC/n7CI7+E4OcoMD2h9ynrNMHr1xxJ6LF6ApB
QEQTNFo7TybVZ9QpqWbtzNlKUcBH2BMdrBZ9TUlJAGKmqNqeeCRoowZJdj/blgXGjFFcHBqtvkIG
wH3MeABA4baQk6kuoSmqmNckfkg45elhkvRx32J0pUo8yUZ1OlSilJooF/EnPectrvLlazsSH97T
9yiTN/up0qTcS94rGXzXpeqTfsnn+MnGSzcKZk0pTC7lTtYol5ACHrHEnboKyHfbjXMXigWbbWCb
7+HGiPBmsnh4KvycSY32k3S5hSmdCOipf5lc6Z/sUef1UK8WjXxAcmkj+NFCu9ASJKHlfg07aS20
oo2WUlrKj46ZhMtsGp1wDp9zFK1kNFNEfl2g313x+jGCZPBiGArCgwomYQytaDhv9P+AY7dPo3rX
icOWtzedG4ljGpy8fZOv8XRcC28Gy5Onag1mvINl1hhC1FNBWjGkScWd/D9lmtJTd9n77ch9XslC
Qgy12uDeeY1CTNT5XTIcwU8x+rwhPIR3pzo/SwvucuBluyQVzfuWrYVG9puJs2+fNbmy49hRZ78y
gXEAeqpgoat2Qk7/p13XQK1qEU4wnUyb/Xwke38P7KW3Mx9OOFHgHF/1Mlfi/laOX9P2v+H0AW3/
RJ4h4a2RH6GEpAMTNcxtoZ8Mqi3uv8Wf90TQdKPAcjVR7RLMz8Z6re+4IcdePJG8QoN0A7pJvm5/
qzi8UBD0r0kELYxUpwhv6YhQuZAXlZdK+S5CZ3PHCuuu+iJGgcIEEQAb6SBbxjJvHWJMhFZjMlsE
GaUzDCZvK6rOoFzIBscumIpG8n4W/wPYxYhuscbX1NVIe766FNN9OZOcgeMJB4hxMKKrnIKAE7ha
Fg3Ey8WjgapciOvVQPwEuJ3wyr+nGqHx5DW26+7G89FtlF9BgbX26JekPsIHFU8pPLeXuqHPOX5q
Z8pmQMy161gM8E1amo3UK3RQ6z5ofyifdkNHIvgTAkdA/8GHYKF91NfKyJmlChrMVKlIFQKNcJA5
DoUjo+fODrOm5my3ezOsMWQvgrJDlzEyARR4EcLGNEoT4zRWTyKa9FhcisF7mQt4QMCB9WzvCd0C
jEU6IRWx7M6QAfuMhjN2BRo3yOcL0Wjfnvn3nUuZbMPL+w56/GoiPuc2tqf+FQinDwKp9yJnqFTN
9RHJwCCnRLLHaeVTeve44ETK3P7WwOsk31mdKvnn/w3S2btBSc8MYbsjvpmgT/fXGFmPz7oDROaa
AdOLm2ofJ0bGKeQMU0KUH/xb2uMGWs6yyR1ldk+ZwqW97ro89iEooHL/+wYRdov3Sxnh9e/K13Wl
5w/DVWJ8HiIbEHOCSNH6dTUNIEjqpjqyl2zgvrmzHBh9M+eba8sQ4st+ZoQk0PsKbKZnR6Ym6fft
EsL+Tz/MudOCROksFWw6/0fUf+rIvGDwZflstrsndscNiB310XLfdK/n9hi2ATmNdY5XX9dSHhtn
zgb61De8VXKp7wOBWD7CLNONa/Z/TgL5hhN0C99DINAKq9LyYnss5KG9rEZ3GZLjWe9THrC4PuFt
EMrnU1GgCEzZyemk08uwUq+Yc5u9sM4txQSouAdOphWDCR62Edqr8nxilGTx1ru3AVSn7Jd57my3
5YB5qxjIwH5Y/ToPPDpCkX2KbAZyQT8Rzt+gMfKjBqk+mYzhr+NsSXgSrVDDg0Nw6Mqkq1O1RO56
jJQlZXHX4s17kE8E4LO30oiGZb8HV5VFlitOQMepp88irBgxMLGMXxeiyg5TXi9A8OqYksXq1ZIC
hWESMW+W9mdStuj9m1XKKcjZ5Q4bcXkkf4dfTNlZh+swthhRh8S6WOLDg5M0FxFwi3KANJ2nyqEQ
Rkq6SKXkKwAjxKwnh4gfezytnOLfP8Ds43P446vilr8uLCIhiKFoxAuawhTPGxQdTkWXl4XfF3WI
c7W8q8LeF/EBOFr08ZBy+s6R5xXOfzqylVPu8uH8z7Hh71Mw5HUJZ0peyKtyZpEwwhJAifmpaQ9r
s6jLhnxg/sTMN7MpQSd95Ec9k7ad2NHGEy1BvofBk4AGWAd2RkVyxCxf51UI7ohiDt3q1fiUwGAN
ZoSKWs0EQpIyPjzivoutZ7EvqkN8oBRMhhKLKu+RB1x1tV4N6oBaOH0yuckX1Kd4lUsnXK/KPzGU
E+Leq/WLaCRBU9sI8mFFM97IBv0lEBPPX9UQ1eniZC3SpGW5U0+Ai67Qau+S7eFuMMdWEBZDI9B3
HYvFNUgybD0BXxWlEXLc39EyGEiKUH7OBbdJ+4XCkRA/6PFdbLT425uexpZIUY8OiBxfSG3n89xA
LrR5qL0kI9oZ6+uKjcVvAMx1OdUAXbmZlRpJ4LR4n2tP8FYhCCz3SpH9I4LBmklq/Ef/oMPcZNQq
QW1nW/JqEhiSfn2sdGsQWUQwi2QliVuaw9q1AIy/ahT9b4QQ/MKhsqQBf3kFBQpZ9NxaylHD/4EV
YBMDDPSH0qLPda1mFXvJSv7en7UAobWbZv87Hr11oaFnL/new3/CeD5GJN3P7JELB+ML0unKZ5n5
YEIrszjwVCEcCLz/rAievR6nn4wUlT0LCxcmUwlhyiOaYlVxEk1H8htCWGWfY0ZBhC/ce28v1kXr
xIPpYxyu3JInm87CsgB5QO1rQPL/t8d9ix0/va3qyvLAGuT2U6RpAuITciBYixCBZChx/9teyiQ7
IbhTL3QwkvYaB5DDkvC7cWBycahG1mvdI1d3zfx9IEr749SR2wQDmTtNwmEPcKG6DebHW1YjAVT4
vB9JZFm/uE2yl0hN834+rs+zjPIhJ49ym2u2LXejGQzxjmW2Ew+sVTvnOBDEe6H9/tcS3cHVyETy
pn4tU57kaT9JRHdoMZ47vds3Qs6kCx6VI7t6nSW6KVEk4arPbvB+JkgvciOE7nQ/z540kMs2VphU
UOFQppxaM7frPJoxF31c/wcV/9Xbt+65jl+cyK1qsWKkyal9aPq28nPTBn1WwHzi5Deg83F/vJsr
3fdi3NnOzj87f0W5TGVdzG/hYhu2EQcS3q1ag52yExlcNEfnh7eEFBA2TgsSN26ZZLpMjCrOq/GP
FB/3q8GFvCodL1m6t6CgstBDMSusU2XIPQ+NV4zNYPUYqMXUdIshO/wkiFHK98xsTDnOf4E2cX6L
jRQwzcT2bTJrnedDY8D0r/34TFxhQAfOWGwy9bz61CcUZcYIb7TBpH0X3kHIEbvlJ7MqGZ2Oa7KD
Fkq0yAO5z4t07pLnkpaQajiKkNKcKEwgPE0sN2W4pJBWSNfCkZW2pfVCRpQv8WbiGSs2rJIg+dDz
xZ9v0g9TG6gwevjPl5I8hFiySw9W0z2RuR/qOdHsZjKtLs2OhWI4D++FC53PVOaI8hogGiCv1/XV
5cRxqx6D+qUzPoYLORgC9ncn+fwUq4LTvVoKAvGzcJGomwFUMT3IpQb/+xiqOe0T5+OWzt6Q9TH8
+WRqGVRZW0QJn1Ax6LjwGJC/3R6QARG5AMqeSq81G+Mb43ixTlSHdT3zNcvnk/DYHlnFE0MFnJPb
BnIapsPlTP9BHNunbgaQl6uhopffAvpEln5xJJb26IMUnHP5WBARxVIc1Ho1NG8oRfINSDjtOvVz
9ZBIeRs903A/CuZyVZVhrZ26UTKlBMrwg/fzMq2ULEyqc63PY+VoF3bIqd1YnxxFNjDWHa/26sJU
rB5jFJaIjYvutKSrsROZ4tm15WqROBjlroSaKQJSw9Jv+fRwG+fZIWAtxX0UImV0Xpn2e9BrS7Qa
3p4/ERtpPlbVLpZo2irg5OLLDDJnRNWEvtXppwNpHr/tN5w5RPuFAwBNSx0spSb4UUN3HRh7fFBB
VpuikMKCsAQREdjZQkN62ykCTh8ngKx5nBjGjz/82OywO0v3SJBJmUGcLm/yLaBVYEh10p8Moqgb
vPuGcfwcIiTLfCN11V2cu2sXWVpB2dmjY+fVanAzbZNLRWQEDLavMlfR1pxb39+rxyf48FvCIJuA
eRvKmveIuRocu+QcrIPLlY2ivEIJkXtsLCkCRX/Y991oxupUhSycpBa0YbSpAKxKRrIM2u1CDkPt
IZOwbA1saklYVaw5rxorj821IT383M8VZ+367m0eE5n17O0aOYsMmzikQ5MNDmO/lB7Ly3aOZzEk
RqX5KEayI/TwMCfP3bp52sebYZWf2tKWHKI1Greu1NYKSOWdfSyPz+AhJ3LIPdwdhXh1zriv6+K1
meQJVssdiftbFse6WdSr71mXS13Pw/zj23iNycKNCrqoBG4SyGmj9obe2ydzgQf1XNs3qROn2cpE
Dx+f7JWhLAC8X/JrPQXuCrQf5CsOOMVyr8Hm5RUUNPE/GrKak7O/FVQ5YRKth713NgPiZuR1OJRD
QYyicFhmnlA3d880/GLBhVBjIspX3gE/Y4GuHauc+D+JFdEIUweueyM8ZnlhETGn0qX20p/kjVGA
MUs4K0bgat6v4FYlulzDt+WpGRA0hpty6wrWdzoYCXKsohkOQ8TJyfh9ltf5mx+ZHM3Bx8/23/QN
GOr97W/fbB6pjR45ggspN2fJYamAZ7tw25zOlpLeAnfX7Cfv2Q/D4P/OTCXBOwTxhIbKrOKxn9HC
ns3ztVKPi3VUHOugMiGWdTgNP5epJINID67IPjJ61PslPz7ttw49/jRMWoZPrz0WJPRfPQIP/BX+
GZLX/dRz8ooOHobI/qGaoE8wxi4Sl4bK/zxCAl/5Um1yIO/oMlq4MyAi+BY25rWsLRLwOboDZuf3
mb+tbCZ7li4bp08kXiRlqU2y1ozWBh6GUaVZ2p9E9j1CnEu8b3vCf6atsMyD7MZwbfSrb63uvoTw
3LLIzyVw6N2oN2bJh0/O3bwkx5kemmCI+roOBKaJH3zpIAuOonF0RZtXV7/3oFn4H2kIk/mh86Qw
3avKbmdDKRXfS6REBwba5L6uf7EYW1BAGmtGvAOII25IbNeRykUsiu7H2Zj3hWZnTevWVUYyM2fj
ZKT5djO6ovAwMQNaDOf+91/wD6m3i7K6dNcFOZ9BaDbBH6btTjxEwfLcKWPUVr++M/f1IDKrFclO
S3R3Ct02z6Jfal6LM/DY7QAyPF54btuFWUzESePhuu6ob5YAH4uBX5soyjN17kYbbOMpbuzEdTn8
UPvaDNM6gyaMxeVl5YiziDx34WMx1pWVfcmo29ABnNhKbpr2Xyil1gPs3jbUuwN4LH0iIAFk4OYT
zHfxNGuVtfdkK43T/wZzjHV0ucDSJJJy4WFvMrTB9WuwMKO40f3HdpLdKCVdEJE91Pe9Ma5zjzgM
XZoLCTCXdOKshlQYsNY0YctCoodYytSXhrUp1+6SVOH/be5qVWagMz8KM4oRy+WiYGOFcLFVUAIF
Nc3yAUd57+/Dq2kKScBvBLq73r3cBOnywaHKMy9WvuPxP0vQU9DJwwwdylfwJxDvUG+ag0tTGMK6
BAeEd2pCgmY/RAZZ6wy3mUBQDiFyjYxlsEloPAAKYoP1q0KVtTUh98V3bmDIL8DpizUufMRqNoPy
aojNZQkrAFEtEgVT3MRxBYRNjpzI04hqlD39ukFjpc/DNmVbAb/qvcDAymxA+Ro2WCF8TddYDjQw
6Eg/LlDqgrtlM4lMmiQ6Ywr12NdKf1i+44Q8tlVxbPjWoZunbB09QFgHAscYDeTs6ERtSvUCwhbl
TD0zJWJ88kosJjtelNlwGT9WjQv9vE0HmFrw9qeWcQSY8wsa56cnbSTEmYxP+6IQ1bi2LDDWSrYE
numGGZ3g61Q5+H4xNX9Rl9oAtfAPB191EwZ+P1pLyw10vkJgNBMXSU+TtRvpIzLzYoCeV+KVLacf
kJqYH9zNayxMEEfjxXhodenfT1ALyi98iiY5in72WcFIs8L++lEeGkD0KBjmMU09eqc5285dEu0s
uNgv1UjjIevhD/sm/ZU8oczNYu/Y3sqp3vreLoFqVXHeEaKx8Ao5bxatOra3cfHZpkM78BgQDdnR
KdnJZDgFkpiKRLBNyjkktjbY3bjh7nCpC83KVmzTI1hN19ofTaihPobWcv5I6W/bes1F07qdw189
OoVs4n+j4qMKVXD31D5S0EONIquVhPfcl/+YDjrRp5k5AC68eOXkANS80de2aOrsli5e8z4580Wm
vAw9T/ipFJBY5sHGoLyMtFqimAWEIYSEoYlpb/uGIsHh/GcZSRxxVnVbYuaotuWmfxceJLscEXqk
qYEYx2YOW0n46cQq9Y0W5I3clS9zfFGF3H70WqT+sunO4RhrqVE4O2AimlvpJ6x+TTg9+9f33wD3
xYIcOhmstpxLT559EhbMfZOUPUw6ZYyZ2o5Zs0ssBRgDkrswKGl6yc/zaacgPNuAwuRlxjVbymuJ
Txj2HzqlFVJfUBIW0VbVY8DDFbTkaOcI8kINwu2/ND5wqETPFwQ1lXHw9RIesQx0wTGTol74c0fz
9aXaC/P/LUxYX/FWTUko+AyPyAGKnCMVGwKxmhLOCPFyi44gnc2ygQEMnmk3F7QqfhQf3vcy/YPw
Okcd1cgK/RXgZ+sQvt+ToiASeFtDbjk9exKrNXmcD016qjOTlM8pkZOUbXiTdcADMn3nwIbOmrB4
TaaYLxO9PSKpNud9MoG6XAlKkkzBZeMDt7S4mNStjS4Lcp+QstWCbZu63GY/IRoy2eaVZcFILt3j
uaVVBdBL9sVyXIp8eK5Ck0IAi1GWQgNW8AiNJBvOtok9yhhQc2y4s0sAE0naKbVAON0nQ/OIY1YY
c+xsiD/nNdoFk3pGYUdnUFy9pdsrwxsjY6j+Jk+Sp3X6NpEisJL5gcbKkgbDHmtoS4KfuV4dachF
erqFuiQ4wgI7Mdgik2F8HANTIivanHpwyvbQ63qdFSm3YIQhVcX9dbUp+dhbGZUicp0trRz/gysz
PzIcVr7HjOonQqpwB7PXpcwz3eqRa4J9IGlGgY7TtHdzM1c7rVtBqkMpgOSVNQBZ7CwC/cWygSUl
8AkA9ZHu2nSTqGQJT/0gybilKqGNieBXtPyykwDXsWQs6mKy59tPK5TLGsLPGnn03+/eNTNRz7b0
Ox1JGMcjJDDD5jTNRchbFZvJ6/6Rm3pRyCI9WxM27WdRfOjmMez2XwQoVFqV3eXS3sHGo9cFZSoP
aq1zLVp1gnG5yJsC9xMa/XrY4dKB4wrORfHjp+Ji6Jt5MlwP5uQD+XVTgY4f1wLfT34w86ZYAJfv
ziiBTfA07d1ij58I43HuAocCEGQubzwLKQLDROKGv+pCkSD241Q2CzwPWYfJ+hDdiTjoLNyu/sKQ
nuOOR2E2gVxfUfnlmVjUNkZNOhzIz0GGkZQZyWYnpXuj70pGES4RlGymMy9J7X9DjVn2fhyUWAFq
oOSzPM2Qppl1GrhjVjKKRCX3yzzXKKeVEYgyZ/2beVzICSKURzmXIUqMGsPVb157VVn4R4Deg4Eu
3hBAg94bCOc0F32BPqPSoB8vBeNYg6aV26W2Bz81bIFMWEIfUjTUQhEdhIVQ0E2JMOBIlsqPbRbj
SK91qXdCubOjciyzIfP8s49/9Yms4iuHX+fr4YdKNNZWg+3sv1ChdLcVGd1KJbahMemgxENk//hT
VWvs9IYL1YnVsjkOYGVJ5O47PWtEsfTu0B2RL2dwaPcurhioRsS4y2Lpj6z6Zglf2iaAZvcsFiY+
kRrqpWCQ/yx4Fpwn53A3WdIg8YAvMiDf4jZfwCUYtXMWffuv7Y2s27+ijMYixYWTeA2lDi7UzfsH
UhWFtu51Jij2YdqgTXgf4rJz2CVut745/Mwk11bIEzqyDBwLqr2ortOo4wW/3jMsO5eKrPczqaSH
3a9zG5vATr8iBk6Y6aqWV4RknsprXAr2QgCD4zZY3vBLYmIZgqVeXVXlh0z04uFtQbD7QzPf/rra
Ht9PzQ4LO4Tulrnpv60YOtBAtjd/Xl6Q9Qay+WNdkVfZS1NAVezWWDPlhJVz6PU+x77/N8R0RDeB
C0QUuDDSGJ6N2mo+AwKVdoQINe3wJhOetaRJuovhQnCEuze20BinPcBXGvcIwzkS/MkKrI0npu1G
KC0njqBev4iPh6wq8CJsOowqKa/tnYqbGSmXYMuxtqIITOaLqFXIJRxdIh1aTJ6gJBqMTgP7U0Uy
Yl45uK26hB1t0DxbmuDXMC4ZVVaVGvScGBJRCEL61yqZP5W3I/yshagcarQ/YQFZkloRxOz4VPBf
3X7UPhe+A43rljSnTKnqOiNvTk2UgR7rnRXRITeAAtadkTfoUeZVRkEpcyoTC2bP9mdlIyhk5B8s
MTrrVG/4wqYoOZVNjfKkE+j1dsirj6VpJr1MkehcqblvvmzwMn1nqGMq/ytBYGb7hWy3f+FiFzE7
wFnXh/XfZEKFnu8XS1EqNesAMi64nwohQ8OgqRwN6NIqFt4j/EQpYfFnS0L2D6vXUd9MiV0eUM8J
gPI4WrMA7vjZNERgrXMEO00MOu3fg3bEwF90rdTjeT2whOqOj/f3VVUkt5QPALaYtt7X4eWdi0IZ
R+L3hP4M+1FgZwazfm7xxOcL6wKr1iFJbdYVtrQThq+GEsDVSGWXo6tw0iVRkAuuEanm3qr5VQHJ
h7QdIyzEX+IPxmun1nh0Edy1i8SUAdvtCLmUeFmRkZvUV6ZcI5tm/f9CNAnIlxrFi+XqC6KQEH++
J/P+Gj2cYSSskQfYKOGs8YfZlgRM4bnJ7ppJhaEzc2s1grao3KzOUSJqj1oSAgvSx/BJmX59y+LW
9ScfnBe+iYSz3962bRvCW4qgm6ltTKDMDejUvHpb+qRn0tqflpq4HVuBql+gQl82TOmnwMn1UK0H
1KCo4OVcN0aHkeBva18+XO1DWyOLzGklZnfnKwMkNn/JrxkjNHYvwPV4uBQ8aFF24Eomrk3Uu8r+
RQ1oTXFASd4nRG/iSxCYm4pMoZOT3ykfjHpiHHmvH26LBuQ74Q4C7h/ZxjdEB8nFOoDPgIC7X/Mo
qyDr7RKXjBL/5tJGNtlktTDXJ2O9WGkCTkrcSSgxVdD2g9ThUtLdT0cMpcwP3JYoVeT+Ulbl89W3
lQ8eRAkQiRsqQ+6gTnk2r199jUzknFBQKfGM+d/FrgzA5oUj/3JtIgvDiq+Ei23utkE3072SvoAi
RE3VastYx85hPyGhVrW66o9kcgUr+cYagRFi4Qc8SKXPw0cucXOXGOh8/ukY/lsNXTslxRNX/DN3
wASmYdoqs5ahkmuzax/dVSGtCcdzGtG+cHRO0I659rYJGkWN2xBsqrDnx8gvGdpjati/W3GuF8DE
VFrq7YLeiCcMWtkMEI18GDbABnm5cPfyobjph9Vr7SpOAls6lfkIGaObf6ywFYxQ8LThYED7I1IX
gAvNHmVP+iiDm32gdcm9lFh5QfX9Jjh2i8yge16+gl7cmtT04W5Y3cBZUU7+ORTMW2Xa4H2KXHIG
jiOxVkdeShT+GxxqW8d5OjnJNOtMcdDUmeePHHXGtJj87V21jvXj940vQN1jnO4KZxSx8NRtX+d4
TI4t5jbawodLNUWdxUScbcyyN10DeubVuxHUDcEnR3Qk7tmVqt90ALKcTUTGn6/H9AEm/iPsI/um
500Hg8rflkBFnJvSy4ZxuzoVemE7zowqVI7HQu7bgWsSAGgJuI9CbvIQpmpfRBb5NdtFilNYOwEf
J7AUn2wv7xVIPhTpLjT/zvETB0nIgI51BcREruoN5g6i1sk1H65W/O3LzEeIGRwtwm62iQYynkOe
HSikEcGU9D2imjTnhtRVkp1P4NlBsSyj4zMgBTgzm0PY88Wb0IKRc2qaDTqn5C2w9qDYPkhNrlb0
lpib5Cd8DlVipIJa7N0vST52utTj3VkE2kVROSAOrGAQqwgd1w2bHSBGoms0ny0xSMmYAsryjt0n
7E7AeTd63+xTC0lE11XdwnhbdJtuAsRQVB2r+K6TykAUZWSU8MLokGG74jv6LMAgDeCq1LdmI/H4
2LaZbhkNmL1XJzCVR1nBenKj4YlwwezCHHCgF8qJVGvMUpaOBok2MT0tL3istxtcbXz52FJFRT64
1B2F8evLtiakx2jG938Ncij8de1/c81a64uOY/R43n9fP/YBXSy2rO9fP1sMd3CmTPYesGN1xaZe
ZPRqwuYMITT1t8QMyIUWXX8oP3vaQICLeXYf1qAOgQKSuAjk2q/JQp5AJKUw3cWjj+N6gQcYBqt3
XMRY7Uny7O3f4c9jovkLX1O9RqaUcNhg5m81fyNzLUFl9bYQHRJTtMZuVWfyUKutFGqLjq/ZueTj
cO6bYkPqk3AtbWf9Lr8Cj/bgK6oeYNI201qDzBYSrMVOsugAlEbP73I2Dg+U+oOKflOXMhylSlkH
7na2MWV81stqF3JzvYQ8VH0LA5rjWWR6NUiwydRlGT2huddltweoHSZMtc9wP/NHmn3Ke8E1wIrs
pXR8RwKOyg6GvsktDohUNvCCvzqIrxZOoUfsNO1zmrZ28gUUUJGQNa4O3uDk1+JHxw0mFKTwpvRY
ZzgDZA7s/GAVIg1o99pNq6XFQWYP/iJj4LgIXx5YTpxTtjGjFLT5g7Nsnt/vNHrY2YhCmGwn9QJ2
YYxvisXquVdam2bEAlhmhhjhDWHMI8zop0fzEAbgSZCI5CoasTik8MUZ91dub7oDiHDguw+0D8qb
5dqkz1mZvhptssOgPAvOVeaa+kQKS4KB3nDxOx3g9YBSdO5bZHb8w7PUtIOxDH+b6KZ8HJEcVDKL
yK3nrjV+fmE2VKpJ4blTmQV/m8HOu9FiJTkaTb4D6nrTKCQpcBS/2rbVdEA3++NvIKONWYW6pdnH
tQa8jM9oVM+t4IQCqBcAdsHy5y4PzEg2V5iKRyy7WbQzdfskZ3bqA9/Gkq5W7oj/O0dduP8WPWSS
nNudUvfcX1xjPNG8QuwX/VhNxspfm1HSTRAH67AFhUgcZbRZYzJVpmIkxKOyzolhEUCs+G22a4FG
pmbSXky70RykBLHmT9JRuby6twIojAACRKJoidm57l82XmiAJElB14jBntFAkdvw1xOPY+bLCWs9
z6EkKOCJKrWuOWK/FFQ5C4x7wwZ4iHcYowT+ZYPEe48uZdThmuXJzeq0J5c3a/iVemKR5AfQ2ts4
iOUus+xlSI8ifG+6OLqlzdwbzWlZne0b65d9k9jeW4MHq4zhNMnUSAXT+7uD6o8h7AXf8pmoJNn7
VyvuRMJTN7keu3JlF6vIFjJzXvMnpwUDWnvEiqGYzeG9RPbx54CKF2uEZAltSA0CvfNPHYFV/yQb
INpE9KwbnYxMj/p8pFoQlR6JlO7IkKjWUNk2Szua+P9ac4Qu96vjeK0plQAmQUU1/lJX7urWBwTL
EuPZw9ejprsaygqliX4K59dICum3oZrcO++MuAHkz1ajaHRVI/rKOr3bQRY6nWZ++ClKgNWcJoVG
nAlHusGNgEodxZy1JcOyINoHZpUshjc9utbcA9oKP0GTOncL0ifVCXSAHm5HCkQoinoGyWmljYkl
hTy1XUa0bBrNreuop7yGNNTO+YajWAvbtRqtyDmVGzomQW0U6Ih6DlTFcdjRfn8NOvGxK9lIJkTq
Z8f4GKhzxfpMhszwSEJdQ4DL6tPn948QN099U9k8sDxkUGmyI28lhETam82nh4ppzb8xms2NBwLl
RrT+xYal6xaivJ3RfO4tpd/zCaIukzmkyxKVMKznxNz1b4AkImtctsx8RoDwCQNujusS8djfOBvW
gPgSbjS6HEfOSvI04xiUT6WCC10hPMeI93UZZ+AdqtCCIhbTsXcMNIPUfMESJisM0eAxiumK45Oj
tF4lhlubMpqtmvEKROIEoUNjq0HV7Pj6sfZSrDX7Q8VD4GMykOuH+af5hbPvoRGpdIqQwGDhvzWm
BucpNHZsmp9cXS0aufxCsbcJLCbLtPuxeMDuRmiwgPx2+OEKRA9nhuBojkBsSCJ+s3s7uYTtkFX3
T3G+z1wJJZI4K5A/4jBF+4zD8bJW5j1jj7Eql+lbdcFvjyCtMhrTc/dfJm4iF3k4O9mqbwu0Pt1e
Oc3c2mTuH0wkcUrjy0ENlnzj0MEi8ENYcJCyTcV2KB0A20M2uTejrtozvYa5PbWvRzJMUgeUIQM5
+/GC+eTLn23Twar7FmNtOSglhlGpb7Yv/60uBeaw4BUI6DT09goqWGmueAyBRtZRKkn1vL01uj9V
ptrhzrAj3LpIFlKLwY+E6+nM4bFvB5+72V3WjIabOjBG/o1Sq5+1R0dxqvUL4bZpL9rT4n3FSROh
uHcSyssntu0jkBeA2wlL1usAnTcqz6smqgAq5tZtXxabiEBcl07zlbfAbc/nHfXanP132hK4+aGK
SKNjBEaz+f8vW9zJ/+BRpnmoJRVdqR2KblC6H8nKQRX7VngNpiy8YKYu2yg4Ucxr6jpXHRABiLlC
RpLmETxlKYi3IYyeWN5wL/dkpHxlRINBNiR8G3HjHMupkPeSIuPgFs7j6PP7MHMVlkp6vCO3xEI8
PBob8z5uMZK0USkr9gMTpiccM7z7tXIjWojj489FgtMdMUO0Ss72RuSYLqoIX86YZ+ee8Y90oo7F
KpwszEC/5onDLQQCOJOF81D57A3/OQHxRI8h7pnMmya7E9Yv2EL9XWtwQuKKd+vBRZV6owJ2jOyu
nwN2zo4y0jFZoezUEugDQBuyLjTbjLHatv7o+FNjEuTEwndtucZn5O87ixfMgKLCGBhgsGqwxzi9
APBQ2+3ZKFUokKyEGCjPLsWuMT7FGhLOgAUVrlPk5ST+O5n6y2A/PivnZuvnDYCUKoAdWQvcHztA
ltu3TFU3rtsxwXFdNozXZ3549HWw8vf2GgZdYsvIXv9qIBRUlC+DgZhBc1Wa9FoPtYVrdV/672Sy
csxpg+pzPSkiNAg25Oc+sROYY6/sV6l3BGUhAN37yJ2Wn9k7oNpGEeR0dUtacGYmvunvtqY9SMF1
00RCb1LBNix24QOJfS8Ht2fgIhbpcs6S3RSscof3hebpLsQ7imN1M9ViWJ7QvrOIIjKyqjeNah4y
rgF+gpvPcfYooQHy3gUMdh2ob/jXjz+7JemJoCfDDM4/pr7c99vu2ea1ZdauhvYzok7j+9aRDYeH
KWk3DKW65PNkn8jZpkRNIGI3epVIUkGYE8vneZ2oLtseCfSnx14HY1YkxNiig5fOjhdqYjca7M33
Agg89bGrcjVg1PSbonJmK724InlppPAm3xV+znTUsAY6P7gdNAIG2oZ5wjEXgPnQYp0gtew6Ly2f
Ibm1ZfMeJTp5NxvZOQGvxWM83FPJfHX6owy/g+kHQVVSv55hdkuhFIlyzXWCS4V1jNH29Rg2slWV
8KDHbXtqzXO6EVEbI++121qbApM7D1lcaRdvyefjLsCmFLxsgTR3KYr8+jF1V/bjYKzRyhLXBqhO
336UpgGukNN23c7C3sF6z3pDzFFO2b/oA+ujtOIkKytCv/J0poESbvbf3uj34JZrqL361rQktVIv
fXD80F9QoZKrmC8ttYTqp92tjpZzTBJawj6JDzMI1qB3I2vQUtdWdU2o869r3xI/Uos/x7vhVBaX
TRbH1qPlHrWr7cFNUi/mK5ZLebvfEdf9cSrMuOFVlP2ngNHU2jTjpLDv8nG+OpyrPbifZIP6GWd0
2ekv/L19+eT7QC2BXQUYNV+QIOZYsw1iddLrmdRalxOI7Q0uSFu71psC7uHazqzoZj6Dw5hQZXLg
YA8sl5Obw6J3dTvkUx9ibj4BqFSL0PJ4rE/Jk+VplggGWiKjNQg6vD0gc9HEdNWzvAPSfs26d3s+
vw8O5gkXzvycOYNF5WtakYUujiZ677H1ezG+/m01XbJscZ8qTOiu/UXjO+mpIM5YLbgEg+HnMY4S
QQb4jZn2CiOqNKq+sUYhgH69Gs1rbN/UdUV0gHupq2RPdoiwztJzm24sJciB0602sEDrmk1uiBou
pl+quSdupboUjqyaGzobiCB5Iy9KSOe2BTlAGoWVf6zsixvnh8P08IVuaY/4KSpB8pQbuX+YctV5
XXcL90XwCUUIU1z8qk6AyQztv4gD1Tx8xM1/CWzJDLQvnH3anfg/rKcaN26qlTa8Am2QNGOuw6Aj
HX1MbKJzbAyF51jv4zFdQdrbkyaLPjjSYLU178Ojbm2XT7iz2XTkEc2YGMfjcOsIq52gpTkmIHcm
cMlzB/D/6lX0n5nzdsHEbMRUe0caQw1AB0QOoPhWt0hbvvwhQ0EThP0mmw6Z0yydulkXIcu4v0g+
GG5gmLmYnw96W1ao2AQ7u5v3veWJsalv8AZIDLwwbDm1xRCinXp+SjMGSMUDPePt2uoSXP6yxmGE
ReI1Qqkj7lDE3ZMGJfHkDcekuCsDyVvnGll6TZJS4Yd23bF5+4umeYckwnN6KP2bI0BiUATVCTkK
rz0eOkB94af6Q2e2QyAa1sfqvuM1BCaBciqOTBTKfQ/vz5/odjkghmYZz6EIHmJZIDBBOLevYW49
cy+Lo7XX0myy0W1XllQVBgqdiwfEUC/JSljt+JxRIPdzVtdqyUay82x1nPdmmm99LUS+uHpb4Oyn
Li9i46CAqknV7qf/mdbOX+eAQ272Z1HVkyHHTcOiaJxYln1OuSN/kon/DAMHhQhVW6BAdC4xu8Ji
S+gxMyL+UCf9Ja73N8V+gUNjHlmW9cBhX2ucdJSyks34zsDpktY6dxtztrXx83p2VnM6x8cYh94N
LXO8qPddxURjpMPAnIzbqedY3o0qf8bhvDUtlB9egEUoHu61oC2QAud9/CPX8LPMyKBvW5ZSIs+V
27QkRKA9Goydw1pwtggo58CkqVZ78PvUq9PStD6eNuqvUAPYwpSz2XzJ2nFVR9POj+x80AihPiDe
1/ePWd70ur4ZcOYaFf/IAmMTmSDdDK0yfXr2NFsl1EvRnyxPOHOWM7rOQVUpXPFgp4LbDmaRzNx1
mopKT1+iDkDjHyKu0bosr+1Yl8YYrRpZhQKX7CLFWLILAfIETP2HWxCAlGUHqKE+t9LUFsz+KC4E
MOuxpGAZa+3K7UENoa5elZPYOkGlqCToLbvEwqNwUJe6m4gEonuYKMCjDud3Cj+XvdpChYuIdfSI
vC9veicdmH/9qW+OCJ5UCnDFL1+bUAzkO3WreRaS90LiselNFKanxT+bpWYqwAA7P7oJVGMgXkIe
abXg98ocWTCzXwSeM2eYS6fQQKS+0vzJrC9wU88FTOX4wAtA2T+/K5Eu6TRc+pSo30GTP96b0oNI
MRd0LCaDHiZn9mOFvjp+ZJR5162K3OJ1/IqSkq6RmF1MAnNLXTigvtbfJLrKjcLQSu2EB+NyLubJ
cxjZ6MZRwYVGFQlTruHT96zptKbzZFPHuFt6w4787Ww2oyByLAr4umCHiSEKJ8YsU6YQOEbsJRHo
aBtbGItn4yv/IuIof2dtJ5MI893kAEOj8CFr0K/RgaY5FLIlfLlBHc+0GqZhdZzy4ayZ+yFWecRP
yf+HIqZOELEcQT/F8+uRT0kEI67Y3J6DdKDJG0WlC4kBTQvKEFrxzsXAM1cuHhM+bfrNXpE2UKqQ
PIiow5RvOUvBrJf5nTRk6edDVrwdZIFlmP4h3FmxaDLw5P3xUsPFlMrXHnsfaLF3Vm9WoPSrz1xN
FArRDqJLqxb0X90RBUiHDv1/OyZ6PpLc6RidNqkd2gJG3TbK/XhxTdQ7rLIO4+gJ5DTeaodRGTDB
+CrFPy9gQhDegikMy+w4ZNzwbJzZf5CNMCr3g3MVa1yQcq5DkDuzbTqFlo9BztrqhgAXwmy0SwgK
E4FAoJ+47GX188w/1G48WzVnJ89qr2GmpHucKAetLVI2UdQ0k0yQEPTNJRHKbG9bgNlMa2hQkC6r
/MPAoVbmX2QJvOMvqBZR0O6wJCyRzSixpILwn6E3WrXtW+RDMygsbiK4VEt1p09vu1okSvBHM3zf
/zYluWqKdOaNketeXDbn4XVXMTwsEu1JvGwc90i7UK3N9g9+7fxTcg0rIjt//FR5ERe5zyUxHnDw
inV+lYKFhWqT3XM15bF44+/yugvxzmYjh1xK13doagCyQvKktfXtQUfeYdKjNF2Hi5yemwUzPh3i
5KfMbAcJZ7Ov9SdZVC/Xo7fr4a8WQYbazKcDAy8lqWdr8/qXC6gBuhoHsjMHtlo/3JKaJJrTZxj8
kaxMidkxppQVTzFGKGm/e3imxLBJm8dHC3GDYR893SbrqdRmBWFUuBg5C8PnA/C8j5ebs1rm7Xgu
MUrPKyKVr+plPXx8sK1X9A4S+jgqZTDZuTdj2lpfWK0xEjpOaSq7u7lGxucxF7iTFVg2WQPQ6K99
xCFmd5p6tZ060PDl6+TqGCVosml0QX1LwZ69qalPYXQx3Hbwqga5LwaCB7sve0z8LtrN/fSYZhd9
mpRv/RA2yn3mw6feX7K2VBXy/wkwoP3jPumf3ya2ch/N4RVNoD9drp6ZQWm0qYiDOS/NAhsXLQ0+
i9jtA0XQ6OnvyGgCm+PVrdM1DMifx1MTYOf/RuBtSsx0gNZmKzLmCsxKrvuHVx+EzlB5vILuePFw
LqqlNpG6bIXNBVql6QWx0aOJRd7EN3pu17Skf08D5U2F6bWTfhKyR96NOKfS37R4V1PET/CAIUqJ
PiW6U+m4T+7eJyYH3YG688+PNmcLZRGwmn/T0nibf6AbhGfEU9JhQay/rDW7MSGit8uhI20lnhCy
YSbZjX2ig0RZu5X4+CeqFfw7bAEaHMdWzqp/dX6QMWBoKHN/DT0APHlWnKL7kifYHEh2gNSk5S6W
ag+KmUmK2jgXAl3TK8bfJibUkK+IH9o6nXCPhDeksXhoZ51G9hGxoLJg/GKVa6hggk20l7H1BX3c
4ose90R3LgqgQgA1xf6koTvuatN7iswM6ewhRT+SUInMA6J35CkCPTVIeeouFbZZb7FRnDcMxxrF
GTh1oUkoQA2FVDiwIRTHaZyMNHw8Ja63ONzOq/bpXy+cXBXDKaPtyIZtmXxkvIb+dDzIAD1xsO1h
wu+93BBBr+r1d6sTCR0oBT6sqOPifMLSxrR4dSP1iYfIiV9acAM8mXhH6q6Z8uEv2m77PPMk3L+G
LkPwzLXiPov97N6OTdfZosLvUldfB2Gc8H3yS1/ji/k9wlIVX9Yw1zOKrNcYhOmvmttVr/7LvfUo
/FVWIK7JA3L764JlsmDlwM/MH9SgEjYVRNKRlmtJ7IJpYnA633WFC2k/6RnMop8NAsVQXv0EMNCv
pmm5BDTpVl/bA50GmehiQqXf9D0bmw5VgqWVdhCQkzctM9gd0u/RyuboMKXu6Q00MBOzuxwtNc+y
e0eYDf5GWV3bPym2S1xSw5DqXzT5uxzJKfvxqjNU9bE/3Rq3ZjWX8RTvMmCKeQC+MGqqLi1LCnT9
4OOVfKG73zI4ma7/KD42H2lL9I3XP9DpfVhiZTa9APXsDrPg7z0j8faOIYyuS89Jxwy3Fe7fxtXx
P2TqIqoiwNgZzp5HsAgtycbfNCxE1gOOOYlfEUNmgHdisRUhnBvtl7vJBcN2LhIn2eHlU8nsb8HA
a6cgZE9/6MhiFKQVUnrRLxeBOELxBnSnyz+2YhYyztLI6XcEBk8ctdCe+7gFXllTxYlfioHW2jxH
E/8xOj0ww/omCG/lvaBHQzZoDNJppREHfqfyCvDhHsS1hyGs0q0E3UpkGNHnHC/TyZdLpZleRgmt
oKj0M+2iRhtdeqgBV71oq3KawtD0cFiDIpHaB7Zyv9ZwTcvoF3/kbl1faghFR5pbMDbHnJMjMoOx
fYn1PDSTG5E2gBxhH6NQQ8+KKR+fH4TiTvSzCTvZkKtcrw7yObcCeRGtFv9DHk5cKhlZtO34/4mT
+LgwTdZflg4VwzQVPIPrTIkBVFgA+VShInA1gHuX+X8tjQsm3L90hLJRNEDskA5R/3OZlI2OJzCU
AIf/aj5QyMipaDa3NSZeXBkCd6cjgIplHoE0b4RZeAGxPw2rmQIgMVpXAUoSf8u1RxTzNTleInyi
UCbk/+SXhJU6GB3sKieMseJDTFVHSVb28LEkhZTeRY9/aElDNDyfE/FEr3oqgvM7pRCX57KAAO6L
+kzm2sqIprzQv00n5pvAOPMBlbwAulk88cs7W+EjRDXDWRqZv912lMqsPsSgGgICwKfoZS7a3CRl
oEvLKEs8I3MliYxHERPB3gy43PNNwjwaxYtOQzYiHFaI4o1gAhGNIOee8iBF7/hmsRrveyXIgm+3
ye/IkiSbC4jI8RSfdf0Suqh7ilcARPxf0UrTY/wVSBDge61IYf6YQxpLRjW3oiTHXoMwzF7nbdFN
NlydlMWtFp1LOs03Qsv/jpVRtkN8ZP8WkHQBBPkHanFpq7/ZWmJ5GPd5fRuGuJJKB6QxBLWowBxw
C0m6cMwRM0/TS3zyAP+dE/GxdRDo1wcZ/iymyGPHY7T2JuZY/FgoHG+WaysNFdWxa/RKehOPgvjp
Nzn6lhRGm0+R8ro84HlvDKpRph2CoizA3AVxohgyrKeg1DfpV7DYHWwyiEo6eKrDTXPV9IGyhHRB
sKp8+I2PN0+SREVECZDxRDzFJWcYcyITHa6yYYy2wtzv0zJe92WFcr2JE2v1akmLZp1D4VC25+4x
wFEYD/wjP1WW16RAfR9OGkLXHkIbwHpIrMZeajwY7+kH510xiqVcjss6LwOPlW8ZUbb3jwmlDN8X
tfnXxR8Tq3QqoObKxz+0v3+3HnzRgFZdkh6eUtJF7dWkkX+TsG7ZEc2vBTpYjru9HplBJZKgjQ5P
L2luid5l88ZiPA9uZpkzVoMljV2P98in907Hfoxoey8VTTJrJ8ErHVMWpj+XzKKtXvt4AWyjxoSC
Y6+S3Q8wHc4CT/Asq2VL6bWC1zVyOHA9kUSq2ftrLjTfKEJOgn7BYDE6KeTRNX7w5hfpiX/IMjBS
NfkFWcjfrxDxy4jZBAUjzB8kMCF92lImggq5hC3hmnnj+gqGrCNG428IMhVAE7WPJMsa87W1gQSF
cRSbVCoB/6PTDQJAR474Z9oLAx3ki93LzQXQpWfGXph9hYyq34HhbI9xIPFj6ZdYv6Y2mQk9q3uk
KJrSFsADp3IoY248n17o4NzNnI9SQgUTBMmwsrCWlcT/XP/y9SapucV9DprHEqRsnF4GZKPdUjAw
s7HW5BpBCCCCshT734Ah9fsiJGqoqWQz/J1TxCSOb+sotq3uatQQM5SAfWKKfEKnZIrcxhrtmH7F
85tkzC3Mzz9Fxp2z2eEeMAHNnxGhJXorM2GaIL15EEZUPFLDOIIpcZQTNQXO34XEApn/Cl1Ypylm
1uN2wbjLfMHnP+FysMfQkwA55EuzS67mrepuiwY00iGk2nq3zYXix9bX6t4leDMDrlLqs+IVItak
TYWVfI8lZOq+t13Op9ODGqEW4mdrY5MascAzTwz9NcTWrQomuG1pqhUHM/wH+V4ffpAXw1SGAksU
fYtKJwgzmeNu779/WfDf5IbVd/bUsvasPcLJHjewjLo1N1G1cjNBEgt38ljJ0jTKdM/0oQZgzTy9
SQHIuJ7qf8WIZjql9CCK2BeKjMxzekUpcOj5TubkRwUvzbIht+Ghdfh+BoCtHH8B2gDiYjYP9aku
3cBI7wBxeoex2tvSUZLbdJlmuJwFpGe2k7k2tp4+l4xaZw/6fV4wywHhHc4TXNLrUf+HkwrczujU
B7n9aoaxQiCQC9TgHo48YIO0usaDLJBV8GGWdkczddJ3uWG+Ks/GmQ1wlUHyMdgDp2FW6CDG1KUW
tBoHxRm8cwIHsWNJVptsMSHFUtbkaAUOeoqeuGElnaFCw44mMtYuPiZMssdwvCYxXQQn3CDRlUFL
T83j6WdDLM0PPWNfB3oMqWbiFv8ImGCuXP/6dULnxloX1PmtdhdkiB9sy0WIOWrGn6qJOQTNn5uq
VJsWCwkYlxQDiY7NETkULFbNPKC7IkXj8GHR4OgaJvjL2EA+HW+0VdVVhgcsh0X4aTCiFNIgvCvF
VejjFdJusuBBIIpWFnBKTkFKhEQyja5+jOu7wiBq+po8ydHRSHD9E8ISwF8t99ZS1tpMa7N6rHRF
aoQHl3sGspHrkjMs3jNP6PzND0M390kdNYU5obEyXjxSqg77Hz08p1zdXVacBINv4+gWgjY4ZExZ
Zv9VEIzz9+8hhcMINt9Yn8+VH5VrZQHKTMdmqa/gxtfV59B3pZjB71Gu9EGkIJ2ckO0czNqMP5gW
+wtmNYFjU6IGLieoxhtYSWnS4E1UrLuOgK+vGxtfxTD6dhJ+doIEpBNd+KQls1UQOn3EWD2LfzUL
oFMokQMLsdnWCqMx8eIrv4INBij3NbO/Taa+h6Yx7B/VQVjb1jw5yw372CQxYSHqMpb86H+LcuQH
cgyYYxoCeMwtQ5McSI9TbAaIyY3FRdTNDWPlmEC8trM6iUnsehvBbujEoJXdCBXh81ZDw+ay9yXi
o22sE9i7DtyOj6lrG5/tvQ4JhcCuqwHChxV9yP+DBMiDsr7GRqzw7b+cIfn8Jb71JeEa2mXyApvY
N2/hFFuCdrb8mrcd2Ob+Aomn7ityVFCACMANgloo4rLKDu3yIulFz70F0wA9134jpuH6aKW6zWUO
EWIymfwFv8iqpRTAYX12kiqNFF8YXXxrbhv+S1OX5CN4pwYA+KKdE5LECMCHAN+KB4MJHZfckZ99
TqI6MN3dStUOu6UD7r63Vwat79cQHdH4GclYpX86CEXAK2VBWhjpiNFDOzjYvKcVl3eopfwIp9kR
C+vosM8VjqmNiXFUS3JIYbUMLkcarZin1MkMTqulkWA50rVJBue6tCHAkrN2uUb2uqkZrxLBk2MT
QCmSVaz5uIXDaq0nVUaagDiYhRlvedezQIDzEE9Orx6EBjXUhW/EzA+WYeLZEJ4NbQP6dVLpbrca
Tt4R+BlS0GMZOiqPTa07RsA2SXxpczI3WjWbYopPH0ph9inQIgup/tgbaoLsIhsu0TOBKyvH2FA5
Jxt8NN1xhWnzf6toCbHHRN7wkGiVJAxChLysSLAvtXWRgYwELYf496YNoY7DLXOrS5nFtt5JgUY/
V2R6XXTgali5Av6RHFVIH6gju0JVN65TG+eHCasC0TsSu+UMIXMzR96bKZj1uZtGpi/WdxL7Yc2I
samLRddAkAxfB4Ck3loSZgZTs7o/BGnc262CeeeBD+FpWt4CHTzoHtfHebP1k+xg4fClVuDEXeED
Nm1PsvAXhu8kBFw+EXxO0fQkNaU0CuqkA8gYZfSA6j5HsSOGtmGAcWEo7aTlaY98CpMiplGWiLc2
9ZsRjrynwXTdCH9H3aS1C/tzgQamjYxx2N56CqHhjnbfIj8WOBuOJKEIoRipehylMVw7BN11UYUm
wAVx7LumfzPoUaOfsoE0K4Xh5kpQRYS0CltD/zQHC/+JQp4NiFfxL7V2Hx3zcSZQi/PussYgKRI7
QzQ3ixUQlPBT1cwbReX7edvkQLUxzaC9zZrE7x74nETJ39xVN8Xdpab1AdE/efKrY72YMNEPF4nk
PQ1jDjtuKyeSuDDViM/TafKSc1Hdhtn7X+n4DaG/bz0RQeNpaJrU9sLUYCFviDkwWb2HSKjgLKYe
WiWEQpKk8wEfYKKDd0wpVmA0PE/UdZvMPL/z+lXLoWgPgck0xM8TTCcdtXsJ9FLIHSNLlQSrC7KY
GvA8Oo6x6t0GumitcmhQTAcQwUr7692X5Bl1e2GVi0eBRzBLoU7nL+ztf0BicHuFvHm187lbfUiW
htsfNaQiDM8LV5fBJsxigUpO8MsZZZBBfhNFCYGmw1HX3GZNsjTWVoMvSqN+baWnhP46LIDKdyxr
gVeDBCWkiq+cypUpJDH02gzYRleADofSt69ZnDSg92E6eYg5Rtz594PPFfmrxK/ArLLvBt1WPzRI
5GMAR1fkuMH1BUmLKylUXMUcTGcDYWVfH4G/xHNqgqeue0ymnTzhM0AUI73OLcIdNlPXj9DM2Ls9
uE0E0H/ecePyjEr2fzvNu/Ex0skby8Eo43tKDn2WP6n4BkSKvbbvr0yM0PB4JhCe00us29bUG13I
bNOR8ZJm22OxKZ24ktSujgr+GRoEyFqkNycs7h5f21rSbAxBgEn2djehdVwQHeP9Gu3Tic2+9eoc
0XEd6cLkPNw9we5I6V7V3HdiwvTExrJARahPVCbqrk4he4PjHkhicYpz7XdhM5sY/BdLrVkRloIv
eESc7S7ipDAAnnbXRRiCiNyAA/qx5HcRD0iBHnsyINN111Pt4M6V7cECXw5QiBj7vC5zdFPZ3flx
E1pIZLxl8xpsXiOortaGDDEnpcwM2zTqYFyQTWn8PIeRv2HIAiMk82tXkv29v07uNnNUOAFmHNca
3lMslWifdhmezuziQpUm3AMmhFCW3+W4ooT6KOFEjqds1+/3vw1hbIxY3G+Qm5FtANBBRjsN8Vl6
pBAI7WU3V1CpVhvgIcEGT1XSVAq16GBz+PogGnRdFy8WsPcd3fv6br9ASXNBepgD7meO8InnCLNQ
G9NYrBXeymPJoeCIRtbaD/5jJPb3lds7i6LnIViZ5hKgeEOkL/U8TeKL+KuerYxgiOBzUn7MvY1a
uSzT+Bq6xdaycrYC8Qj1IDqkoeYdyLDTXXEBNhKFNeozlgaPk1/+TyzAHEUvGhu06LNaEdQufyvL
vvHIOoXc2GNyulWoSdq7Bq9jhiwU2mbI+OsoFZy4kHm0aZRQy0xys78364h4eXJcKKLcw3en0YJ5
R8iu3hg2MLqBpTQ0aTosUtb6LPQgIaqHArLN1rEpw1IKRVQqWbojmfrYrAnaQn9YqxqC+RxBk4Bv
RX2hfisjP5i4mGh6YZXGGSYXx9Uln0QaLAvovdOOE3e48ypPZU4ATmTOLVvk1NtVYwDYunvUS4uY
uVDbk0WZZM1Tbv4Ui26T/EV++HhVcZWiHFj2s+19nrTTrpOmAMN2bWll5+yPNCoG7cKkNUzBBMBw
ovkkpwCS+WQKlPch4pZf3GJte5TNgpviJlXpT/aV7P7GXfZsBewUfqTWJLMrtiKqhPhBEEdtwgFJ
9+ESqCNz6cKDh4+mI6rbycpciQ6eLkC4O5f5ELGvMPfxY0aA4FA44WvOe/OqCeZCve37hzqjv/07
XpLx0XmIputtlRvxbGqbUz1G/cDao6NUTtBogtbAaNNH2hQ4pwTIzgNWZy5cSvh9KKcw2wOGLXgr
UjVohJC4vAs06uBOEOZYmXcXu0gaJnG65rUqh31xrcZQ/++dv0KNyFhvJH5VeT06Je+2KFhD4VMy
fBrKuzQXRY9IGkYaCatujt4kbfXnLKCXq9vNkMxqKWle1XdPDV/TTSpKeAEuM5d1D6LdyIlWU/d/
uVyJfPzihacrs66mk7SC2skCCIivRfR1hQSsZgeUVXxGEgycyTJ+rI05qDEWNCGil8FGbth09O6/
1Wqh0ihmPaGHtS5Ifpgocis5tbVJR8qL/vNVXEKnfBurMOg0kPc8/LAegDzoyg4yHfs+bTJuXF6b
wbu2iAKMhA+pRCRBRunUpvBALW6OHXhCuDqyfObU2AoiAFGonRu+4FKfN30B9Q2+i3k/z5eTc3Pt
bLA2Z+tSnYoFkiw0LmiRBoKP7lKEBd0IDgIWjazw0eoAM3G6Uc8QPOuyiAsIHYKeG0KNlOJYTdBV
10IIODuUTjq9IFiy+HXzFcHxrd+L1g1/6gWe+kditi/X9qwtG7R6k9M0w+I2X4yz2nq0Dg9RsggB
r47t0KBeUsP21AgMckF0qNhrMLdqHnc2WKhlzECW/XHSsVHXqPP7f2mxZCiMRGYvJnJ+3NeBdYqA
Q/SQSlEQ7HiXVEz18LP5Z20gww5KGV4sRhS/Phn3g8fLzlOR6oLoRooCbul8QVXv6kNBcELm1Lfi
EUB8El4AihhUoKP4tBFtAvIFfXPPF69SqsaGEsdtOzILDgWe3OwzBsCyUDeeUpRsRz9R7ky1Hz90
EWNBod64FM9BtkhH+bEY4nfZc6Adm9Mf2mgi7Jvp+dkXheCIRh3rOozTu1MxareamjSiN1Xr9EtM
Me734Qkmw481mAj/e5+mGL5vd233DmGY4dmeI1qvEoFwHiRo/Uit7UuqgSS2mrN+KIVjpzkiw0A2
KHvl6SBCh18X500h0ASwgdGjtM5tjLSvUNdreaSTfQYnFaflmEVNSAfHpOBSB7zNTwEMe2NqjwBc
KaM1ibdv3zWzxaO22byyMnFuEmwotw7VPl7d/Fz4oiJlK7ZY0tdXFzUSP3w8jA/qmnzIsaSWPOpr
ixdLMf7ks4zHnV7G0nBxqrdgLQ8V2f9YW5YDLHTDnhUUJiPaBheCnY5K8d2HVEvTB+vOJxyDSiId
xsLVTz8h4P9Lu/bX4RwaYiKNcTFZF2rK8z4+k91nXa8ckYY3ljFjLFasi0UlJqIHJvfd4FtYkbwE
WZkOYVXGHZkKkSZ51MuiPAE9b0vAnb20m8QqqPtlCnRDHFLmW6z83XiKhhxKrUK4VLny94F+5st/
7qmSbaHNe7vdY3c8OmSEDI7PbpgnEtSa4x/Kf36kFaEXOsnbB3aKL73i/lyJdkO4E5PqJ9dh3qWO
tmeaezLksvLf2s4PYp02JEID9skJKwA2+GS8oTJD89KwTgCUF0GXNLyIFmUk2oTbzso+wkXnOLG0
rus2lTe2XQKgcStwYBt6bpxQOsO2HuJaQDW0d0W7aFQQ4/EjB+PFGo3AI12DtGwRHbbo5ajpY6FX
Q6HkBz3hS3Et4LSTxWuQpe35vfG+oh0wfNNnoOIht/o4HjP63WWDuTSYpmViqmL4mOJ0SgyK5G5T
xFivkcN4qaIHeiutsGT2Y6DsapBfktb+yrPPczntZCFfUYmZ+L0eMSKJp+8GsKfyGxo/I7IjEQDZ
r7b9ewlG+BHkKHveiJKIq6OkTH4KAJ7TAqd7PxyJ4ZqGNRewwJbr4VqzmeCaZgDnjhnKmtRe6kT8
sX4dMJuGVyQwm2j9edPeeqbH8nB4ZW9ZjVtsAe6iAosQjglCs6KaVsi6MfpW0x2ir3Oz6YWK/0i4
93ssDAT1rDBtUzEV85GXCc6BYUX6o+mGKEWXOA7Nn72uS6M8PwK8Td+dbcP3d11fBxpV7Pzan17w
3Yk789nCpwhrbYyXsqVrd3fqo+iEY4xxcIEGTcnbWxzZEtl2wIs+HCsxtnd7wWLn3yzzyw9vhw3n
vittTeLyUERGyFJ0yPxXnwijPCSIKQziTpSy3UK6XteyN8prYgT5a6KK4Bw4xRV7MOAixyq9ZKcK
c82MTw4FvkoIp10kNjtYcMxUsisG7xOIaUFlyCUUhFqROlVKvfYn+AWNEuVP1J4s6Eu1zA1Id8rG
jeZMMNItjHmdFSfR+eijOHiidhcRoKHGRQYbnYfZINT5LowYeDrBgjyUFV+bk8BA0QbBe30uUusT
+k6noEJpk/m296eBhWh6MLoY7PWZZMF8EKtH82hkyTs+25SvRBhs4VrQ1HuOyo1jIa+1UPJtbHCj
jF0bUqtHm542QUSZMjEKIsMZX9ZBuGDaX81bXcet81x0Ly2zndte/8heMonf9cvW9yRiDDAZHCSR
0TAUTo0XirvTtsIISw8FV8+nYyic3zgX1InHieDns5jWIq64M1sFTzn9PcVkXhGzEp6irzUrzIpB
V5e96VTkb2xEOdGr+hdJj7CqafOcCpBCeO5kv3DeBTHaNCvaotiLaWLx910+4jkXFVBi6fAHi+mC
n6SS/XJF6ncjskXGvWhmxPQ6EprxD4h5y1tfXOu7MRjsexZJKJ/7yeuBejquI6B7P6LMm2ShEDGL
R6HpTdmKvn7K9VRpqCa5qY/6iNV1ua7CPqcMxlXJdO/RlT342JmLreUyJtJoWf2CMUA+89Lzh+qj
m/spdovqKi/xuqr+0tI33FWqrgxfUPhi9081yslXK4ktCVzRoqsY8PnzUVF5rlP4ViDHZkd4glTI
yAWn4wdDc0jOwGT0M2KHDGW6utQtHceW4p7WXFCl7GcQxANe17H0TcbGPplV62DmFQQl/c5EvHnk
8RodGEPJTFOEcd3nXknCubYFBJcvHRSqRb57C6RgRK78R35d5PvIMqO+5ekVduY/XB1fdmykbf2O
0EYkOPeVMUI6r/HATecFWrLgMl94XDYGEKih4ZpA5VBKjANFqU4CdDlNaFBGb0vPEau5Pn6Mhtxt
0f68gVL1nxof8U1kpLq8og7s4de8NFto1mv33nKpMRETcfhtof5TyLH8NVf3oT05Ce7UWjUEuhp8
rBL1trMBU4LJf78HjgGpzJDtSZYEArpwBoSqbP8votMZ2Os4kSuRPxGbqeDpl8A0o1psv5B7M+/k
Il+FzilO7b10RTrwQrUv4iXpWyztP5/RXR85/rcl8l7hyE1FmPePMtg8lruZQRvLMaXDU7CAkeww
wk+lEwl+BWejsRsjAEKr2uZal8XV1kvZFpvBzN0kwz/Hx2HgCB3yFjHrXLhnD9HYDakHMJn12zg9
n4p8XfUQYcHeDbmJkvbvar2kNjVpgwQtg0vVw8pzYHu0EzQalVgyioKDeeMnfYi9eJvetZXKmCu1
+AVBZvwuol11YK9tBSvjA6Ybd7HkqIP+N7nu+JAd2wa7vVWFhYebMX0SEImGEpHd7J8kjLl9jbFn
+Z8sH/Cjp9u6dzFa9pECuCK9jCVSr9V+aDH8wwgpNr+ES9YyBSow+JEtx4M7yEDkMnDpHgZE+8FI
go+jkmP7161DlT1NvkoiPxkvSHuGFyWYJJOsMdVaLHDV2Il2MIYpaO/LxzyuMR+0coLBEAKFNAll
fE1mzALb0mDCaEC9z0JQtemHScNRMVVwhO81yBUxO324/Hjia1y/CTUUhn2L2EcN4aUI/OU4n/F8
d/ByZPV6aEP4g/CbZFI37+Mv99v8WVh9Do+sg4RT4EjKQ+iUO/4L9MPhJzKwPYo3N0iGQvBZvCkT
e4k2hUATQafIntk+timmK/h2VLk5Zg8Jg0JynVsDZCopTt+H/Jnd6FN5nhsq17GkqQzqiEJ1vMJ+
nRt75SlfSIOC7FMx/vzfVmWlSbX7I1FwShq/o+cF/ySO1P/DJglrbYMrjTBFwZO5f0/UvH1b2nz/
K5ae6lotjQ3prpl7mO/8Bhr507HNIcPo979+cKntQZaakOTt8kKXNOqOECjTlMdHcVRepfecOfOO
sx6kaYlvObHge/WPAPmZtqNptZ3QQLnORbZRZckdTBtK0gcDQo+VGAc34RyOTF62y6Y4AVvFUNXH
qj4XwNZ71KtEZCPHLtVJPuTOtax3rcydfkfpalkGhLcIpSvTS9xFE9umBDZrU+CArzntdfE5YnBu
ctjR58lKijBk9aDdqQILdGJ7JtWr8fBzqELje0IJkogs4+OZ2uvQ/TAwN7O69m26cxJSSFieq1Oy
sA+ZZhZzwZ+navoaCnimtB1K5BJGVILts6p/1lVwMI+0TIo7As5qlod9CuKgDYU6iPlwlZMsOb8+
D82uRu549zEDHfDDq4UoTtumjWgTSA6OzWblyauaveks1gDGt18AmiLliFRtk/wCvIPWnXmdoOxL
eytrDB+G60+wGj33SiWBhUYqctF+UApX9izz2aXRmN5n3G/6wDKQGKnbtLZTt/BN+tvmRSGa5RMO
C15BfMyVJzGKy+QDXTgAskP8loyU2sS4uiw4muw2TpwAMqqNcmJkQHhQ4wOg5nXD9Q7NWQwqymof
EVJWQhWsM4P8B+TpLqCclioKtN1pUSk1u62kgS2HdppxuoNC9nqj8p/uMuTSAvIS814eHSJNkoGr
zxipppq8g4Tii8CsWUsLCF/qlAKgj9ngH9OFUHcdlzlNWLXjTmIeiAxOeaP2fPp2cqibWF+BGbKO
UVIge6iOKVvhxZXp/+bQGpXdigL5WJafu7MKSEizDJ9rtHT4VIWCO6EbpkqcoQIQ/7XhDj3rwSQK
P+bIuKsSAcq5+i/bXYMxEi5LAKt6ocby0mChNhzBltPetbDLm0szetMb9jnc6txqfinRz3GbyvPi
QuokSDC85Ykf0aIvngsMzGnCW3T99Difv7N8/dSXRiT0Ld1bNIZpQMyfrkY2lao/dWcKaUorZiPM
Ipd0Vcs34wrPTk+mm5KC6XCMBQouNPlIqGel25TRXApoA443jvVJC6eVDd9Pl10NN/OQKEWV6Fi9
t0HupWIMW+1tHcbDdr9Hk5ivoOkfDKbCwiayPuHPRowH9kxOsnKLmIUzG3nDKFexxYXR5SDTRrrK
uptvFfG4k/o9YyzMvqKrBEHBwNa8lhoXPP2zyJ6ZOpucWy1vEvw32ohYfqn4IY/wElxLCUkKroLt
1ecxWppme74SOxsiSbnPVIxQbKriiiut85fCGJRHbdWUX4nOFpPgMYA/OZM1mnOe1bDsHEA+aWxu
OcPlMBEwMg7p548Syah3y+Cyr1S0uN9z1izy5FhR8VClAXuBHu4vfoLf0SADlQhp2PEY4HdfmR0P
o1W2RaRt5vXb8Sov9OLnuExsH4H09iTc+2CUbIpBnXmtQSdI3AAa7kb6jX14eRxw8zcw6FZD6I9K
aXH7gg/vdDnv0CrTiAtqfGwHjjN2Esi19IgQ50GC2CFJaLSGerNBUb8iYal9Q3BZ40FQHTNOh8/l
ZEY6pzeMTrzln0dG3OLoHKwJOw3IfzkF5Z/G8aLkoSoknOaJDtuJ81EzeomwomDtWslEsYfsdOvj
EtNNhwI02MrEx7cE0qBtITCOZtKbOImbyhUzrglD2GxqcQBwHbOPHzXazLLwugr6yhXsvMun9uvc
61v4KF6ZEvfsULFwtB14QvWW36yHa9K7wwtA728hsCUYrSHHuZDFps3FXawA/r5Nl4WxlamziYcf
tQegsZI/nTGNNTrWkyjZ7LaiJHrPDQWmbPbduwNBl5aPJFIltqOnN2IGbHnuwt9ECoao7LE2CZrz
EiTTFAPOElRkHN9Z87NM8Vr5hJ1Yxm8ZDpELXgubYv4AcOWmudJA72vLHohdt286ovtqzzDxgEVw
fpxIf4jp5eyOMcWVhGLDVWYkmBSGxDUx1zZpTGCzXXhXP1qzMXeVxCZN27eebhXTTZP4xej4NTEW
jeMk6bh3GRSYTMRkTeiO/xdc6BssXOVyxirfXpOniXD2LOE0yirP1tKdsSLqwHIoZme0dAxptCOP
ItMlxD+/hsEYrx1KvNwIr5Wwk7lNiG6xchpoB0xirZfFp9xvOmwa1d13+Wzc1vIBTiW7Z3AP6v57
rlzEX38Rda3gMYQ1A0qajFPF4BS3nqHVjGVL6SFona8Cdhsi6EKhNSXF9O3Zy3uwSLI/piQDhGFr
AI8KN0+WbpTxKYheaIPNTDgbalmeih64vU2XWoI5JWvt8kON8kSrwiMJ9k/77jf/kuY/nJwmWZN8
kQ31sF11IXN6t3isXcTl2pKk4jsMcDy9uIx2+djNrgYGm2lvXjO/dmPvItli2V8HdmlEGE/0U7nP
GIFBXO66QNTS96L8ydeYoaTVSh//MWVWhocNVTGv96IN1cDBaGKnQk7vvLGJvz0l4OcXAPvB8DN3
1zrTZ+DbrUff1N7OqlGHBiS210ZAMW7pMWTZ6Hg7sb/Rn5kCkCs9FzXubyD/15fjMQvvgq70I8EP
YuMptFLKVmvUSuo2zcKCQI8ysDRP1lZtH93asxQxXK7ANbwAEHRit/l1bis3WOBqZBlORpshzZRQ
x9tBYoW559rRmI3O/bLiDSO+ERMZjbCAuKIuLBL0tjLXKTmzJbfA1LPTcSLYp6iaJJEYW5jJpncS
6PDYpJD9gsGszbJSvCRFXPr4pC73szHRPPSbSh0a0a4/SquG4EiAG/DslY52OaQ8ns0qPP9ITUQo
oCWdRNCjcPqRRWfB+m0m4CIbHqUK098E+FJbjOlrC7Xwg96w+4jsGUgdlmSK4h+A6sRzy6AorG9Y
jRyRleTUMM7dXPLTHtgNPK1cQaGpJ3MuuNhDqN09R8avj+KolU6Wz5/Cy5ANweJIX6YjmZgK2d5m
pVLJbwNws4TjSOnr8tgzKLa540HlKQ4k2QGJFh7P9WbtjChqKNrtnMrPubXy7e5SHEBAmFan8oQL
oW9aRJ7QmOaHWoW3Ldw2+3R14KQqJ6c9ctKsktsaJml+73njR5ds8G8350BDxN91OiAWume1laP0
Ks2+CiCnJP3Uq1wVpmOb3tYMFZNDkIkUrQaojiBs0fYS6ZZYZ9slMYFdCFDsC+Azi9qLO/Ed4Pt7
6+9dQ6H3Z+ZBArSzHiGardRrE2gSE1uiEHwTiQ0j4FlM3Z3WBrvi/ixXwOteyABTVnfmwK3AWXOX
Up38iNHb+raoFUTylBhUeCf5DTKNZ0UvA9c5hFChERPg0b1sJ0qLsalHLSyym+jTBCzHNy01yPOR
1SuO1fEiVtURVIaMiKJqSWLpSD5Pam6K0EflyaPSpJ7OQA9qJJhiFTLqeIYS44DMNxwVNcoH0Ixb
SEKD9461IiZWd8lwyuypDknKVnJWdf+7Q4+upfZCixYti5QRPvjejHTCj9Tb4eCt54HVWDQYxiPO
BpRvcJ8wgvnNN6BSVaqaOr2QY/93Vt5xqz3GpqJZ3ZgZRv4pZIzdfAgv8ic9NZnXB5/Cn3ILr1PH
NBiosGyucMD1d3SDDSpbWmYYlIUYxYkzrZr+hJPlmYBd7y8zhE4Un5AILmt7c9IfsNcVrimvmAXt
c806JeyhzKRu8boKAkBh8oKrdKjRx6H82a9jJy2h7ARvejhBjorbh+kJTweygB3JmCaGBP1TW231
hXV6blNczjHHSnGb2I/KODwrquVwVs3Yo0TVIDcmj9/O/Cgq6nJtbXyon+qEXdADv3W3PRfrFOTu
psfgh8DHUsNiSZU5oLNBmbj5pLPjNOatHOpnZ9BJFaPswbbbwrV86nL0Lfg6zRV6Av3//sxh2I+s
VcBeFEzmf3Q+nC5UQOR7E80v66AfS4ZPI90gPv4IX/JRgDqsyuGhjjZPdioexmcoIGp3yM5wEVUt
iGX/PXOLmzVTcUS9qOFIJqxKdTzmfRt/nAe8CSXVViuZFBxUMagPFD+kkvUbujniCbmLkTSFlXf+
hyjzNOEQqhZTdtlaSY0GzMXG8428/0Z5XeTHxlrhJFVaCU2pHqR+xNYDLEW+F9L43Il3zO/mhWtc
fSiu1SnABV4PZfWY+AzPtKksLt65pyCoTmL1rc7X5Hs15uISPxKJAsxfPLGUaE+4334D3lDedevL
3qhiasga7d5t0EGImjxmP0fWKtV2HJjORSyScPebQIuDgvYcL4xu7pZjt0ZZohjLVu6D2jb3PML1
XxoXZwz5DJIGCtdp4fOJFaq/B3k5+RgoB3RBKZ8hhdBvmTttXGu61RreOZEojiAz5XkDJq/ijd8s
N2D8EZqkejrcOFDcGRRs3rG+k2CckRE9D8oRtI+0r2gQUxN4lDoY6VJjrj28Gcx6l1Gorr5/NP1z
Egy/gRmlsqaRZmISuaI1YNU2B3hmRhNyUF3K3Yf2nAQTPAFJOyxenL8qxQ55SfrVaJrX+mlEml4d
Ox/RSjjPltg9OFrAEsGL7K4y+LNgrvZzVisztryaV9auZCq+MnDDk8iKeaU7ZpRRV2eMxuEzmZtG
p0NCbRE7FJmEFQG5gb4M/oUwYLezfmXeM/JFXcfucxfBbsQjW5obGAfWPtTXvrjzzRSxHjPM13Lg
9Kc/2gGQ4+jKZVde5EwD4Cz8dCXsZRorP+s3kRAhAdcnZkpDXHKfWSj4L36eiaEmONnDhzhR384Y
ieTsrnDEwd5Meqzd4/uylHAf2bAGsz4uQMnG4ywrHj28UyJyQKZj8SF1aG4Vd9qvLd6QFUwX43GW
zHv1vgjTx8ORpbllkl5C5M5Ms6ENl6lDjLkKHlzh4TPX99nT/4hr7bs430sPcIiogy5ZFOuyYdbX
TUvQrPVZfe6uJwIFIq79c9Tw+g63FiuM2I/nprgzy30qTAh6qKybeSl+gyEXLrZ48UNboEBSUCGD
5E+EJZt7e92BJo3AKOaI0HIlj1asleqfzqh4orvrpuZxfU22hEx9AawqJGU6p1TU80JALn+ce4gS
900Vg8MUReHpxcGLMlrsnR0iIUO7ECp62GbxSKapioXEWE3xw14bqNIglTu6nC31im4Dzx2aMofD
EKCm6mZA5SBZ3hcuYtKsN0gmkCjAMnOUiEuc43HOJmSnMpbgdyh+GwcU9c+NYLT4j0k8ytN3VdXf
Czka2NAl9QZ91tpTRrAYMXeZNA9na2Z/IKdF14dHe2Mh5yoZyuxnWNwjCx/yt5+8zx5kb18Q4fLD
oHXURrhU9y4RelMnriynaB4fjN0EVHIUNU5ssdGJF7Jy1dkUL1/Gzxckm1SL6wVD7ZtWD+pktuCB
vaPJAT8FySXHDD5RpACH5xmUIWkhsEeQOfWRgNAqbPMxzxsHdnbdvVQe5ydR0NXcbXOkcXBm//mD
xs1d/MeeZNiy2xKB1C8yyqqaPOs57k2iP2ePlDr7zwDDZ1STUmP7xCvrAxSRwZoOV9Ni9SFCTMLM
J99CULBtlPRJxpOxA/uGT91C0+eg7ci0dESHIjGAiXXDjBU4wMFUHuKk6VRkQKM6W3WvYStjyo3t
GCk1ZrBR2UfAq4yeRGUztDtt73BtoqTUTWM5CFYyo4BOOY0IzUEq92LHJwd6Lpu04xOojdHS1er0
b6CjYOTY+DfFH6gqe7OUktbgGVqYTT7lpycLsKLd1a0vhWImbYYM4IqSG63L6GPza7x1bexCydSh
zZXuRYFTxj0nL6cEBTd1iIPCWhcyyfbHKmk1lqOiyiTEbtYVIowOAU6F5rdihr1g88O1EsBwvNTO
AjvrNhsr6NC/Q9yY3hpbjsk3VgfjrB9Ou/Up0MF2/VNvvv5UqLv2WheGQAAMsanWQs6nhnR1lHP9
UPwlS7FZJOUOpDiPsaqoyZ+/MlfWd6krZDfhSK7G6KPOTlWm/3kjEh+k6rn2CQ5b8xZRikL2Zd75
9JucFAFb5JyrwBrLr8zqHvj4nWYKIqk5yDAXvgzoLb0j1dtdrn6asWUFdNcWNeMl+rireGrQRT/N
wB19d2myEMvB0fp0Z/91AqSLJ2H6+iuzTVGlXCdroPtuqqiryRVIdqXK0kfeTj8Bjizyzb6pK0AY
3gd83twY6bY1e0c/mVtT4PljIDqh2u4xKCMg+UuGLEgGs7pgVfoKaYvQKAaRjRF77EDp8sggwwBo
SWTVcuTcrE3SvhZu/dPHr0tx6fYlJup+a8FMBHo0oW0FAevXYZ82bWSus/vp6yc29cpxhZd0nI65
JjjG0/DM/A0BHMSrgXcnQxdIvEBA3SCACEBgFaLeBELgnsnQkwOJmlgfmBPM9lX4rgFOQVFEZuTR
Rj5xrqx/7UHo4McWZ0abh09GTnJPchaGt4humaencfHrHiiCtUBT/oVQniEUgKp2hJNMKPsATHCD
/wxC5pfw8pHU8M1ak76ej9dx35v6gtFff6tUlW+S/E7i+02s4izGdq24o7hGrrS2IobpJ/Fqt051
kJ8IiAcCRNJ14a71oWB6EpjC3nNOkmcEFeDMR2UbkyL2lbNkNonDA9d/JGYY+gQguRbeMJn1hyj9
4dYx8VB2GtuGBejjcQ0b0bWZpsVVvgfjLUquNEFMu63Za5rx1YseqvwLU3XZ33Eozzh17uDgaFE1
4ITFE4YVzVgYvCLSDkkXB6UQVqimJCRv/IcQhRG02dauCd6ztsBRJRo6uaHDVlTJu2oOEvFa3x8k
b0tw/cv55wS3ZCDLdO9x66BzQfY03XvZo6q/PnTvS8Xe0z19SRdj2G8Jcb/NsJ+43c4DGDpE4AlR
vaII4lclzHCZ2eDiQ0wUyiqsBKfUqAy1RBHZ3rhN4r6fvaYS3O7ofmSR6GqlNKPhrOdoanx6iXGc
fFutDr4ZHy/W310O6vnQObAHPHKFUY3+tCILDReIgcgb8deIplGn2XSOwKKXKhb1hrmsHrxEUSig
bSG+oBs4Jm+tAqSEMgLFgXE85rmyZfwGz3HqM6ZITdY5Xq7rSmIi4g5pNX6jM43azQGVjud9Oxgn
tni1B1QOBBnkTlanesV9gzkR4YCjFjpDEPXzDZ1T9pWt23h0eK2s961M5lIA6t/7oHO6Nn0zNfd6
5an9mMJVgwqaJhXQ5sJkUzv/0fdPO25yyWr/5G3/aEQwviMKtXIDKSTBcOHyg4K1lpiyy9LQOcPE
KQOIgfDgcIutA9b/hkc9sAJ+Bmq5xf5/v4si95oI4fxtnWIkuTcX6EUDwMsAtWO+BmrRRNven4Fq
K75fC+A0EWKKq3/qEtn45aU9d/fapcOX5/kChsKT6z2kTICoGT4VOEByGOCWLoPSNilB6Zc22oTV
oV5fC0qgOtFUobBdoIRLuJcxjjQIeRClFkKyzbe7st+pFeOu731HhqnVuQ1uMqufMMmMI0zB0AI4
mVXzGAfI5+U98/BFIRTeW5nOuSwdYF2OC05zzzRTWyX12JYpuHLaLC8emVf5cpQCk1ayYSBxcQuA
fotIcMKMd0iA3BljryKL1USp9cqHHGkqVz51y6+tn85W4jSyodw/NrEir6++jJxW0HK2JEckG/a6
IamsN/uKLLguX/y+RY1NFiTYwn4jTHd0edds6u+2GH9CWPyJbmPbQMtHypqEdBxn3qAULWTYLHgd
TY6fCOWAy5igXbQ3JS5f1eJXUPDS7uHhPz9LTavmL8JVYJUUe5I9xvucKrdN1raOrheJiu8hcFhO
9AmpirRkhwplqULIBbImAypJ9vMd+6H5sccDhPno20srYVYzeSO2qzwQRide7HM3OBUn/svEbb68
TSPBmgDMYv0k3+ngSunVnuhDywDI5hXWWhCOywIMQanhK32zL1brssH4QmohSizkarnrbqb4FU3L
VNKSY4LGKySddtXfDCiUKF7SfkTQX2qEXu2kmIHUE9ESIwiAJRqVHT8o75q2lI0piHXQEarIDm5C
TzVvZgRbb4K93OwdcJm7XtfjnnkTvnGxHOhZGJU0gSgifdIlCkN6boywpPs7zWwKS4EzLCPjHN1X
3ij4l5Qgku08hUbklBGgAhkw6phgRWIIlVMOQNGTeL2BpSjrWRKHCH3u2zKXm6j50VWW/lp0QZjP
bM6X5TcFVq3maaaqV1IlCi6nDKmqMahlNcr1kvrxZLxeYnuRyWG1uYPuS1hETulVG3bkjRnznzSZ
bDChADxmlk9QTxIUr6yrmBL49vriY9tDgk+8dpJIWrws5P23JCq+LvieYI32PA1Lng8TvZO6K+IZ
neGhitPgvE8fheNFwKlUHZbEBkxhMDG7IsZm9K2C2v3jX3VlEdvyC9SVSJKbteJUc7+1NUkjZ7KI
PY+C/wieLG524pwdXGraKQj6hA0bgdIfSeovW/mx2hSV6kLQxjDx5z33LkIuxbGHsv/VRIyPL5vR
gKtfXLjKURxkkutxY8JKeKr2pRP8DWIwQjqrcvbCGc92cgeNrJQVE2eFEVmBgX/0HrAzdHDPDzXp
CKc3uIcm4j5lu4UfmLZUtFg3L/LG27UAL2kuXnCXA/OvP2wZL6WWk2wo1C8MEXGelh8+AF8VV/5C
OkwuVW++sG0TWpre+0KRw0nwiagH8NybB5svOXcO5JX2we3GeAb0S9VY2B/yF+oiO284MFTKMsBQ
XFPGA3G+YPBtay5jKwzAB8HE/ST75lA7l6/At5jwA42BVZZXQJqkpZVGyx+8/ybTNipAq7b29tCj
UYOV9qufNPn8ZaeLS920nmSxFpdTox3biXLe/6O/AZChwdBzLakmFRqumSTc/aqieO6LFP52rpNb
Uv5W50QFIC/9hI2BeVCDrOMab6E6VASBqNqkLXmOijRGM27m/RrPmj3bXqvWkxDfgjOp5SxzNSG4
UOhDGmppLZQpZQLi0BAtaGs7VxGbLrXUoU+byqak1OYfi8qH5809qqVRDjgb5C/HYb04KVhQw18v
z34scW+UFti+tG169i0PGvXQUBMrAeDRXpRobi91oqFJXGqTNJj3lHuYUIaKmUpvx7RM5KJZYBfC
wPKBY8X3oF0Sj3N/b/oOTfTOLnVQvT4vH5dh7MJB4UJa7qWWyYZn9jIFqs7JmlgcxImp4pLwIZsz
5cOm5bKnZ6sSw4DDvJINoDuviei8gAjOCIZWCyPDpUCyM00NKrXUZf75X3gkTfeng4UnzjjIJt4H
1Q/D0bXP5vKSFKVJtSThN3Newwva6aAGCcsNFA34fWIOugNpSKXuKxo8TeCaquJTIOWc4Y+aiLQg
E1kC6LuDwh236QIgFQTS04isVQX/gITTrGIibFGZ+yQclQg49UVvOT4ymDnvTXpX5pKd/ZPC/xXG
kQKv++ZSj+ER7ORen7byu8oQEIZZfCvj3zYFMI6zTJeisBV5xuWrtKpjF1VrFL0hYqIrGQFrWEFu
+2RpCTKG8rydKlcZc5Qv3kKuu0SDqWUXIzs77+8Jc48kmG/UeQkkLXFTE+85SkrtnTU2z8/L9dXn
/sUcnSEDQ8O4GsqrC6OpT/gZywg9hZyop7rojnPEwf1eF8Ijv242pzNlNj4kNbmRyLbUzybAJT0i
FEwukPgyVgWkn+sBWBvHfdyRRqGut41nWLAEBYyGOkzoHbc9DvY1L3FXBzrn79oKSEfUmxt0ULvz
jHbXFMk29VUGSjEYGqG6SQtElm2fVnp5d5gCx51s/ISPGfHHpxVgVwqRtv0OygzV1SqtECUOw6Ni
YaE7H9TKHx5xMgpnyNdyCIa5vwoj2UKWkdVIVmfq4w4Xcf+1ti08uIaJo3vFZfaFtzMEzKzj6NcT
cNV2Rfg6rWOCySRkr9a4aLPwfN9nqUVRtHyZlPstSpNzjeECOJSwV2bA8qc3s2IikBTLSFwrgR2e
eB6pHdjAG2rcoNEZGC3Fl9Q6piawLIr+bfA7bPSjzL8hqBPP5p0BSbR62q34xzLFyvr614y1hRqh
nrh/2iTmLo6XYZQYfg7gRGaXFGSLzULp/o8o24efe+Zhp22+p+CItD5MHfS9n3l4PBVDXTW7FfFH
/0dEzK47dcZckwOvlCf51vqAI2acO+PtAf77YYnVXPfbqnobizC7JlivDzZY1hLZ2tIqutzbcEje
SsuMTpy9nw2a4xWR9w6ayYM9h0LegeF6/1JIeKt/7iCDwjhfVf76WUAhDlcwDR5NJsxrY/O2qP/W
PKFr+thNLMGGyn/zENenttzOZW3QXtQutfdnhOMylUlrnjtaWxI911yPvqHBg3goJtfmWQlGPyiR
dsqDXL8SoLnvUFk1Fbvw1Pl7UTUeRrhJSto0tS1ZitOBUXtEuzALl7nkhyTqepOL7ATgT4sWrcKD
yg51EZBHJouFRSd2xEWcu+x1PitK/cqQ3m/EW6g2WMm/Eh7ArvxciibhzgjG3AzZFKuUqgUr4Pn6
ZV3CHNrbfrD1EThuo1mqxrDhEDObBUYGaBQh7pJx6ETEMVXhllKKpPa4UeO6LQTCvSk7C04upGka
FWObg2uIVQDRECLPBcnGtfY1YGF7fcx3fO+xi9IRUmiRfCtJ5DZQDApVC0SOblI792HaIRsSpPwn
d14eq7aVjaKQ1POTFzx/vZMkajzqQu16wMucwTCtsFDml1eAWXoA/tnRQaMgSpvPMdpe1ktMkUjQ
hIFP+NCK06qw57FkxVwW2FzLkRtfh/byN3T68XNksf9CQuAIBHO5fCBje+XU8vZpfOXkloBeSAzY
3Dmgw+n1RZiosvMnfXdtz1CHSRRuHTz+7ykAupeH7ZtnNsxQoZJ9iMP3tT+9wSjnmARf2Xe+q0hy
C44ebDcCpm6PVbL1H5kmBkRCeJk9a7j9sgcMtERwdni6yWnQfXVcx51jDM8rXwD8FYyreyA/GVSz
Dy8afrSxq946hR8X5PPKGZMYY0HuPQ8QaYAJKLhYLen5sd9O7ULgxmasPmi1jXhkCMYqWtmWUapx
zp/2TXCWyxyxEjOUQNeQUDdDY4FYQ9yA9lr6M1MKMH2o+3nhVgy2nhHw35PGxF+50nF+11WyQxu+
kSZRxjEZ20vyIUM88KH0NdLB7oJIv8hTSvhyCU+1yntA7/INDo4NrhGBERYv3DZXTAAapk1xKCHA
NYhVL5sDIAuqJcOxFHAR3QQBzskgMZwwgzO8pNHuWPNSPwU5xgxMyYzPAaXGrO+ae1FQRdwETer2
lVCrYUOmkOaJ8m9CDx8TdQ8LcWHZYIlIuLjFZsGQBt+nkbVIFR1aEQS62Q3XNuIo0hgNUWuqc869
fT+GDowPFbIktDVrHk5MMhL3W2kHXDm8HCOI6SzZxX6Nz0SVJ80OgkH1Kk2t7NGPofihpM9PU1ux
KsiiVUKPOo8/7ZN/ffRsz5zdc5GC20Jt23GJQMtn7xP2nAaSRiXfrERxbijRpGfdxmEZyzsae1c6
0zzdtonsN1lwD3zAjCI2a5975ETYo1TjIAE2c+jtK9la4+GI01CxizmATGx1S97MnDFNWK1DJuNk
t/4xCkdFA9gcYfqtvY/E6Xav8X876IYOa3ZXd9X9+dmuoIhZU0kS58Eo7aWimV7P82XdzCD/zWbx
35bn1x9Me/NyLByDPU04pcWvXzV1kQD3Q4AI65LVw8IbxzBs6tWK0jumGfCbrcYbdhv+Jyf75r4Z
v5yNXQwNk5W73NlOOAoTN0lqTB/IbF7wEiadUIGU9TmLL/EBw/I+GLjwEJKH+lITGE+yHMB8TWFF
Vx06DZqagL//BEf+2MTEoy9JjhNT5sCxptkN4WaPayrSC2K1e56nVT1po5XaPZmFEx5/s4szj4/p
z9x3Wa3vrLERc2Uoqj6U930OICznBSRAfs+TJvlVuq+jaWCMHA1LZC3hdt8L2ok01LeDvNlRoGU4
/xCSerxZKSpLD//h+IOKT65mJ8k7q+E3WBb3vstLIshZ7ROf5X/VeglZAU2xF/YSq1qBFhhk3g30
QQCfdVy2yL6npJy6rEPMpnPLThvzJibKe4wZz9uxiM0C1F5UGMKQ/8Hp8A9TGEk6XUeJFsxbn5cR
2AuODZCKQhgvTExD+bTDdxXPzawDMd47/WWGVXAoU2+GppMqb2k1SzZUupdZgbHPjCdPt9aPbCnZ
GfBLnUUIGEsh7pOxXMofLfniOevaZcB4KGFC+TAFEiwMX8RcCWQlce80lC5whZt1mqoxyIZbzLIN
6u2A94JvrVMoa+Zo686moDTJwJgWYb1eJhA036TVCdSmN6S1iJHITmvqVOorgprQNa0yTCEj+pg0
8PXdkbg8JO0Pv1TTRg/JEjfZLv+GLZlm2sJJ0BxRkoCjyO06ltZIdPEfclV3sOW1orLu/vionb/h
h9edXFEPbrWo7B6rJ6LjTDOF91/VqRumBZ0RhUJqqZ0EqaO4qiB5odzlg9dMycuemuQBFkAZBGpH
WvyY9/pR7nEYEFnpGln57XE+RT/4HUk/yTiZLyQvsmpezf9OWWL0TBdB+hmpqdBHRllWB0itu0i0
ix47+hrgZqDs/fUeO1uKN/iCpeYKf2x7VoJiSl4jBZaiDUxkmSd2UcYOF6l3+FnbCBwa4y7T1i2t
kRUc6tAgQ/rAcPj5CzJKQuJQ4e44FM/g+MiWkPycL7IWgUZ7lxCvGBo0v+8DJnjoMpwbfaz9+PZZ
BS2Ehn4Sf8qpP79rdwU6GnuC4AL3cm0XAZbh9LXHlwMwhM9NtsAwf1U4MTgBm4yxNLL1ByYSxmYe
Eup0BJgrDfjORraw1uNqI8LG2XXlI7IB7bFw4/uMxaaTk1ujeD0LYfQc+sEdX3PUJQUrJQfgSINX
V9rOHzYY6wk7WcV6YqkEC8P3jK+5XWTBHbF7WGXsQDL7a2AzbDrVUV2n+wAD6ip/SjCIXQhC0iZ9
TFihZtsNlWYtbCImJWNQXkiRZomq9qvXTiPxcxtCb7ZWvnB5Wklnhn7ekCVltuRFMKjk1IFLGQup
c2OUS2oWaiLxLeCOLVXSXde31CXaV9SzSJIiH2QiatQo9cWkR2PgHiJJj5KdhKv7YUgoBqChgD2t
fqtL/zGBWDRgWFc+h3VRecAzeAVMMYTKPPcnG8cwIY+5WWnqovKvXWVb6hyokTMowIk5anttfw9G
HAjQk9k+rd+3HZBuA/tahAwVg2PSww8IP1JWR0SLj2L3V3Sppe88sEQGT/XxvEL0U4EQXBRibcm5
9Uf0wcxJV/qxqnsDt7lcnBY2ziynJryo740+XFxdP/CNiOMgJLL+N4eeNHs1SpTO7EEVsNk2nCUL
pBE81ys/oSzsk0ktvltMIgbRgN/1I2KWyhfAORioquVrOJBICEFWNZ6aTywYdnQ+7q2BYsMOMiv/
SfQ6AdsAsOAP2QnEzxKRx0YMYO9/HRWDm3DL+jlLud1pkZ8BmHS7Zk1gWCqcjZV8J4vAAV10qmwL
7k63JbCAduWbw8cKcF2+XZX+8PmCHm+J6AzItEkh7nFQwGBpJ+rdon8TtUs9gvjVK2PIzF27/+9u
CoQUGooH7P0yswp7ss3uNhnVO1nIjhAePJfXaWAh4CSml5/dvC9c82GG6/pXZ+XYA4SiydGWaMHq
bz9kMvF8qEUnVdywpp/YevO3JEQbFYnF9l54DjPzowmQaQFHHJ7hDT4YnB+TzXQCmHc/F5+K8n0q
x4w2cL3T22UyY++WUQRelUtHEQO1zIYOArYEuHcjTDTmJSD79imwTfwE/E4kiZLw3wIFy+Qe9xuQ
d89gVlqwx28bGjWl9rAnI/jsKdZy6UESz119wnEj0SYdi2CbI4Dctod68EsM5k9NSYRiy2AUn20w
B6UkPnUoMGrxDGP4skqSTftWTRGg5N2tYBUY99R0O8FNa7SGs5mfK13NnS9xMpi75LaBPO2EeEKH
2RoY0R97JoIFsQi4fusTwhtczt6OglFjBLRQNClW00fQlioR373GQzKpN5dHZg15nbZekrwiJI6h
IMa0sFmKv5UMw20LKjf1E0qRyDCgDATgr3cRH/ZtaQQFYdCQqc8WxBPUOhcGB9Wn608c2yHaXL7S
AqYLSPBwvjbw4zGq5xr6wcNHgCdWFMS1rp36mAWnsWzlI6iiNj8uIbOGSvpnV0esiA3PzD8nBbf7
rALc7OHVjBf954TuCnk/qvgU+RTX29yeUAixH9h1emy9nnvCSVyG4j+F3vf+EN92DleMh6UGTz3a
louJoNn0cZwR65XTFC5T6M5Ud7jFgE4CgYVYkyaPpRWXsLkhoCaVEh53+KYwzC58swMKnmh3Py4n
VJ3aAFcIqvoanQa99s+NHLLm5EL8VEnwLGavYtf8earhslfveh9OTLxupw/zW8kbZldiFP64Mood
ecBUMg9MPegPtc5GqHu3T4iR7k39F6PKq10Z9eV4ua19DWUAz5V+ktMPzFJWqWnnAXO0oi8ksC+f
YNxIWWKPIH9HJIjsFRl5RWfBvjQDcyhhOrI2coVZfnjPYSMgAe+nJmWLmH7KdL5kj8lZb0quwjjl
2MCb3q+9ukXppL0bVeZe3U2rhn1fFNBxFPOARTnmJN44QpUlPxTgRd0Gg5Ajs6vdQbiKoqGuf0nC
dP/SHZ4YKPRAsKvWsUSyHX6bzfAaqz+9uWscdIXJ8UIrrXaZTCblLoC+CojbelhK3PgIvFfrxCs/
4OFFQaJRG3vSQtyMFFuGiMt09ybaJMB5PpziVYXbWqgJLxq4xWQ/f2jSicsaWsv6f9jO1T/yZ8Hs
PiGU6DR70cLvmKWAsVceGQiQnW7jBN7t80LPyOXvHkTQxq5szmNks7+c5RXQAMLdVTC4MzMT8Ckz
fS5iKgrOtZVQNheWXxtbKGDN+uP01PPiLcGz2LftEnhDYUOQdcEasIN08ofNGDuy3Dw54OWGmRI5
s47Qr8CHOp5CFZIcB8AqLAFKvlNKBE27EtVGlZeyc+EXucVHYvGDZbHgOcIxa/wWf3QzkhCvdluo
KjgFsmjyVwSnKUhbmvdVqyXrP3LEc4kFL2a5NUBS8NIhLRAGplMxO/1muHGrZN3s+Ns+YIrsmQez
SAwtki7pxZh/LHUmtOemcLjc17+1kuFyHeQUd3ny506dMB5V+UbRahWPRlNg4yEVvzZi9zuABKuD
EannmtujCJ4HhMK61Gy0cAF9g7K/AsovyxAhfd1fzHM+X1QRGeF5loXLjfOWVu5gWvzKfpA8aEFp
FxmPGUeeR/jjWNsR3lMdHD9XjopsgOKTYAsVzNnhYRC83m+QapwRo3rDLZ6+MVgjhuvoywbiKBjT
Yftaa+z+cxF0A/kBOaWL/dF7EYIA/xcA35Ar/d1zbzKQm44svd+8qWY3KzESv3E/qv9UslCN/pUd
hoAO7b2ed6U1ygFCreGe9HpmX1rf4IvLV0Q/MQQxp+bsdgPyXXlcIpuao0GTvUu13SACU3EiNLvL
YOoApY17ZLB0HkYJoV31cpLZap1Aix9asjsTaEzvLg15/GvgS4rNdmvs8zWTVb+2+M/lpvICs8MQ
xlq4jinTWv2Gx943hr/A7AuziB3fF4MKM4C1BUeoJ/5jBsYSRBY4MSoV8dmCW2Tvj6phurNQlnep
vZvQL4coYGbN5Fp+aZqjsDbuSDv7MhIRrjbZ851jxS5/Emn3wH5cfP597h/9Mce8VXsNoGTa5TvP
LvRnUhDVZpZf4eS/VPXZ2DHgXR4XXd2el9ZERg4uyh2qHu9Jc3kZNQKh3yqYptNRB95mP3hcjtsj
z/u+bqZUZKPB/QnfgTY+qZ7hyFZpE+dy319I830sHo8G4Dhb+F2IbnlRY4ZXDz7Jg6A8dEq0gIXj
zPl6urELIanwfiQWKdlHbs9PyiuW409Z7AMB66qdPahVegyYpav0cnXgiU438LLRslwb58TakQux
8z5SJbz9dJJArhx4/jGcLO9be6t5hFY7/hb9ybEMhdiqLYCMMbNegel/inKuXwtABmkaXPMcabC7
uYxpPHWXnKPJN/F9tciXStXytoZ4OQJ5kO6wcLJbh593av8nDoe4NVs3rTgaCQRupdRRcT13Nl4/
lBWVGvD5hYV9QrO66ooZtXF2FAmqrCE08/QToDKszqMSCC6QB6AsNSvZwarYheeCF7RpQooyoNGX
28DZjPxpeqLlYwQIHMx4uYbmlzB2RGVtCwyvCSil9HGZ6UWJXkk0QUAJlre2sVGEboOCepumq/fj
YEj+B+hEk561K8O8p2NdPBaRoMbtHWHv6HZxrhHWC22sghKXqG7vm8+6dGcaTiinz79bMamB02rD
rGnvLsLjM38AHNGSCZYfKjXeS9AA2d6/XyjB4FNWg8DqP7NjerbJyvHDZ05XgiT9d7BtqJ5+yWKI
Pou9A2x416zoJ7HV+bPgxMFP0OukoQHnTuOJsygOuLcxReuhcfWKuRbuFWgPZSY0RTCXKAAl3/fw
j0WoPKKPfhNDFcF7/MlQSTeYG0kMD440RcOgY4JpA+2TYRg3/lA7q2rmKFtRMyVzrM0PuEMopKez
kNlL6yiuUfbyeyPU7T8YYV5zlcCCJdJ30KfCK42chg7wyrv9XaTqPNnW0TuMvx0JjR/cJmaG5cRe
0owDRPEdEaTIibDC4t+IeR3NRCWTXtI1HwBBcaQGmuvuGe8nvdrUp1S+LA0wZXX5jv0tjks+AP6o
csPG980OEiJKToH34is4gDAQDmbJehr1RAWoH0IqWWBThZZodTjzWRlZqt/VwPb1FpQypxqClyUy
ALuChjnMpeDogg9fuOgazmDyu8b3jZel+toFdIQ63bDLiPoKHSjCVU6dUGi6AuNEVFV+56IMgJA7
a7DqVCERThGXidb7qPh3lfvvXfEDWZTFx4X0PIuq2mdZh4VfyeueB4DUj10Wb7eJquNy+eESaa6E
g36kr9IYf3s3qrHyrKZ8ILv6df4Vs+/52m9IqezFmiEhPPbIQAJDGN9eDofNDqHGCcSUbS4AR3Zn
+HWcUm22Y9w+HKl2te5VkiPDdtZZex3qEcsU+seDGjmhfDjn3nCIX0aZQjGYboa+/2AsL2PrCKAD
t2elzEETQLVYfrvLi0WOLlEVk1wCQ0dE2vH5XV/YMiCuC5t+vxLanJdKEgkQz7IMQQcALC2Etfc1
ZLg0qiT62CwkgI429M5CBN6HYcfbOzbUpAY44801fySHssq8cSoXm0xtD8DL1NyiQrJurDTcSReh
DqwFl5FRou2jTyuqk+aHY7RUvlfMHVQvA76UPZVi90JdCzaY3SymWKrB9xqwZIhufneVFKboK6Bk
BAVAvemYtpqem5YhnwqiRzvgAOuCqPTq4qHhraIFhHZj+AORwDbTNbmasNXNN1a51u6ZDk4H1DVE
fTOULHXyM+5hwUeNv3fpEgffVqME0UZg80NsltQsze56CXKXwuSTzBwNj56Q6o6HSXmWDCa7rKqg
enPfTlQFDZS2SBscSHV1LJ4o/UDVvWN8Rq0v0TDhB8qRsdvwjljYe7byJgVvJc2r3jb+LDEgRtfx
GW5TfnRLA5cGyAXaG2gYhKOWOEXKGzWiUOG1yL0IMHjhQC1lh8PNPj5cYyARae+h8WcftXyIy9as
WSs3GYihzA+GxqZaPqYKVb3M0DwUj+iu6/jwssuC4+3OZdAX77c9dho2ZbiTF8dxBxf/yJUdyie7
puc0WlP4xkoBJOYyU/gy0B92TQFb1ZnjgNp77oyi/1U6GghViRKrSUOn4WZzGVoDXuS+myo6Yfme
r6Rpj0+SLCZH/I9GIQzEAoVphC3gOas5ZKm+P7TTf1GB93N/+sDsNiUBwpF8oYrHVww4hjg+fADx
jQB8dC514yOszsjU5Zxkznd9auEAwFveyUqlyPwnvTD0Iaok5k/+4USlsm9yudsYtMezjE5CI7WA
TSz4gQl5MZ6n7/smv2IYABCddVX6R5aFv/e7mXMOthVhH1s8RUFrqb4Pj21gKSCdiBnhsiX4UBZ6
brmTST0rApqDm65VuBv/MCn5yEs24wQFtyq0pxC/+7UA9VoKqNGTdg0soA77eLM1w8PFMm+BxN5H
T6G1km9V+VpdT9ZBiHB+3d6KBjFmgjjlOrpi55MbOjFXzNEKzNc0QWO3pZSTF2IkgUWC28do7Gnk
dtx6kQP/WpAr+hhwcvFRQylZGMqsNww0MpQIZzShOPIlZL3AwihD+FZR/ANK/gmshDS1Mz6P2XOB
H+DPsfIXU59sQShYI5NsDBaH83mXRDNek+dS/fs5jOCb3e2G3a1NjNr9rvM2tWSOsW9o55GEE/mH
xYU28682IYEwPFsKtgx7EB8yNuE8RdFAxp9/JtZxUkIvuL2Ms+J5qntOaEPBpBbCplN5YrnVNVVc
19oO48vf6gPqLZInulLhTwD6TOwoEfQIVz/JXKcbhKw9Xss4XwMUYSRqip6sLoyzLF+FfNwgrU/2
qk02zM1amCEdbDiKySebgPT7msVTMpcs0uu0/vHc2DorbFUN+/S589fvNY5eEr0qMIzUhTgHihWW
jP7+3YBg7IyVx1uQ5HJ3kQjwRpIdn5ox/vcCvenawsP08P6j0j4gf0S85Evgl/1p+wayjLVbDvZA
Co4RTvuktyBJrAS4t7ynug7BmM8SIEB6NtzaZUuLYsW/XQ2mtik6PcHQsNGJRLhD4orkd1v3pFZr
0kCYSJvRoMTDY9jCnktxxe4EEuTprmeR8DIjEvfwGH7bgJCtNw84DO9wSbmeUZ3FYfUVPaeDCjhQ
Zv6Pdp+4on1h8MCVYqD//02tnPoOUDPDy2+o46VkJiCt5/CX0RY8IqsJvWqFMECSLfKp+2kTprPq
GnnRXSgz/uCYDviSXQdkMLrmsefDg1Cepzj9QG70XEHkf9sGKw1wMNenyMYIwojxGQTev0FeZByg
m0dMht41e6xxfrxkVPY2dCw/hh7kQlisHRyVkIjgxWzF8Xj36OvkGEsFpgIDj8+/f41QLm9Mf86h
zmjUaYATg1GHNd++IUfMp3jm5GZ9/CO9Stet8qMwEWU5+D0STh0goTY05/gk/J68QXCfuYEG56wU
YrX/vY0thuhOJMLPrPrYZ5g/ewUOF9Iop13bcnnnHgAMZWA42q27T9LYK1nQsZvWHr3oHJ3WaTqx
DmyyYGV+QKWO0ZnRWCIgv93csDFfQaRVnEZtgw/BurKTOm9d1FNtCqLD9BYmtvbZSVStemyzvAoQ
thbpu+0o6J+2XtixhxIoll60Qd6cMVqA5nHe+Zz+rx6q8tieZadv9nyFjydvimsZuIUyllRABI0l
KmyHB2yAXnJ6M1953Sjo3l/lHmRlr8+IjiFEBOs/XbxIyM9Mtam1xyUhoenF1i61eRW3u6bifh8l
6H3CVM0WfY9CgreftTgT+3Zdbu9zoBd4FMMSzmn6onwZvYxo8TFczLubnHobMcNHgGqH2dwsaKQL
RVmaZgW9PyXYCtokTY8nJhxA74LY68m5M88qEMxm4z0JcoMZP03hiux+FTayo/Tjzp2LFkAcDyAb
ewC14DgHB8BnvC/JQm696YDrxiQbtgcs+sn2vf11mrt43lHPbZh0i2vhh1UvMjfH17+e33YJuFEs
XHI+YsUkKCuZLMjBM9Y6xOkbDUHOF//h2fBvJ/QJHuhLUOgeBXhtu7HgFN5H7gM4ISoY3MGPwTyh
TEYhI8pIxPr+BHkOMqAyHq/4zGSnaxFmDX6Vit2V0qyZ4wwLVePf4mu2DBA0b2L8QOG4zt72T1HJ
WO1lTImAX2le0tsFOFn11xZawrmQrkchVC622phH999fuBioFo3eH329J86rU3uql08feH2r4G9m
0Zd5OtXJ8bsmRb41dkGn/VhzidfJAsfJBwj303jY29IPg7k44CZztWUE57F4+3rvEPkjfpq7u29b
kMKk3Oi02sHjIjnR1AUqkiCTI+kP3OSEAO++sGJV5yO1wxyozY7XgSknzZHQDwWuFqjuOwRP3eGE
kcj7/CnOlUCYqfWVR3mQXB5/WJ8XnvAnO1+m23qdD0/O/IsA9DV0tlJtyat7sfDB4paXGnUPXRgW
b7gFWWNFLemEON1a44oMObqnEPUhcMwiMpx1fPbHZBihLVV/MEvrdliwVKCwSh06NgceVmqhkRa1
g95pC39SA9mnlEd3nBUhWoCM9yczj7UY+pfP7kwxB3JI9mvNHVcumZGnz8VWRP7tuBFl78k/sj3D
J8QFyIDxeqJR9E9iyliQqpTsyAmCovX7KgM6OYdh3RG4ewDAQQrRE60XfssZLqc3Lir2B5ElOahD
TTfk//ymS66jaza1ALm37DozFE+e0ud6eaaWixJiXcM7b0MK0echeEhiWJOYkZXFuVTHjykEBxpU
Is+y6CSyHUuQ68i+euTp2hwPBFSmOsYyce5V2kNtvYOm6kQtINpyaDmpGUEfn2LPCWvv+t2Za8Hf
XyeNmdZoc0SgGAx7RF37F8u3mtkJUhyw3Vz08bpT3DNETcp+IDEAgVDKkfhYqXv8oQuQ+Bw9Sc+H
Ba3nttSP7WK2o/iZF5viS4rZblOJydusALtykToEmLmixJQZWsDQk5fK0WsTwpNAoXtCGz8Sg+9p
cyKb0JmacljYlr89U70lfaqMCnYBkoq8NqAikVfr+u9nqIz8MnKAukjLxPQNnYShT6+9UoWIRKKc
nEUoes1DU03rrYZ59YJP1XkbqwosuKcgrbrHZjT4cJfQacwzTftD2IllsA1pBcOIGmHhKJj8dtGR
kXWzKaxNjCSSFUU/kpmsj6X18KnuauIg4weuLvxFqcZI4OU7JStSBOCYT+LoqVpENjUdLtnSdodh
p7MseU2EAV9ecCLeqMWQTOU3zVZyyVfweYu7N98aMxIMbc9HUp9/oEQ9hbTA+aJA2pQKfJtwwmPd
IX8PDoMNMFn0ROWwAIQrQLgnY+ssTPJ5fr3SMxL40SmN6Qs7O2HarTGrN/s/YeCk4zj/8JOXjDvB
vJwezzBpd0q3GXSJmD6RTCASWoyTOLWM+TREK2JPhdBbiPw4yfzO1IAFDyhKVWU47KvGNRfWo/n/
3pLYlYGXE5Di+G0coflDHITRtA5SCxan9fsjl81hXLcgdQZHdSUP9fmBaRWChVdVD7QTrhG55miX
PEUur2N3eEEJTXtTGoV8rKCy+4VLNpD9NIlJ4o1DH19VdlCxWOtUAh/cQM8Gl7SLywNoLmAi94+w
ULma8HHuBqMRhFVGwKFg23ym9YX5nwpxrH31BrDLLM35PL2sZKZTOBKeBmrb0fBYHgJsKMIwFglh
0Q+r2rFFpDvMQob2+xBkEk57x1PGMio4vih6dvQ0KgIUvu64mZdGKzGVAD+s1EnxymNb+7YHdKug
/l+4NMpSLkIJnzZIlhCTT+ndpFJ5j1G1H33vWXoCuW2Vyxg+D9MvDy4tmsiePD3P9YUqxkEifucq
UcuvAel9E3eFGUrZ3giQGF4mc+H2Mc/KufuBl7/kZ2Fd/M0WUgPTIqGfrzQRuz4gsWwyufWblRaJ
pEbmd6uMvtqfx2EkKSDR+TRhYxoFDnu3odKwHqXzZyINNDj0DdkfL7FVlya3XFmgaVG85z/yydKV
RIQ6OgqaT/iyWRqBmVqpBx8Jrze/7NpEjNUe5EqA7wNxlMAX1GgUQZ0M3+GZ27juw/xkwONqd+mr
GrLH34brBQ7LGlXTkiWZjjTmetuatyt7Y1JSyiamr3wFS2guG9IW/ZP+Y1rqVSYEL7hPkprHv6nQ
Btg2XRuBMkOLvinSzrNe+MLmSVSpVl/ZguFoL/EV5eHjTPWeIWFWzlpMYl3mfwOK0WJ34vgcn4ug
QfsvAwtCjT0n2Vz0+QjmJioX8x4V1GT5esDuoRTGrhFwapftnrwaDZzTONlm6w/h7A4RjyrE8mWF
bH3BvWMoW9EJEOF+Uuc4t1EahJGei0826/+BeWgPHFi2J6fWiDx7w0LKiHTl+6KD7LCQEOXN+7sh
TE/qjl3Y1K1GM7uoRL2F8oSuRnFZ1rtNeWT3BTD6l8V9gvt3gNZ0TBGcMVaMALPAlOyrEL29OuIj
/4axVlsPQkKmpt4g0lr65W0TNLB767MAXO1xeNzKGRCIYL4UQ/G7/VG+WL9T/C+0jHUIlexdRwOo
UlzhTrMUXgCdJ1LTdPuDH0glshF3BL3w9Eo6iG/POHItdBaCyEUTx+K1GzQzx/QjBBDGoDCVEtH/
NzVe/WYZPCBnV1sICuNiS1dINV5zw43zQZ2Iwt2yNS9SRp/E5jK1XiVp6EgO6Nf5UqOUg0vb1ZpI
/eEkwkuxNJA8qzaRJGbbbUHIZIXxocRxF35HjniHOkM1lJwTnDh4ODGnIl8Sdrlg47zbDlPlCC6U
J78Ja9MGGU1zUSg1X1evkhVVd0eXy1hSP0zdfGg7MB2WJtyAjJpUQkKb3Xe8sJLBre5c138oRjUO
9YY/zLar5Fan9gmL3RUE6GSBIMaqxhYgeWuKv2LkZhgJfo6TIti9TRWkgyGDsbZERFTyDYdAfx4b
1Gv0M2W275BHwnOelxhd48BVKrxO83dIKpwBaJbidAcIWoRAZx2f0iVVyb4N7Iu8MvXQ1Csg5D75
uBXuOqu0NyvoxsJ16C+UUmpKDOzG/KNn3e/TTGHMusMmSneT12Miqgvw+Yy/zW6VK9C5VvAuV97m
uJz3EkDXoVgIFM9I1I4QFR4ZSmXj7Bgm/8qr+SYOcyDYtQBtxBmFSkvKzlM9kqGelgCSy+ZpTucO
3cCOKp11d44I19GcOwX/lEkZLopYvo5+DzkWmhuD0h5GHCm9MdjZ+LQeuhkJfAmWWNFuxrYHnAz9
vKHy1ugSe429JPrefx7dvlFP9E0uC7pmb9pHSLx0AMlKyGxWpZJIQch1IveZ5V4Su3Nr2aVJVSTC
oCsIe2qwEhd617mYi5OBni26KJF3ZVDADq14M5mowzUy6tp0ZTOhBNGAlXLKCUB87r8BMwo1qXC5
Qg7RYDrOoRw3HKOdwv/7gxRfjkqp0QJlca7JBT0DbjLLNpr3RaYv/donoz8aLTZv2TxMWEnKC/rr
iHpWZdalo2EPo5W5XVkSKLixCHtOyw1cDsIYs3IxvvuWba+OPdOP62jDHk3ZHYa/NaRrH7miwPjq
z+YDTuBJe+5GqxSCAuhlOajpE0K53wPnWyHOlGwMQFXpDpD1xbfr6ci3YU31hs64QIr8gGJbPNrH
YvqmN2evsouoPXNDzf+YENNdLhl2D54CAZL0+YQWgYQS9JQiCrGWGhlqV5KFFywAMemvX7NDFJOo
r22hWEoFNTvkZ4IxL8kvsfwDVj3zgNBE9mKe5pI/5Bk9fA8IkI1vIpNBN+z0SPWN234AQU65+eVs
kJngSq+vIBk47CmRNW5lX7LBb1GgejI5/RJF7d5X7ahl3rBwVtNYuIhbAELgEkga+BGq+c7vwnCz
iXG48VqIV+LosktwgKxtiUrUH4aujxxDwvBrDpRA2pCFUrgvyJkRyBaYIGDOen38nzTuBbkdYYFP
M/56FErLFcrBdKZGGh4FbNTxpzwET1oXRNLIo0Dp/j1c2Ivw8n/p8edpl7mDXx3praRAWv4xwDqr
nbKKnG5KDZ+65cb5j+DPEI3ZBIutiOd53XNYbCpVB3zVbd/DRVkWdB4mC/UStAH02ElAC/gLif/e
oe57QVrK3EY1pB9euLYChRl9H7SmyIGgnEo5aCr0byro3FdPiBMlS4tUX8ubryc0fp59XvV1ydXg
X3wx9qW2p27Wf8+rpqA62mYmOjwSdScV2HLXtdl4WCPfnzv13wKDBMgPhsYwKqBUmucF2i8ZwZBl
/N/9bAM8m6bUNVWTi8TIvvxxDcXM7ZnbVoqjX2N8J1HFBoKxJ9pcAc4kq7FXRBIpGs3disnVHuEE
Om61wuNEEXD/gFzii9Sw+0MLQBfCNjvStTWPSkz2dJtQsdypUD9jxt+8rSenv5Af88sirFwoYyIP
D1oXdHE9cNRQSLAK5X/su1xf7u4ZZj7FdYIZ8sIAhuUW49LFdeYj0Cl1Z5aYXFANuAhgSA/G4kQE
88QrbPlPH/doHBpYWmvKz+2Wb0uPqmFtg/et/yEWl5lYvg8nE/SCsbSqoMkOGySNBcEPQBXHTOx5
npsjRi4IgEwLAT+J6y993Djh5jV3WDMMWjC3vDf4sJUeb2wHytR/mfr002iQ6Y6jJECrryaQ95yU
lI8CSoLA4W3RkgmosQW4SjYv6usNw4ut1h+mwlbNbQ0XliDCxZrJuPBUX7D9oa6teE/RlPJcHmBf
PedXHUzNH+JqfByX5aHImMHXTUmY6U9xxtgL1me0TeV6gAvC94z7XLyCpyC2VJepc1KCZan8wSnP
E28Y4ZvjyOEBviqJuMzTjNaGNog1Sn0BAJs0N20NasR2vuXC46iLToKKCw277nwEgpOWeFxmifiW
y8sNSO40dC2bS73T/3kkB4wzGbQUcbZYOCw0gFp1yQOho7tb/hsFjIY+HWOeVdRTW13n7cB77j55
cRitu0hxuTWq/ds+O+Q6zmp8Bzdr+aFbn3kyYaBEy+No073hPRR+VNZWcCD2mxg7Rck6X9CBO47v
igT8rBpQhnqGt8rui3hoDZLyhvEDT0PkDxwNuDZ2+qXV38jN0yWVmu9hpfwqoj/fuOrTBj27ZDhB
7GerMnj2lyveBfllXS9oouOYYb9J9lv6DWqIRB4nLhhMZYReMKdeXb3Ix1yB5/RKphmgm2p+77Lp
qIMaCMijLEI50qHJWopRdFU/1uLfbT2NXQxJ8OxFMVRHU+Iqa4VXQpyfrs9SBn+OcQjnrFYkje52
6KWmpV5n0Tio4hLmyLer92nswoh/6IbY06XrELavDQOCqNeaNy+w2M5SnVL6eb3qp0YFfvs9xe/O
0nDYrZAmeFLMGIHq0BzIhXkmpm6cQMHIvmgDcjxZtzymcsKOpi76BXVxPjJUUOMBmqE4GoaRUjRX
tl8Ty7P8CiZf07cBbvkwH2uMVWlOhEbduDfE4aDsFvywWsdT7X6efcxOdnbSDcPh40mn6QkhFpuw
PBn2nvJfn56pO1quSGNKNiHMy2tRS/RmODRsGtrZaOd/U9jW3rVr7cXsJvbYPfsHkhFz8oiZMA9k
SHIIOQIV0E6lp656hulfWF7+t8FOlB9CZ8jfjlu04k47LrwCxpXaztbjfJKZYnOpGHg73xmdyS21
m6+faPKN8hTgbq9NeLrCbMqFxQOe8fBtu2y8WgaZHomGHzLufpNcq0TYGy0UNGp+bCshnKxSyV1L
LEYUhixIVobA0UNfdCwTzXTzh4EGQjWFhrwUAQNID4fTPQjV4Xj/phYqeEsK+OmUvjZgOu/hiWfQ
nZEfJaZRSsdkxOlSlF/UOT5bd+JT8wV/r1by32lyo2VhTDMMO7JOa7TVFiLDgzweMqEtOz9YYyuG
tSqmQwn0DdNKAqF5EbyIFiTOHMInlUQL1+Ju8Wz0uREM+BqjvdCLJ13pvv8vSkP7/XbFARd45Lx1
HcweukF3FBjr2YE97i758wqA7rH6YsYyJTL2RobdzhJczgBgCRS+ZKZYjOGlrn4jGVHSwE3bebRd
UFrhmytLWKtLs0jMe867SeE5KmSchucxRGzq3Lzo5NMhjH+BJ6RMqcupaYcXaR05aXFpcrIPmK3G
TrBv0xvaGpBm3KKL379936LxPx2RUXHiHto7p48yd7MzGnjWwjMM74tS6aWfnRqW3v1/uodTDDqg
GyUwlUMq4cjyXgLiWRl1Xzl2Fy0Og1LvByg4K+WqLBs7asdfIO8eLVhoXTTILZkiIm0dcWHrz1Kf
4AHx07823COtyrzFxCWWhAObnwx6Z+8jViQgATwMngC31YdNp8wjzeKMqojY5vcf4gjtzbk4AfZ9
OOVbqqhJFgLxnYMm8I3A7vHF7ljYyJ4QD34LJsYNckru8iUQk/DL3pX26ObTm9owE4ib2cq1m1ca
eRRA0Y8arVh2TA6ucf/EmC3LWZWhG7UxzFx0oR+K8MBFHUrttIFbhr5GlEHHOWdP5ORCX6DwHSVi
KLGRXM3EME1Xf786uWNUQ04VsV9nQQrVp9Jxp1SQUw+Ur18tTG+KuMhWYE9ulNdsw6ZJJVCd+xgG
/6SBowcCSgkuhnGRB1yA3HlKC2nqM0QnL/ggjVdn1Goq+Uy73ba6R+EQzbza+F5YJHsEC0VpT+iy
gTakl33chdjhgi5G2DBHufN/9/6btoyEvanNgZdrQDpSpI4CE8ayA1xClc6goWf9RWtcwf6KqsFp
bJPZWlPRkc+mibpsVJXIKWmiWfKJNbdYtiuBf5oyOFLpaTL3Z5Liiirs2WXsSLDhPY4q6RHw2esr
XI7Y047SizJNE0ax/6V+v6mgYmQJY/2h7XlmlACzQO6wcg+R2IzHVoioh1vtD9ZMrZG/QBJfKIvN
dRGOg6hGlYUpoKJnkJymKufsCAfAkodXyVqGH8LUPy7LKcF3crIgjdK0SRWyCmvaCi1uy6MsjSab
YjCFYlmSK4SiwdyVLvcxRztAWMFiWcdw3OP/EVUElsoUjhK+CzH2KaEmEeJQzjKAYAdqKxdwerTW
y9xae0T6NhdBQ+xwCNZJmwrD85BKIry9sy5h4WFplxDInX1kmd3cGocY2z9PhmVHyzA2DiFQXUmu
Af3Uek7OpFUIIeCiZ31JTagc+Havwyea+inxcJ8iEPBwU7joP5XHo4bHNGiHZSAYCGgzKqhmVN9Q
0PGtc4V+BXcddqRauxKycfkf8T8QzStEDnbl3LLL+IpTnnLOh6Eayyp73jt5BXWCYgkCLF6RiaKU
eSu2rdKq8X9+JFFQ0bF09En7P+Md0zFgDyWnR06oM/+0FGtIjEZkJWZGRsOpaisFDOZB9dFOWQMC
EgMNmttxS5X7PkVjxHBqkFybJ3WCRhKPasDH+lgg2ufL2EsmJEKY5ColALdY45pgcAwGC+pprOoi
O5N9SaFDdS7OyL7APiwKXc/TKac/dAk8XOu7RDuAl8QEZbk+73tBpGTOSorsogyCPb1WlAFmQDdR
9Nj+uzqmfecWZsDmfNBwlU6QDaJIsmU7lQrRuYR7NBgSpKd3J3JUYThg4ZWjcpHw9ek1g+2tshI9
RXWbBewPDeaJMeCb72lkH/e208bEUkYC3vFe9HqEfi0NsCB//lmYhOuURLO5NFqx6ZxhZMX+XF4Y
CKcW7xYCKxfsNnWgH38GQTCRrjMX/hGEWimvXf6UaAmUZNYeFbRtlypMtW0z4tvzTnZo8KFuAPlo
+KPG4zPI7ftLYNLbsu6TRqTQblh0BhEp21LNEYCEBEQwdUg6YTlfwVSqPhVVfZ7MFWj/OD+vJ3R5
c2l4FL1azegsEWnQBvT81d/1ejx1mRvKeyDXgTNI/woSylic/EJcqn9CCqehkOxrZVSPW3xIITq4
8K0KETcwmLWAogsCwf9knmrdw9gS+pROU2UyTK8JctFSbMoxXevruRNv/IMJ5OP5j/iPvoBIYGtN
XwV5txF8qm0SfekLWNdT3OVFhlIUfWcbWAlZkcWpLtHVGSN6nPb1BQIFf44/nRNChJlzBPeG0RUs
Dne2Ng3I2T3zUh0msquhkygy/T7ZTKiA/DKZuEtZqOJlyvDaq9TbyqeEKZWg0CVpgk1c7s1voVmw
v67kSuQrsXiu1jeNDw8GWasjGjwvkD1vIywLDxtjSDExIUHak22yJ56rsU0kcyn6q4C3t4nxzRek
9AlKt4mZBfBmCznempEhsLkt5iM/VjOJ3Hd2KKlOrfxyPF4rUpf0tCPfUO6jMSuwxV3Sd5/VjrTb
YxGS+KvSn+KD3/wXOJFtSJo8GQVIdjNT1duZIsNxBqF3tkEOfhyAf9XOAbagOuJorAV1WdayqglU
/bGngivZfaDda29xFWi9O/1CcWvknbNuqB1vk5VfXOmYwadkHzWsgKeKXBsSPhzBedVPJZHiSTeg
wVgDNIRcdr58MqRBFGt6JtY=
`pragma protect end_protected

