/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
aB5EHAkrB6NT/NTMoBINikqg8EwKYDaK54FjPax2CptnClXJaFSk1P6Y/9u3FWJjIsff+dSOe3bi
iAx0iPp0pZj8xWoo7D2kuRg+plJgYo3eEH77LyOgJ8X7XStkvgjstpA8MmqOdtjObA2+nWfOXV+w
qbssx3RmnSBBdhARD6rqOFwTf7/3cDuK7QTo3GD8GmkOY+DCob0TXNl7kc1BlYaNbdaJok+U9OEg
YjjGCk5uikHjY6JmbT5Bd71P+OPQhQWHoUBkHUIrhbxZIfDop7LhnylOAsOUmH6p7xY7O9pS50TQ
NpvG9Wsvg8pUSyb0Hyecew+1A6TcJyANzCU7xg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="MxahWTeDMTwz2fyFkxR0OEw6OdcfpBcLNutRaEfsJI4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1050720)
`pragma protect data_block
hbfFuBI0Xp74waLCAt9YsNMb6t7I3Q5ZkSurTo6y6enHhhHJ+9Q3BKXhTpOUNCV6vEF2bHrSnL2y
xP2dPhLzHp9D/KdFK9UYQ2t/PmTBNwTIpcI5JRC1UyQr13sLiq316VZ4oJMujF5NxFbJa45GJNtr
lCoH5rb9ljth02pzHDYVjBAjJLEcqn+Np6hnhNgCjfNhfo7Bxz2lAKrZPoJ5z9D2PANGtVSxDZdm
s8pRAQHzMG0dp/seQgJ+vsCzla+0T6QHvY8OQQlRvdmL4mo/des3xrZ4XCl+wGcscs+po1CkLFta
ZdcNofke/dnJgjIrFkuhhGUstAk9EjR+Ubb8y8WlP1ZuM6ZOtiQgwZvCg1qInMxR9UKtCwmuunCW
JHBUiBIeGhmpIzM3U8YHWh9bV+HE1sNS2tLqyd0uyltlJfGEi26iiPKWgNq2s0aufqta8utjMCRH
CdwHGuaOBIXC/slqmcEtbUD2mUE//jaed/RXCLUP+QBpTXMcCPqph4ketT8G43SdqKAn/OwxPK+D
Br8x6I7NNhZ0Xcilk145t343SXW4SGmKvzDcAqSOG7La94LLTEGiRSQ/wcdeXWwz3qxqvPi4Isz5
NtcaO9o/rZ9Je+ACzLQDtEmghct7ndgkpr8H/oda5VqZ5gJBm1mwJWwt3j/qlWyn70AB1fOZAgkr
7xqZTdIpSKH/Gu6ZGLUDk2YkFxdSqgd1zMHAvt5ecVkB35AQitWUqWqn8Eb0/OpHgKm9wAebGAv6
fQSu+vjpqyfqjmM5BKmDDrFw9fomEt76i+X3tFBv1A6lFyIJ4+9AHNheU+mhvRtUculA+Q35NpQP
1ZqkkrlF5JHLVmYTOwk/IoaCPyeF25MLUHBP6esQorwB93IGMMDtFoHQ8OFnqvKD9HyQ+3BOTera
/XK8kWNapD8I0nj3eMolmWQ3/DpifJFQpJGFPtPcYjtBqN1aghf7OlQuuZDwYjjBbgwv4cNQkPKe
BMlpFYowepBvt9ZU0oEJLKu+6phtBmNRX2+zPCt14zJWghzPqDnozNgRGzDRsmMNn4lNgMqmYh5u
yt/UoneBV8hnGjCnKDOo28njkNJAysMLIaKi59i2U7iWLtQaejKhMh1+wvMUlrGNfiTasM9ftjqt
IkVrq+FNVgxdqjYpGy+xfGDVEQYEnqJT3E9rwnnXsOpr540BguaVfZfqDKdQ8VPYL7cZ3g6EMub3
OA9Cuj8REDXHp7yF9+Kv1P0+CF+V6kAiXuQ4l2Be3lrGlpY6T6t/2qOeOe8I22VRt3BjQmYA7InF
/9lDvgFtK8scNz/SPNIquCZ2VolSsvQoAVdEuQOK8uwy4i6lj1FirK0W6SMeD3DrlZQChRhfNlHF
n+k73u74ldA9NUDp1j+4zlCPW2C9c7XOKBUsEzHihpIe/5YnzJEBYtISQjuqksI8papt5GnngaGu
SBfNKBtDHbpEX8NQ8MgwrPmEvhZMqF3V5IB8EutPhphF7hSkIL+GEfr+0hujdRegqtrtiatmwC3z
Oi3popWGwCs0rfpnOHVVfeDrvfpXE2v7t6yNHzwc0n9bBIjrHNSRajdsrt7sOvMzmgmcI6BlJk2s
9y3yjaXbJFunBsGDPglullOV07G3WDD3AdA/otjvFbxB3Sl9swHJFGPRVYJD+W2TwiGo+Qsa5yLc
u/VWNhi4ynnbH0x4S+wr4Dzz582AgU12+8JG1ds+i/fhCsyEeC362QSxkc4epwx7uxIziW3dkK6E
CTy0UmpwtVc6pMM7dPFWnV3EaAzTuV9w4cWVWQvtWvdYk1ScdILkofwDIt6a3XP1uyd6QAGKBjTB
ornqb2CCuBgVA/TzEtNj5yVwYV/CuZXwMoWmgaGfOBpSotuYRR8JLR9JJYmJSGSXIjcnRXS49VgV
17zDtMyaMTn/YsOXh1G3ISqbQ9ygmb6bFZxUSy5j3SB5t/hU2Ex3VIpjIPZZXmxUjylrJhpDxV8E
vzT1n7qQsIIcz3O1SYF6joqsYiX9cuxHjEv9hMXV4KwWT6TYUWatOgjyW9rVpsttKRVHiKYuu5oQ
FO4Ee1kqu6DiAfW2sW0rMIG8dgdsdRuRhKFsJP94C9CRBjlBAMCDNk6n1lSRWfMnEw9x5dOnjIXX
lPwvalmKn4mJG/qDMLyew7bjEiE3iDguUEzV3sWK09NblX58xWe+TW+ZvE+vaYyl8yMmRLyN8UpD
/aIkGOKqI4cdaIyWdqLQDrIcDKUwOx8w7Buvzqj6EnrTSOsLHHmV1uOXXHtmA6sIcuu3zAxy+0mi
RfLTNNVBTUOeLJ3EkA0p8EHXmbWNbyjiXv/JS6Iu+iHmGuLc3fFd5mCdeW2Me3A5biZCO8Cihwfg
Hf5iT4ZrsZYZuN1C492svfhpDS5bCnCPpMFFKVdp3IB9R/i2ghFc10tYJZZ8S65/k698Gu6qxxVC
3np/EGCmt//6uUUQgn9My/QcUJQWbASa6TQB4qVjzCpYPnr0UcshQFIzFImeBeHlo7urqynehCHF
/UV9NNPzR+P0k82tfaBoRBQllsOMGiLEFnWGsyjYzolRdPDVUVU0kJ2FeSuAwN6AwkPLDabO+pbG
crKPHUztw9FWloRbHc9l2AxBq4I3DoDQk3Lk+2NH9kaXsjvzgbWo5B1Xejr+fW8AiSgPFMQHS3mu
iBSiIgKQD1v9rnaREbF60sCqJ6RgNZnjwBaPzmqoWzu1+I13UlhJShRNjphB/i8KJwa9gxNpDRN0
v1fb8rE5cofnpw4ahyu+b8FjT5EY5bkBiEyf8O5Iwd9W0I4e4nSPYIdOiXkqs8VaymAkhuIWJGO2
XaNJhTIL6D7QN3vLfG46M03D5b5sw69PnR1ofHy/5rjOwW43pEksGHgrgj4KmqvqPVrKAzux/jcU
jP2n01aoqrPjkma+otOBtHn498G0bZh+MPsRk4TfIpIJ/VZ066lteX/L7Cb0Bkz6YaPB0HbBfYUv
s7hY5Ax4NTmvosG6h5Owdta1E3NgQtFB4twFhT7STuE25/kqgP0kHD4trhMW6VL4fp/N+/Djl5u5
O4fFwgTGWwpge6J1LOwqSXICmo3Saor6gskUWf+hABjNlqNKX9D5WI9MvF3QcztGxLgQyeffdSI6
1+4Bhz684V4PAv15v+sLgkAvJnm5Rk0dL/PUSZwS6yybAlwHdlcrsaba0yuIKDvRIIACq/X1Dcpm
KZAVpGrrZs59isDT0KABa2QLKP16evkkcA5WPXomBaMJX6KS93nBwO405VF1S8q+tbMusOQFjg4j
8byclGx2It99PZH2nARquRZ+EpXtaJB9k2EaOpB/FZGMipOxeccKmkAvVOUs76ZuNcETLPuM5uVG
swx85q/BjLaOhC/n4fJe17HmTFROgsgGyzCesnxqUR4VGmIWQ2kZBtsMpCguiTUgIeaoaoMtkT+9
0xkH+6WiRiuIUy461N/wDdgmwQCQtQCDOujVeTsWFqrm65FTd3FSUmSYmvSAe+GuYOWzfq7XGNc2
mUNnC8NDQ1NlJwxBRSWnTWpXA2TIk7h5snj/I3uJKNGTa8fVS9qjVP0/byOfcuS23RuleHCFS2ii
Rc+7j+RkP5b9ZCIbxjOr9MS0FHmVoyRg8GFLHvdbAeCfLHq0vW2xxYWxSJXQ7B+cRTmlv1/rfXIn
zmZYJ/y4opRffOgvdQWXN45oplzl7Z5I8K55MCFprozbwYdD9IUj0D2xEVh1rxPGSThl06o4gSbJ
XiSdz4Jnoyps5McFs2h9L/o/+Wy9gWMC2Jaqlrc9v5KJmHGpw84eePtOs5XppNtma9iuTfMtcrkq
2gQifDEYlARVGeE68tgQFEi/+kH/npyXp3diXuZxFiFK/fRvRhjJw+puSpPHRSmD62TjwuBBtxkE
0b75raNkRRaABiwGhv8feyUCG8NlR7gLtGQ6HBUjvccijvfmPs7VOcBk+rnEQlkm0sXzf4gl1YFI
j81QkkMM6chRmsysdiKG7TG5jdEsfwJ+g0tuL0TsIW/J3CL+FTGgZjga1z28k8hZ7x4LxvFklG5Z
/1+UkN2IpCoj1A/oV4ATeQTj4lTPkX49TM+F7FsKSZpbEWoYwG5GYTa6H/3BQ0XWp/xR9vWHEgqP
OQEL5Ig6ED924BJWRj3PTH//EGnMj8EW576fS4ZxP3SCZ0aFDjvnDkK6lNCwjsPM+BNDgQE52gm+
EvAmj22YNWeFmWRqeYhO0wIwjpXp3djY3KpCVqKFqRBUHMMeRfvfR/ndqwWpsTk/oHffT9XMG14s
BR49RB/d4dHybsmLW8jX5pQRe7f2sJUEtOQuiTiucqfajkuZ3pIfyW2EkVZYmmk/gYWRjllX9+ux
Rrm7kmXrPFfFzv+t2tVNbxLCOGB1Y6NvEArrWDI1Th/e9Drx+dxj/unFFJPfeh83DF87+9d7bsKc
z7qC9gEn+MbAleXYoVlaZxb2QndWnX+T38zVvbvQBclJ25Hu8dSrVW6akqb88xmZVq+/G7A8ZjcM
8DOY+RXSk7jgIIAz2TLcdBf6rCqqquIF1PE80aY/3AviLiCfDPN3+RcuDW0w08y2Tj6Xw64DiBma
pghbWeUlukFhiSJ0Cvgfo4fwBZxbKB1x0iuCp+jtJQhO5XoYb6A07sRMvKo7Odb2WIZ6gV4qzymV
6iY4JLT6b6+vsutEwJxOU7Ar7YISp2iGjzlxhyFTHWY6yTck0muTKcHSf5gwMcnrI0hWpjMSE/jO
nM14ufzLkaxsllrRjg3mi3gi8jxYN56Zo77GriD22VsehF+Asep9ofAiP9C26a4AMFt0Hpm8jWBW
u6YkocDx1P10EqClituXlNf8r8lMbOfDp2Sr3VhFDwhakUYKyOXEbXsbFjiv5wny4OjdNcvKiIOc
/DB2jQuXaSZ43IILE5YElNxUx5lVLfxX7dBqpzZCVNXiEkv4F+5A6JEYv7YVxD0BU9EB8Q30/tu7
F88mCbaCzppPWSlxTClMI3WsbzNyxni6e+CuIjeuiPOxAo7+HtT8C+DZj25VBYo9PXpt7NEt0+YU
cshsyJIxqUcvlVYaFf9tCyQKsxDmoz8W/OshZdKe35A3p8HzKgzw5/eCCOTOAXkivbamvl/MW6pM
AFLhEtZfWmY6v+Chmxry5vGaK4Udriyp/I8/CqDkc91jPB+kAcRYygDQP7EJSrWnysRgYXzhO6lm
9snJ1UsBWHe2IyMrLwIQpoiOFPIZGuyWkPbREnofuTgcpZ45C2LWBO4CdNCqOEOUZxKKeFRxsIWy
gRdHaZLtpejnanzMCusRKmCA4CGIje8JHzoBqG+Gw7vHR9uzBM6RwUQsk6G0UuU/xjFUdyhQK7+G
RrgsynZWCFRJyT109lVhtq6BLcSE9JRJ4MzYVsJ/qzRRiQFW8RzYfs1kYXKlkS4s5Cwg5aPhjebH
0lUTitaiZRR9ZNfYFqc8Rxo6cATb3dnccTXBCPNW7ukFu034yvYxlJLCMI4U48zmotQOOAnypK0R
vV7DKddhoj5RJAYisNpGb7ZsqFvat7IMASqhACXLwREhNQtAVJs9OStUHWOUDWRBXl0jqCpvc0j/
k9aEXrIKfO0p/ZL6TcXTm3ENsJrmAMzQZyQSMWHCLF18xMmhRnccdoU/0K6EAR9IYb7It3IyeCBT
nJBh3quv8kGzjptzzBFNCDiAOxqpLblDavwprpSHlipaIRJmda2kzpCBhjCKpmWknCWeLlRt2zZw
H9Gf21Ii0y0vTvya6nmh9Yoe2EfbjQ1INuii0VUxpSZ+jtpKO8oQilPSgDwHRyiqSPfgNtWc15+M
wNkq/tqb8F6lgKdPwRRsgGcsq1fmo/C1K5sfvP4FCuX/gEa0LXS6kpkAlzXE+MUuggxtydaY+hPt
x631grdABypPTFsjbMgLkLKPfPTx2RMKDZAfDUjeotbkfxZVrSEptxP1/BNf6QCmlwJqr1u7SQl3
1eDi8Ey9FPOeG9zU3g2XLpNYVA2ntokNROPJRG+pILvAqEF2X+Mvfy3EOuxvGV2DOZZOJFcgoJgC
FjFb1l45EKeBL+8WVarcwcWuuLehROnQg/J4OyoKuuHxQuWss9hykwGQqBaU2axdx71C2YfaDwwO
4GOS6825UUMeBc6gYt/YzPawFhUkXtJHFNEU8VPrJy2G8clq10HHPNLf0peHbQUMBkr44AyHbF+K
0f1KF9hsMMS0RkK8rbZFdTU1uI18+hoXDGr00oZN0lRX3TF6ft0pIJ9o9w48TYndkZOmcidM96BR
tuh9qR94WysqIN8EevLoP51DjtvSKf2pcEhA7myFtJQwW7BAFvggkVA9vb5mlPtkbK9P2Q5GmJQD
0kuk7Z08K6A8i0qdC/dnLUMyI25qwJTWHDOm9n2TXW0REtkZnOGlQkFTFU3koXPaaj/X1Dzipj+f
PvQXREjCHDp7bOBApDjIxK/fsn3CKjYCUOSs2FoAfBnjXxO9E/yi9EQuZUEePD+VDfhj3CZ4Dfw0
wgYfxXjUnEDpWqfrbjKt2JtesTeGtA8e+3EyHdbuWMzrenRyg/HZlj9Bp3f8xD/5fxRhDPgyxlVZ
lFrxclIE2DfoIqYOROK7RBJ1hZmuFfqkcTUr5EEEFoQAHmbOpe2z5XwLVC3hS09oyAfTX8s98Dw+
uigwR8GmXBTYeQaRATTjQMmzNWVBZua7VFzWCYKlZLPp9J1Lj72hLDRf4m+qGKKmHjnuqvIdDkIR
IYvZz9G+0dv/RrEUgklFMWZcBnT4C9tMO8mzvFpTZkIQ79rubbtgcme6Lm2HOzUIlfn2q8UzSgYM
356gvYjme0rvDIzm32MrOcmZGpMkZZRPtedSKA3kw05CFIGThGGV8EqqrVnuhYhifM+aL7BqTdZE
EMGidLkWidVP60CbylHvvMwWDBRRAj3/v/e2Jv2+ZSoBMIIROOEsPwMMUIMUZ3WYbSUlMQqtRMkW
ortqnjjnHSnol+BCg0NLJhyZgoHSAHjhUJgtXlMKJBvAy6dwvcqXiunA0A1Te1908/20eFmjac8y
kPVXABkqBmRnmPIIpOKNDiBfWlSjP1seRZXMJTah4CGALmCnxPFA0IiV/Ah+8ABKf2p64CISwVwS
/Y+IbEK/lcMwC7hTh8j72SXGLrLDVZZqjQruMMs4siGxFTjmTYbOgevng5DfcPGmJY1TzE9YNxBf
W6ULbyeMWX0wPLv8uaCUJsWt2X+uJxTvH5P+ZNsfsKRua2cOl9N9fLo0TInakAEwT7tOMnI90XA6
Jqt+XDbnE2C4A/ahLM49JH9oVYvkjEVZODY1Vodft6Qi4frOrdGASlnHgWULPpVMw53XhSVRYmrK
4kdQUyNifxbkrc7GOqTKf44pWCvCnT1vwFHCayson+Pfcx4lXRJ3x9/31XWkyaNmcKQ9y7H3aE4X
KhRZZ+hsKYUDdvKtA42BXHlkb2Rj7iqjkO+D6YaRToLqYcgRJkiUSa5yAuIVyGeIT0ItxwzbaVFm
PsEjVhQGcZ7x5dIRFJrNzEESP8m41Az7qE9pPIBLr/Mbgft14c8sYrtVIgplFK0YcHKiNsZbck2q
i+TC2KWMFylJxC9fuM+C0AIUr/7QfqSsXkqHSq0G7ngESLBzn6I6sCMpcIx5Ej0Ky9/G0EC1+za8
KyFPb5KBp1WnH0d+7SsV5UoSDpB/7DfGJZit8Lkav7FDDXLEPZeAPMBbm94+/hqnY92q3AZX8XBs
l9Ix51L/fT1TAaQooDWYivmGkq7SPnQgqEPWo4xCdP3ZoqvfOxesv6/UEpHtowXVrEP/QjcidhdN
dGW+PZMZxos9BL+conjyTezwPPIvPxd5GV2g5W/1FEijX4AUmkerYILVvsYH6DajlGeI6x83ixp+
RtTrAz/RcWD8l1R99J8qK9MGiYMHuloNOKskoO+K3ReczyDTQLGAKYEHePeZ1s8hCzpXclyy+h8L
w/IqtElnkqByiRjVfCP448qVVxckXHQdvzbMrhuWwsaW5jYHpiDfV8zc2az3YRVTHOAdAVQXJN8u
sPUfioRq1NSEHTNnLjRJsZtr5Eiei2KnxID7vY9fq5e66Ie74EBQYmCQz2wT+thjQAbe3t5U9VTk
nm5R0hdgIaNymlT+2Fq+B3cEIh0fFrpwJrBDeHeenyG60GV805vwBSp8nE96x0uU00avV4Yblo1A
jG9MYRTpk+ZxdNxb3pGF65diih4z+6RtTpBfHA8FyKgH1CIeqodxLjjCNxJ8tx9Bgyl0Dujw1RxI
0nbV65qz89K/KvcItjq1KTJm5JPHwqZd8CycjgheycQF53dIvyK0tgCycTIlXeVCcumergMuz1lf
bnCafUS9RKEOwwNAqolad/IsF+nIEGpYBkZIIOsnOUdbBy8tfgzKrPx4ThjRKdSwdE4T3fv4mSwj
qtPWWhJ582WHzu4pHrVZF3Do0OaC0E9+vrxoRXfayS44DfpaXoIopDJg8VUExQKwu/TCIq593Mtt
4iog2CwZA98rP4ySBjK/hbmbtIPo9nia0D1mJ4ZjU8DGfBGCk2o+32PXgc9hcTls735W2RpdVdDD
3/6Py9QvoP2hTwDFLQwPl+HCSFxU++reybfo4GZGPTwgEIDh4/xBSY70HcS15PTtfEiAXjt8ka/H
xDIkK33Aw3Q7P1L4iGym6wjOlBPsfs9j83uYyu3clJCI+FacxLo4vavCMxE+IsdE+DfFaaecCTNn
pfYffZlmFyHpLOg99zRrXFyhl/b80jhzezD06wrw43DnQUxEG713YeKwVeweWR9kKyHEIAlFrnYL
bZcoA++KejwPDmi91IKH0Z/Sj/VZWaUY/Mxp6BWpm3ykGvhNiyaGYMQJ9tvHvAqOt2fMPY5xw/Nn
jVvZ2q823fW59B0XOfVF5AYMFAWNrpMwl3bGbiWUyeqwS5ui3nWhZ6uV9fvMcAKFvG9MfUJLcJON
pX71okKCCBGrHXrmzzKfoY38dqBz0oBSCSBVci7IoMd6Gjz8oJlV+RA9DFkrsjgYAIZ0gOWbbYZ7
ReYEC//4u/1XT793CYQ+dt1fDaR/CaeFA510YVEEG7FnZSez+LbXtZDxNBwgE8MDxeuyOE54BM7z
FtT90gjycR3gYMp0bXDg0zHm8D0tLvGQrEWdCAsdE32SUUHGUkRNe+EDoCz65Ek7g8u5b26eUVyN
FbQOCuQa9fAMB4VmaRyU3Z8xWZ/JHa+TUVztTdvaDUuj0yXWTbCD1g1mFo+w0I/fvRzyRyse9o1x
WV1TCaYpxyyIYuXWzjPS+LtUk4NwnAAAmGCb5aG6V2K+YgXCK2gC1XuttZu2IgKiDPgoRAcZp5AC
e7P7HlDNWBxNMioQQ8dxLAQxfTS/iKV13w5DMB8j1duZRt1dzkT6N7erLYGgYrmCH+QsgBEjWvYB
lXBIK+3I0JT5IDhO3HzSqjd64OuY9gCbGrkdI6qU1D1anNtrlQvwEKU8u646xrExGtlsfI1FvXJ6
0jB1shxg/F5w1aktZly1i1CWWxbNTYoy8HdCLNj+LqRTBFLbzbpYOeXzdRAQJX6LiYoH1tT+/UEa
w8r6MvmMivpycHL4W1EDWA4pjU2JC5E46SPUv7Ktx4DfVQf8pWSVPH2rQgTEFcdNvu6MGeLkXjkP
Vq8s589vEXw/IE/lLt5wX4Yx7u03dRYDo2/FKtlIvD28UageQFAYshGl25YXq8LWWHtcqRiByKD6
LmNhc5twtpO3g2ByevEE6957aKlAnkCuWzVdyX4yrKhuDXxh5K5pSKY5ntfhtvKpnKEwuv8MLHzy
o10pySeYjMaDf0dNvthwBixh3rPCtw2C9bC0gG9UFWYo4a7CBYiFj9VrcB3Qx6Qd8s2tH2LtjCtH
YkppYIZlpx5YfYLFfCtIXSNdu7qeqCLZQ3quuspHGtSmcXkTewq4XsAx6lRUovvBpe6FQPyFvnRw
rEyIvKXNyEL8mOqRHtoDwnSZ+gXUCc0zbJgzZ8aSMQX1VRoqJd/WBo284XAJdPiT6Iv4IgOwBmcJ
UKBga6eki/GHYJPvIBKeOndqVTnJTIXQssPvuXIWfp6CkBVWftBxaqMtMReU0vcOqw6H9VpxNO9z
Rm0ZIdrGJourngidu+jyL6Ar5VR9h+ObczTaEBcqPXP8TF7Zr5gbSoGU/3JYH59L9fG7T6L3o6d6
Tj4IC/lyU8ahuurfzuE0BvAaMwWHaUY0Gj6zj7eAJIzc0xIik3U3EwbI5aXOpyjJE5Yxj8HS4qQx
OyppQfz46Ok8WxWcKB5AvbCMGPsh2lgU3JSTorMq6rj7JZzCryU4DsAaCmmgg5wfRCb15kj7RTTp
4kG+C4uReyaBO4CvgtR40CVkk94rK2Aoi/YOBv/QcQP/4FQPUF7CASkUApgSN5oDxfoVs8xVGgUT
YqXbZ/cvEuZadfBkSoB9sMZBq6rSmYI6VaaQDxD8ODd3eU02NJm9a4F5X9cZLzN1R4D9O/j+SYhq
ER9vOE+LPegW4waX4l3WbDc5o0jMW4h21rFY6hSRDQQ0AJo4m8i3tNnZ34ARiNLYIlHv6s/zQ5/S
BNtkVwRY7a55bQFB4JYkhQ3oZJPfTzzPf31vhIqN6Axn6jNfNM+NaVN76kiyF2fH5upSBqRuUpo/
yzsqwheWunnziiobqR8xo5ruiqv2cnrpGDF9Rgib1M+O0VriZ8YEJ3Pqva3vFoEmrJaNW1PqK5ql
nzMkbZ0mYKkIqOFBk3MWNXwYz+5K0WZoEVcr2RiVdM5ayrvmZJA8/wQanY08GqUZc2AbCuRu7LUu
5IelkJCUYAEJdL23dYUgaPQvKXyFwUmYmRPEoENGB9gRM8QRKPuz8nouUVhQi2n6cDoC41hgd7mF
8jKNneEKiX34MMDrBh2gavrdfBkHYa2t4gJbu7pYTtxe1dhZgNIgllZdO9vl4ipCwHCpdYFD5gmS
tns3VTx5IkurglGzdtoE55tsISoLKaTr7KRQYTc1rqtctRSOgZ/cIEB5ZPG4hdYnUCJr36rb9Po9
YTIxMsBdvZ15p/xUcGgftgLmhAg+qeFFHo1A8PXNMGcxw/KD/7nY4rbmg+biAxaRwY/NKR52ZZbT
Vaqzu9K7mVAu9HdeZX+Ks6B3+1VnWUsUnxlXPM9KiIXwbr3jyNAVcuwFMipcBJhlFXcuy87jVQJg
cRAAYongrpql4wQM9L8oJWnsmEYCg7pqGP/LcF8+DRgNNlymaT9A3rjY0ioFTIoM5s9FfWxsMgM2
WvU5an7J6l2qahQYkBXD6Qdj9QmHAAvEkG+IaFPX85u0SavsAniZPR1jrokncZVb20irk2OkVVbt
KLLY816twYh65giBH7xIlNZaVeciNsN2IdX5DtD8LjHEfb2FSZwTY/FWvO5mCUILb4W2c4b5+7uy
qUSLF+5BBx6YyXSy2jOc1QLhgjy3EEWHvCwfa/E919ElHLG+Nm714F3BaS2fJv/TqTG4zFWHVK4F
T2iYcFRZ5H6L4NOgWWomaQD+0WLh8xK9N5ERvQU9SfJgu41ZaLbCKPjO31LnHhc126RIk1TuHBzh
ROneVwdr3YklR1tyEreOhdlW74K1RJD98VKdkxpiAt88KeVFea98OxHevOqTqnB4GLClK0hlUMVv
qgMFFmBni2OuaXGKspfLJecv3icz3Cy0/uQ9+QyOAnHF+dhHaKWltI0fsUCKnhjWso/BbnVgpt/4
5Q3QJz4Hoc2hi+kU1JpHTaD+QIaeMy9bZ6WoSKdS+Mr5J89LjQPbnkAoWD6CQiz5GZLoMBZ/ooFG
azlz12iCqK+9eMCLXGpNJCurhr0ZBCpjBrTcbFQMmuucFH0wL2RGcPC/HD8ClKLGgGktDLZP7L7d
5JQ+JscVurTObMkyqWKNiv9W2s5f8RrcQrp+Y/rUNfQCzyBYNvECMri3E+Pp16z4h98U7uBEc1gG
NoeQSsg6NR9Ql+GI1zFtkm1HcKzM0ci+y30CKeMjrgXTzQ8G1k4PISQkBMnGWT8bPYEKrveBUmwc
ZKtsanyIZzMPNtYQquzjG+2i7Zq+05yANkxLwT7UL1h/23SwNI4Wak7y9iSVtnuIossCc2wb4knw
aLci7HcLz4gJCEuCLtHTzSQ0K4wFJe7Nhu6rGiOa3GSvqkRcldFzb/Eu5wPx0VH90/7FfhzMDJXV
iCUcrfHuWl91ZjnAlMruDFXd7nz8hdvWf+wDcU6Cf3CG7gs1GJqpJU9eZviAQYZPWLLyXFYWhVKg
JFW+LGTAO6iAGSWoXkuGg1BoB0Jap8cLLF/Y4Tbfwi9W0sso5O5tf9UXhZ1eWsy+VWDW2cTOHDXH
umRUo2vx3vffmyEkvdFatViCHohNlhE7Qt6ONFHItcwfUmzj66ldHlbmlZTEr+b37xmUeWXnxKwm
w9B3D2NH+zoiNT//AZq4pLc+xKnzM5A/2SDuCPuqEN4rYE+D5c2VK3B4ZtyWOHI6FCaWf/zoxOjM
ih95/Ti4mSJQisGQhM5I4rel1ueEF+Htb/gR0Ixc0AXpRX1QACCTxLgoCfN9j9DZ0c1LtqaOhey/
QVvPt+IB0S9/pYHcebRjR/7BC2P7tupjRGJv5jFmF/jxKvmMdYLvt+/662xFtnVBZNpLW0xRir/j
sy6wPFKYrA/TYZ0gd8BKSHCa6mBYrTQxg1njyFqCZiBF71aBImZniwoKOOZREnzkOzr+6x3LrI/j
L6NcZN0Agj15zimlSpeENpu2SqzX0GWpJgbaMcpd7Qs3jNWtX70wS+vn4QaTV/ZEIk1iEpRr+wQm
TPILQEXWUshm7Dg5rBPYy6Ce1JTNjhH+vklEyUYdRGGm+rPm6XtDvUjSEFUp+BfGYTLoX66Z/DtD
3AP9u4Hc4qfgzoJVgEvAIrjZfj8wOe3kFKK53rDXB3SryunDl5U7oWllS/1ltSCnYGwlIXSzyeJU
QzhCsbHI3Sygja1j3aWY/IqpqTgma7xz2Euljila85HJtDM5Wcgm8d5oGIn5yV6NonMybOfE+Snp
CNZcjdPvNQZtNJfIO+VF2bos+d7cTIvc9Bi2/wEeb/oP/yPBjpv9Dw6Faywze+Zcqphu8wUuhjbR
Erm03l4HO+jdnUxRFDJvnIb+Q1dOy5MIFwlJrfKivzzoHi7YhfYxDuXbYq1C+q6l/5kbXrbKMAYk
NlIioFFQpDPlM4WavFDds3XUAM1wcG5hZhaShs0T55TrrEmTOro7q067SQWe3qx+OzyQ2Xrdbpqw
T//XE9Uqzn7vHQQpIIkuQ22OIO9NaOICMTS5gGvc4EmfZ73rXCehp5YIeRZ50cC/PrMYWzbPZ62W
4TvKH4pfDasrKswwA9iSn8uSdNFHb8bL95zhYFAx+uamCelNKHqrF0koaOyj05rZsn6PeGSlHWFS
6TYlzu944E+Ffr1SGeoM7efqBSMfHeH0hLx4GeNRZaogxpxRNZbGCTik0oAIkx2wPgwOhhzmC8JB
P2BKiSpy7ypEZo/S5AdvQSLQ9b40xN6HwnQ2yIykEchxMY0KYV95+QBCVSYZfU51OF4VcuaP/6a1
X4XUlb/N+AzwN2ZGhy+07zsBwPWrNpJg82GS2ke7ri5ROSAENLbvywe8W5UPWYL6eAAOv74L0dsX
ybYWok6NI7CiwZrT4PQihHiTz60rXYQaCxkxR2nZntbfy2pXKDCWQ8Dms1E29CCFkPgacfGNDJcJ
IXeKFFqfH42druBE3CMeMKNdMjbWGG6tCAr1O+biIeX/YwXkk4dRJilGVq9ki4qdIJmVov3DlvZK
u74hM6FkDxzaxRQCF4wQVBXW2tb5LMa8EG1/a9xSsfyRjuE0bB0UXz/I/+un4s6QUT/+O9JCAJjO
fKi2oADm0zHIGnvVRgXnfV1qBv9WqrCyq27prZAes7Cf2gwAdykrEaxrsi3jYGc/ppX1p8WfHwcI
33etdDZVzvbfloBsClcEQaEWjYVHU3oeE5qVyACj1yTZkttGuf9++YSxb9CEHURQU5gD01G6inu1
/sOrfe5+LFzJdzlTvQgBm8A5h0Pu7bfE7xvBVifQ3VK+166Q2N9byRHe2ZaycKGuO0ObQ51ukG02
YjYB/oWaxX42CU7IoNS11M7OAoPNI8ugirzCKBTDjd5fEA8FiPbg8MGlSkycWNNDkKG8pvpQfrxz
AISDh0FW68KbzbkdIs+Y6nR8JyUN3cvgM0w4HY4IudC6FWWsMBntX2fKG7xfVQtshSFeNhddtFme
oB9e3TAX8puUvJbc2tTzynWCGEUP3RH2IyiaNuPYxLWMb6xL/j7lUwLgIvKudpbnpeuC+ZCU7VN+
2CgluXvhdTbKzX+Y0eE+h/7d2CsmwImvqcK/Qzurri461hL9o5V6VutXCMOLTwcA4tkvQCZ7rz9D
AFYa8vNk0qjCWCpXZAoIQrBoteD2M2j1zJtBXvhp56kSa/M3+waiYdarEwvuoSZB87nUiTPtcB36
7Vz9cUL60RcIZoCmljnyK8qf3Pfn8a6wKRnxfo8RiqtrkEB86yt7SaIhfnll7zLxCks8b7ng+uF8
HiUOtefyKgMzTiMysziwAHQ0+iA/2bc5B3IwaorNMty4n1eZTxRAHJDfQc+epeVuXi1TroJcVzqc
EKVhDr532DVO5ZzY9i1u8KktjHXkEm4Wp047Ji6c/QpRiDPoGuJaoBXgLjCgvN5YkBLYmNGFZi0u
2PfYN+578BBADjH/Bx6YzCAMEYWllVbK+5tkeleUU6UZpdQxXPCOCSk0Y/3YoAJvuPLK5B4Z7+5G
Xjy0HVwuL258pSAU0hF7Wk21yJ4BTI5H7HSCSKwczZdvxuq+pspz1vl5K2bNeM+G4qelmHiHv1To
aKrC/iZ0u38TpljTE79peDZmGDsKWM+GUoy+JAwhZufGxetsJQWWoakLyeFKWD16uDCSMxdTrSC5
nA5WAGYi9NBK9AyDA3/bR5WdPiQF9+b1Jbb0lCsBxLwuZY4srGJ0XwavQs1Z/R8yn2Fxltvqp/S0
WtMNrHrzzj50G02XjHOdA8wy+hzshCXgWf9zz0KHrIv1dDgRakhWsliqu9ydnCGcRSa0brtZzR5s
y1yXYopKJHK2OiL5kCQzj4wQzqIEI2Xl64+u8NYI8DPl8d75D9+HuNG99e8yIl55ro/I8eEzhwET
R8tidvQRu1bBSaHhs93Gwi/PI9ayR36qVMuUWGFFjM/LtJuTG4Jr8G6X+wCR54z2cYupuH64u+LD
mWTbV9yafLaO7tSAsF8iX4tFcdLbHTrzQvTYYSeRlWliwx1lkaltV8Jg0ojJ4e+4IrB4SMnv9T6E
6MmwHA8PJYTp+u9KKfDy4dnwAQMkgh5rN+t/6xZucwiNbbyk4iMIpfu5vSuwtK5PC4fr+Ru51OMh
Se4DKtQFXl2F31Uwjs7YUwfbED1XwKVqg3mK73BNSUK5CcK0f9PlatXsmg65Yb1O3kq7ehIXRd5Q
Si3agAGyFml+aYD/mDUxe/w6W5z6kwKn5sXP9T5CcMvSNSFVH2parFjtOLWDiW/3EUfTg4oFB9O5
+c/KVVbpjn+TAWhHLDPwI9s5ZBl6FMLA0Faoy/LwlujOCkb2XEZVzT/R60VjuTPZlt0kjUOTpheF
MxGbowazwIWEaTp2smkOoCQY2KmoV15x9J0ZEsfrCVjC06cZpmbzMuSkjyg7LjJ3KD5z1ewOOaiu
VEvietVa85QiK8YjVgJOq+Y1htkBoNa0NSXBbiXOkq9MwnFKEVSS5YsjUXsrAWGx/mKzTa2AJOoQ
I5LCUoUdIxAU7kLEb0li7wOjE0eS75hKL92nJXOxNeVHs7MfqcfbdcKGAA04emSf7qBklQaemgfp
AgcAZAbyRkz7TRm7hclbLRGefn4Afa0A+RYJfXY3YmyE6nZ9Eq4IqEPhz8w2cI+IxWsad7n710Fd
U+HmDHmMk1WIvAphid2tuJe+Q3evYA6ITATQOhSKYaocZmH9/7PU9cQO4V0YWLaZ82cSxFW9S43i
oXfYReFQg5R+5uuGrORVRR/aAM2XiTIHlhzSFU8TKYLTHpxWz0dqoeEHM4iezhYJ9gIYLlbrYVmC
PErKIE09+SL7HnmqhVHpgjnxSY6+rdHVwBezfWQVv6WlgHXqN424gTcirDrMbJ6WU9ygyDkx0MY0
MR+vz331/Fy1GL+nGsOh1eODbE1gQ7qZuPTXawTyNf2fm128mkUpz7tTyQeZqPjUFJuhUVz/a2wL
tksmKWfvb80ZYp1sNBQMszXkSs9suPUDR/maoQKhH8vHN1802yyJDAn3zUwO7554hrIO2fxGphq1
/EfdhRhQt3AgTAHHcQhpq3kmFdII629Rz3cE6fzRk5QxQtZz4z3zDAT8miHQb0lMD91MJdwVSu11
p2i6w+utlTMb8k9YXZ7F0tvspEKD+jxvtGleaAMFD4Y7wo128KiPsWf3VPt8Z7EpXyMMhkl5/Mln
KZpnE35x6Ii3x/wZHx2zEQNOvyYAiy3LSuAhTSBPnb6FYP0e1Gz4EaT3UcfFMEM1eHO6wYbmrCuT
x2KstCug/+wH7U2bRf8fJ5hQJXuHP6D1b+gEttcMgq4ZtxEifK0a2eLvBlS/T6lSkEGe1yqcomyQ
6zD9sCtcEfpHfg4/GMl536iqhy/yN637tWYpaXgOwgRz0YGQISLvlt2PbHcht/NyaTSk4QmtdUcn
Ey0G/rTS54eVJOGsf+4U8AfGqAyYuyhTTnAEqBZG7cG7HJbx2r6Cvb7mhHHFu7Ui1k/YM4gsRitU
kCr/9N/M3rMEwMyLyVmF4C9Z87EBMImRJ/Y4OH2eBmJcGHTpA84/pbwmHjRFxl2UDx9XvcUqbsDp
WgNbIbZeL65xkltM2rYe8xzZ0U44CtFAqKatohpjOnMiHojRWi2ue4BdOn5SdHUTCDsJWFFnprk0
U+lKoLPupVD2D0vuXW2WIoFRc3+Mcaso18jHWtBgFRSypO+du2oZGmr7C2B0ryIQZ+g8GFxAbTXI
2lNcJhwSDQM9LkbCLRuLqDm/at7C9zo9I4Am+dJwMyHcz+HsgQJjQpMODCjMJHaj6wgXEgchDoct
rMxTskB3SntvE2njAGgLfIxpNb7yEZKpKKuNe7OEpTOH0qZzKB+HfJkmKlRPX/jUg5DcdzW7C5LC
MJa/922CenjtWEotPgbLI/nOj6pDUtMKztO7dIKxW2dFpbT3bGJZMcQTP14GE32LZ3aUQA8HcwbL
8AjU9jbGufmvB7WAD/mtUfzV/ePFnX0YXdmKwq8pLqGtGl8A4eY25cqsN755AZ0GC1dVImSMWumu
XjJh0i2GheazTXM/Hz/G94NmseuVkR1zwFquFBXe/UiXAUUUM7/cgUir/KIT87+kc/k8+IKDo7c3
7T/Txnuie9FYyjmfSK7E7bxTRSUNyXsjK0q7my7J4piKgyvEvSbu6nkAvLdpmcMmitD/WqRgyFD2
Kqy27Gh9EwlNo40BUN3oUgPkO/cs02hUz9iwBFP8aFUkM+KtIK30Uxtg3QsWvNRxaSEFz/A6HvF2
D9zYIe1ugRPl3TXj2fE6hwvqmO24DMFBsQG8CV+YSA7y8xMhftaVpr8jxbG3KuyqcYJBmHr23eVz
jqTFB4xII7kNxjl8yxz+BpwFYvY3nzk93mh7ZauVeSXrMV//c3eDdaHsBpcBy4lwqSkco30RnFL0
Uz+rrC2Kl65GXAB6gTEozT0cLUECHqJpY1f5aB6Hb7Z/mqDFguYTsDDdaPwHSZd3zBfehD2f3fB7
MnhifoOYFN1ksi3Ju1u7ewhioE7qK0Oo1j3s2UKJagAZQ9Fy6Tvl6LvnGaFvdWfsIkILFr/XVUGR
8pftPbASSMXBbnuglGiUmukIzHnseHlFt02uY85j9kp+SZVDydXr19wVYO/7wgjYZQbq67oSswQ5
VnndGID+ACj0Qg3cKMdXcmNwfciyoYhpB39Vo0l6CRmi+iTWJPNt4SzLG8/nnhTV/sKKHkgM+9Ua
YuQtEXdDvY253iZOdiQUziPXkaatigoMo2kI0mJzWKwzJV4oY/QWP+IMAjZFIIEpH//SqIfhe16B
l5hh30qV2NEZelb5A9w4UPQbuMJSjyqZQOh4pJbHL14HMzgsPiSWVy8rnyfAj0ioZjSk1GluWPmm
8r8/AXQkmRwFNq26R4ctfCooEvLlh05nxQZzSBHDzpm02Iu1t3qCsDalR91IJsHPqNsK4syyz5Aj
HpnE+nbaZnwLupM+DZ9QNgHwBazjt+TRi8ESUAhjUSr94JaMaVMkbvpQSBEKiRjpHwMjbBOdsl5Y
mTyLG/O/btGCOoT9QO2ONVl1NavbS4almdQoYaLG9dbI2VSlrAhuWl56AjxHQflcD5dVRL+VR3aF
hE5WN1MoqzjH7yiW2xP1DB8Udqi71J4PfkK4zE2ziDLAyvsWFM7JO+DqhQLaNzuCVvQc7XDpyXSb
1Wg/aF4pR27rTzJ37XNvZx2wgdm3RAJvKMWSNk7vGloV76ggGQ9qYnnoaZM4XQMP7s0wm5hiLDm1
ie8F2vE0Dk3A5TS4jgV/TCL7HuUU/tYc/J+wzYchvj//iIpg8idmy0bmgYSGFH9EKAGsLLXUG8vV
Hqw3YjFdYx1TqD9Jpgffbb/njBkEUYa6FoIDJJ6kNtz2NeQKZCTA6kNq4ToIgThtMGz2tnitZmUP
MbI+wrXQYUOEZhoFCZ66gwXlWnrxAaCqGjBW6aG+wTBxxTHWq2XaZnezXuJUiJHNWPZK30cuGBqz
M0yYiftVSugJpvnZcDMQxp5ch2yia1MjWZ1r0UbSgkPexmwKAr2ernwohsCv1p7ApWygeVxZ5rHJ
3lyG6vuj2V2hnoN+nprFtjLOL0WcgTZ4LogpNUiU/VGSofY50dEkKLEjxZcWhXFy7tGIDRi44KNb
i2vK7K3/vtqYPip+i9oF+nfz1WK4NlCJ5a8+ZU72ljzTJFZNhIBgpcI0W5L4e4c1TLMxotnhuZfG
xzDHqY4rPEMQxsDmF/gs/3Aw0hcKVXkVRBZ2aaMe3yMtPh03/vtDeQ2SoozLtJflTt7W35YgNk+4
bDtdJeQTRreWPpj62h0U5uQlBDS4NT5ctesYdulu+ieGknWY1tZ7NNqoU7YA0+Z25Gs0I2LU0imC
dqlaigb5YL8PDAiXi9Rif187OmNqrT+LncOp8gnNH4siW61DVBSdFmuEmOQ5Kz/MCu5ZFXea8wcN
WcU/pZw89kJg3x6fNreIo3tcueeawKEQ5uMf4DHLipDujsXauY5Z5kxONpHTvt4ELEbClM8AALCA
5mIoBHCwe648vbupkscrwYIVBv9ZantgYqS1J2s4p1HEzqZEndVJPwzAs3jnSJVmyGtcz+vdVxFT
zSRI5XK3imjLULt/dk//tCmhDh0qZ/lxj14RLP+ruYftfEhw+dZx7JEZ9RI0OnvkE8guGvPHYQw4
WIV8F7osnVgQxCSaakJiiwtaq4mv8aA6OSlwuqVzFakBUjIVIokQvFKj2mTJB8/+J2/IlMY4hhFn
guGT4iQWiVJgSp4ci0t6GJYme/AnhQSxB2BLPSa/vOWH2hZoRityu5YBOVEmpeRFdndr+aS5hhCW
NsM/OGCagYBTmSp1/lcyZG1l2a7nd2wbvhOGSKpAKcP5YU6XzZ3mZyttaJZfIMrYNIKYPC+jhMih
piuiNzFOZqWbkt4jhnMlXC9WuQsOzi0FCYE9Yv3fyl0YoQLKKKshTPkG/CBDcBLcBCuy+r3l0+Zi
JFSkeyz/gcA68a2UmZ5bMY8WTvQwy/K59EUYX7UhW5NhpEZA9eO9fbGMeolH/BetN4ed8YONskfZ
k4WuW35V5xVqFBKB5/sAh772vSEY2Xw4OhdOg+fzkp6uRpEF+U38yUDxRRpdODVUYEomRg98EBiO
SShRU2tzSVZTPNcGX95GNE9LhgzwouLUqDGG0/coWp7GmFkdoprlQvbAI4lDHVEB/axfkVlJsKYN
imzq3OCuP7IOcbdB9nc8OJleDSVRtTMQS9B0l47KD20QQN+r5RR5qQpRnok8wBgwTSR2hqYIxZno
1GjYziYEVU1chxDKrORgj7WkYk4IW1ZMLNpCZHulACVbjBJIvdld918NM5wBb9frDc5N8MXhgB01
wb8gJoP9GnUWiWk/CPvllqBDjrtI3z3SfTO5bwiUs9zv13OzM9x1cpgStDxCdYp3vsf3n8Y80Yhy
NAwdOPNIRxhWttBL420DhmksWk6NVUY1HEeB4SBwba8iFUUt6GHnTWwK7nd4p908hEiP5JdLPDrA
Cu40bWAEZvDSiKcRJxpGSezvLk7PXH2xox7Pkfl1c+0qMIdfPXKvx7N54Ol6FhBAEczD/Xhr52Fk
ltgheSCEHkrO/Z1NyEphEQm0EcnMUxbHssO/9WulsbE1Y+TSd2CzRYMJKi8JxymT6bYQpcjzEeBR
QvSKK7NWETXqaKIb1jJImHd06ZuHdwUaPJZ7tByIwwaPWAyHpp9Ppu9QGWH86ypNKsYDO7WvTYoy
PUWYqSd2Iq826FVJdt+uzs5no3e8oVXl7P9Ze5zKH6t6sSN2sKjpf9lvw+LXLU2qsxy2RLLN6o1N
aj/Ssuh7+HWvTyWoK0ix3GcTi0Hd226oCIv05lqfl1eCTuO4mYXQeKekibSeXc6PgJC6gour9wm5
xQ1sf2vKB4TQKhrVvXyKDLmD9XEIna/6HG948ftwAD9CP5zgbpue51oPR9te6wNy4q8aQ8c6ul6n
aZxKThJ5M2u6rwSu25i5450b8Jo6z0jqxo7OoN2M+aGPMWSx7QsRSojtuDynkx8HgkfaOKljynll
je7gxjhoEN1G74gHFcy1HmEaaxDnJ8LpNYpdIUlXQQxHEkXWw5TLmy7llLlOEWbfScPff5bmwGTG
6+0GHODmfBMcUcaU7I6PMBD0hULUstYt6pXKLHjB+LZThLXc6oah2wgiGOF+GrGbsQlYRnDemr3+
dnrCZm1jNIZCcX0Juj6GO4HCkHGmFTtK/VLuzz181K9iHobffJtDnKU/rlMhWiTxCT1v/pw9Leyu
6z1IZe+tbLmvXO77hUDb2xhqVoWz55HS6xDhoohs1Q9ME+L/NWNFQ3A9ijfpsijw/Fqk7/PbUuRx
BpiHvagkEhJHk1EGtu/DxmCfBSE+jl1/Z5XqBTGFkeSKjpYgdjyVMgsD2pHxnjdGF22moPe52cUR
8aMcAj7CItx/PJDxvwn3mm2qlxXLwmUAn18MgcZiZ0vwI2pBh8txrqrMKF76+6sxY3RdHdYi1ToN
XH7i4YxuJzd9XqkRKpl6CFmegiki48cLtWBQmWQHHT9Lid9mk04rb2homMRgO7LLuvVetrObRY65
0GCIWlHG3k91xgbQguTfHZ3pFszjHKJCQ9XhVNsDOoWe1mTxvYiB/TCi/xmxc3zcIHLUQvLcrVkE
dD+wnoATnCirACozlY185i0StYbOUxLE/NCKxSplT6nq0gv/L6DWgXGkAeWkdbjg/1LEyiWuLPoN
/Q8FvcDKQMsx9J86XB+yt0oqL9lvpUAwNwI+XAhdlXgyDFJ4svMqInvZhnEmjerr+38aHO6Wj4Q/
WJoCwDk/2hFulP5AkrMGkB0+zFpBLC80AlWrjwtVU8q/kzQQbcpArCGarO9RDeCkpkTFHQS60WW5
9MHmDF7jFjLajEf9L4MsEca0qKUTAKA33JRgXzdQpIkaqHtdbQqsY4KjYvb153upoomfmKZYFdpJ
gnkSpc52RyxMJ8BKh35+R6etm9rCxXcO/01HGAHKNq3BuDPSWPCeXjtDeuBPmr60w/CGjImMYu5f
qs6iObkNgk/r5PnPuPc46LrYsz6vgyRwMSCMVG37RCg0Ic8Z0ZO2cnbOjVARJY0aQkpA3cbozL2w
6yRtHD+uHG1mQkolw8ixjQm7Hc51k5nEC/J5ESr94zj0XQowAyWdGDmmKOPMxk9PNJCxFF3CoW0W
8hpWMqjH3BtC/2JzENAbFvxpwAogVOgr1kkMqKO3b+Y02PYauRded00PaXxBbJf6D2RxycDZpQm+
uNPjFcE2fe/U4Q9JD+DMfGgi8F1KNeSVH/1p/wRvGyPC5FBUzC/UV3iyJYBUD9wd8FTP403wGlMY
LOUWMxAQZndBIt7xLDzalwlfReW3WAiz5F4NVs9pYW0bzOFsQlywOTD0iIqdiRwov+NGVsEGCeXc
VKkQSC2usFwYSBDTAhJHGccpFTkt1Iu7xRBx7Qvq+UsuJjgq3WHbvkOePjxRjixqSQoKflcj9oBm
mguHzy2ezH/kfHjRtls/L/fhYLjliJpfw5UnEj1pZL183OT/UANjCpWchVBhPDdLmM0iYxAfWj4M
ZfPhAO3Ovt+vJInBFGgfQNxN/zDCOTR8b2XD3ntKZlL9BTBIlsVEmL3LrJTHPbQawrjKp2fv/lGU
M93sYT5ZvfnPyueX3dCXLCtcdPb5oj9AaPaZC/akM0IcCjo2PvFtkiURWv3Q+IEwAgwNks8oUAMH
FTvogmJxUQYI60tdGfaByVZRyXA0+zmVGpCoBLfUlSvuKJawVLxW8rZCumD0l0LaujRLGb0DgbB1
OP4XkRHHQwrvdzUBvI/rka2InnRIaX2m88WUX7rjw0HfUwocxrjlNhx8FM3/KN74l80hS5Oga9dw
q4+WsrkFqH1HWH9AFqAI+R5gNBFO9YDIWmk3BfG1iUfeA6PHYwE2j9L9KXnJsZSNQNx+aw/5sgw8
uWWplmGFUcJN0BsJugtc5tgw9rqJs7DiaYsv6NpBG9Sg5R7abykdWf7QjKs2fex55o57t98oGoa0
77e/51C2cT6ibfERgj8vpce5fbzViMBLuVMkVlpgt+edrWHDJ++rhRO5r5J3/BTSbLQ/TdFnLPWT
gL9wOMAdkuTSKrIw7XFQKFOj7aMlUmuTXjyxpTAsrpxurD5yEGm0h6padodCYCuxCP4HQjE0LqZX
wqiwwA8DBF91y2G/VkBkLrzcq+htHfh77NN0s+llMbPof/g7RVI1O3wSv4F3a3X2AHc0R4hbH8rh
yb7py+LCwxkwJNqOiQ/TzmJ97u2nJbwbsr3ryl53bhHDrr0TviaT/KXh9AbNf2X+Xyt4q+nNsorX
G5Q66pg6qDcvWmas2jmJM9gQNSFGN/CYRABx2+pXD8Nc9x4ELR2fhvfRZL6xkflyrfI4oFXsF6x1
VbZuDGIa3e6u6LKdgYPXONNvHda5tk9i2ZBI4jRgKxNG6r1XljY16i0G5it+DCddymg69UU4+cwv
ZaUARQGGtSmlklklcFFaH2hssdj0htKiCiZWD6LYvhzccBJe1jX9orYUfrb8tzaqINxGAN0IHNhS
dFEvGTdSFAGjhbJqktdPUafymn8ZH648gI3Lk4uk09lB0DWoiPxjED7QJaBiCXFRIT5F1XHi5dRi
KCcrnzUP6GEkGYEz26oaaEFog7XTAR66gVy2oaZE+uBbJMOIRF8peqn0Qlc+n9no6pBt9xSlJT+k
t3DqHw0xdG87PJNK/9FaA2hXvTq4G/A5147vZqcDBpw6CGHvuLisTGy2Gxc/k9m0B4JPYIEFkuLt
EQCwqRbtuPT449qizL327cMdFd9YxSaFQaARJE1nRynid2ZTJneNV2UhNUjIxmXCE2QmbHqgx2Ad
gH5pcXrmjr89Ot/UVTkvKjSGrPRS7VxFOUrggxLY8cdcLvKDZG8Z8PoHZi0i15ZF40z243c6EyxG
LtsKYdZn3p9tLLKPaM8mHLiU3yb/uyR63QY/YRhPDjXjPK5aS10M79f1fA/p1VLomHrRMDOtz8yP
23wLaqCLpT5vkKYlFLnvZC9SctcPb/YOxh2Hv5FPjxjqyzOrSNpGbI0q5+HtNS5J/IrYeCtJuROR
wzR+0wSaHIgsYt0YQTElH+bD6AlAUHjQR0YsEfVPAsP2hXesl1Tg/IgDAVYwkN4ZA7lOpAnMkOVH
nFR5AdoeKuWzRRRob0HwtsLAsHbBVc8wydukwRiSNnxNkqQZf/Bk2X2aguJs6ri08+UV6A+bcZYz
vV4pMnTxONqolrqnS7juEJFVpf5CBFxX9G59Paj+K6+wMhLW8MxLVy5T7OcYVrh41eoA3FpBxVY4
zx1m+jyytWMVhyrWVGJiRfYdUxEwCQ5LCt11rj97iRSoNr1K/OmDDrCs+C8eQgRb+ZaJUcLHGQUc
UgZTUzBwZhBroJiHcnwe1QuIZ/uOs3ce5mTuHoZHsZ1a+a+aFkZw8IN+trEEHI/0TdJwWwhgSqdU
EN1zUmZEpk6WMPbPC5fkQAz/sAoqLiVHio/627NymKvFS0niYCYkwfvJPcTuZ1ik8mh0Lf954gKs
yJyEYKwbPvKRjq1UduG1ahLoQ4N8Lm+w1U1zGQQS5t/uR2bk7CeGNPhqP1YENRUK4B3UfHxQRTaH
/IiiXgrT1Iyi10us6EdLs7XnZjt1GByIz5i2VpQEE5KFeye5GidJH2XNuCAACPVG1cLlcLc8rHA1
oyvGpuU2minlD1PKKolpOZgecVI6PSrij78RXzIE/Dj4oMrcdpa/43kLXBwmsnyChew6urGxhbIy
sHDb3yE/Q8u8h1ikzTisbqRxCUs9CY3+jMH+kffjrbWzv5RWWMDjIRWACgSxG/jrLcDU+HInO13l
QoczKQyQsPNLkJi1Z06XjdMueGJVGZjohcqskm/XIobYbsa7+Fg2LYPrIBz73iYwT4LcHhhxqzQT
ufF20a31zO7SEzyU7/a+fWv0H3Lww4NwRiEL6TI+XnD+acPHuCekGlazmhBBs1TaiITvorI2vXCg
rXOcEllfgbhlENdG6Uudw3GDhHO9fNtRXqlqLfVCCSTZO582KGwtR7aQZzKWeZGd+tvzqUxTS+O4
4xGE6nex9TWU+FkWCON5v4JyQzENuy4oLIFUM+V2EQtEFHowD08QwKRFqVcr5IT0uNJoXibLvdd6
+76jYuxo2FODwHvzX8V457+M20qrGWOQ/R/W9mRFk5Jo9qBLiCj6ZGcYlpV5gCjxesoQE/uW+IRe
KYuXRzdlZhURMAd/8VMr5hlQSzo/uWuPDKVpPGNLQCqjeXwyYEg+0zyx1vJzr0eL2RV4n7Zrn8S5
gzaE9Gd2pdeud6RuRASkAH/P/OeGfHn4vuRTSz2RpSckYeQlbFKtmpCdi2sz4nZnCPIkUtOsG/TX
2P0dIO3Dw2vtqqYubIJZYeG9NiSmbNKFI7rAWKZN8zX31bDyrMc47hueHpv6TbYKhiJJA6TGmYIn
RkKK+KG8JA5sfMjnmpeFflM2nusmppAy9O5igAAXGqTVcXsT7q5hMSY5+OywXep/xkPaV8gSYLah
fa0y/psXNEkvkS3mFAtoDMF9VpEkrCtek6EpidMUxKqK2yeM5mwI2A+nZNBoRUs5KdlzT3L060Qb
UaGleohyjOiT/8xGvgavufdlHcKz3BVj73togUeF7NwST7M0ZnsZ0dhkv6OOZDONmAEjueBV/k3X
gRMndEgtUoQhtvPVNGkn+oZvM1iHwiRIalJkNnOUOkJXUKg/SNW2XdpMd0u9zIUoQ6M7Ume1nFH0
QOk18WxuYBjJRzYW8/kxva7OTlAtTatMSOpPjqiwEncETS3F1JOiVuuTo9kqmbCM9JVhj3MnuGOM
7akBtqzXyySmwFs3SP920CISe6QaS7nCVYv3MWnEtHT3WUHbcoxXlBZc6YZZTG8BervZocg773YD
MAhSCYxHi+hj2+S1T3Nx1K94SJqpQyyJvmri1nMj8tYBK7+Tv++iff4c5TQjiPMxXWb0ijlgmlZm
En+fg0nviKhyp9ZB29dPaHRD50pyGvuUxzYmpahUe77VxveR1JM16OvK3xUvxuQIZl+Kga9vtVxz
pyL2y6SYjnjEAOnHWt9h87ELbfG9SaQzc3Q5A7egIGG3w4uZ6BzKUhi/+kuqal+MPc+StZ6XOjOa
C1Hq9rUhtM9rdyujUm0zMhUz+zOeHxTx8X/0qtx0fClSvBV5xgTYEEvMWLZO6A8tW8eckGcVU8Lg
lZy88tvrT0xTlgfvcH7f4psgQcH3CUHtRWLaogU51Fb2ALFK4PW1OUZpLS167eETfuKzQA8cVHnc
/Aq5/SrMJXTniuPvJKJrRNnrBtDdwhlkjPyAOsklkhXQRAWInotHGN7HEzWGc2CPGIi0+lfoGdpO
6GI6kVjtk8X4KGwu2qLvtk2ohvGrUEmTTuOmvJPWkPFyJ8kUegOANXYlY/G9JtjT+1qRDg8R4av/
6maOSxcC354IT1L+Lvtvf/1KpWqNBiGsQdwAf5qjmFuvGo8jGgOB2thikFHJ1MUxEyJeL4IrblBk
3vVgnSLGnHJM/AecMnyBW6IVR4of6sH2y2EKaRTahI2dF8TDxifkJyXv/ucE5aE+n6Lqs52RF2Yn
nHbAlCbYKojm82QJd4yu3vYsRHpzreaLKEzB+pECoCk1x9ME9eqiK73hSjedtKhHmN8xVppMmENo
QuMAZQI4EgBryMF8k8HpIsPw0roVmqeI9TSlNWd1bhckbf92giXNjkfLwKvRlHiPXtni29f5PGSO
9PbFLRhM/vBjg/ZnRfnQTZ0ixrVwczypXPJ0vU2gYgNiIzUooY3NnJxOqUjBzeAUem2KRiiWhLQc
GYxyNUnN5re51jmlaQS6UK54wZtYUoGycHvz4mgksM5hiSpkrkwFvvG66WDauHDB5FUff0wstnfR
O+MbcgeO9C/yv3MqLUWfQgMFpLeEyJQBFPwk2bGDZswOziOW59ojvGM+b3F12zO9Y0m7aPK8o47W
Rs8G4H0jpte3aYWKF7CTO6kQvm13bpiCzt2jD9UtVWvpJpdqWKfWcasPYwU0vGGeW5Pwkn+MTo3W
QWSmM2RNdjqa4qG5sUpgtazRLJDWgEqxpnlkzV/t4XZ2mxwlUTMpZx0bDlPykMAbk9TxvKEz6HNQ
JVnHMbu2ocGNvvKYgRbSRe+k6bFGPqviAR3/ulKb5FulCkXxGY1zOFAxHrDCg7vThcTsmMADfr0p
LqI0pc9hlQJWHtiOhK8OS5CA91CnbO3fU+qG9eB3gYKmb13VOHGmXq0CvXJUqUyxwcPlL/gC5jn/
4DiKRFnAcX9lIbR1DXXyeDAmflR4MVuVxClPbJNeXRVa4lm5hH7aBMnyZCQ+13tu+6XSzVujBJz2
hS41aAWRM3sREx50n0IbfozoNP8jlL1gdCM/gZDmpM5m7gl6H2jBEH09QFisrJAfwjRu25RCPcbr
kwKxboitngfeS/PMH4TtFQ6SMfJzuJ1+/5Wbev+cvl4LpKuk/dulFzFSahI8wrvDbuV7qVGuNVzd
Qm1c28+ysMRyynSbKCGo4iYvLoeXwknLkKhCvRP0vjeE9BDSY5hzGBM7GC5YLZoMdYqnVNx5sSLl
h9/DGPESAuWxvwEHXWldPKns8r6ZYoot4arKA/WUetfHjd8s9WPW6xhrW9hDpoAB/ZDIuwahAHDW
i0MA6tv7D2Ox5gRKMKQGgjfmcvoGFw7L641Dn5Zw3kjdK8hYtm7MC+JSPbLSijCLwxiGK8Sa0j/P
IYDzaWW3np+9lX9osVdEkBgly+NrRtYf8v8ht6pdR6HYCVctRcZwGgboXCyVtNfMkq8T+ZkIvL5i
efWmloO4n93ez0emooconHSZqDBqhJggVfMR+xxsLJ1SGlm5JyP6n4k2XLKofOZRBifBl9ajWQ/g
9f2LMV6HqMoqkTg1CjsrIxCchGPEuA6dFR+JaTndnePh5tA9XROD1PWVSJ9Xb/gOiiVp8TER3S2C
xYk8Mg8i2tTq1clGI5c4tmR8dySxseXe8WKB0vC37lG+besqBzXpXAHwNJAovBNpccBNNwgfA6+t
03aWjYVi6P7Z3eqmxBgVBy57cCiZIFAE7HjxcHovfZYq0umi3T0X89BcTi9fhAVQlYMOzT7dGUz9
0ssgfa8GqlS4KIobFjBKKeh+9Xr1CkwbAM9IIaSdCQ7C9Td1sjhEtkembDYmxlgzTaUY19FC4lnz
Y/5cOztMAe7XCemR1s5bhoNOflP/qjc1I+gCjE6wN8/K/xP9XaWnSKiS3Zk4jui5Q6Pa0Uo96Haa
mf6xP0/MhhOvd8ZBPaCgy9FnYcDvJ5uRLs5zTbj3TdCGXDsEUin2A92TJzsRzkfgWn4crqX+so3R
SkD7Wd1K/1zaZ9Sgx6m8x7OfxKiVzW23tZYZbwaGN1BoIuVjgqKyXNgfGDkfWrq0Kyf9QX1uyiTf
iOJltvGKZjK50ewHXJGPoR7dFaPRg1f6K1zZNRtI2ToeiWAzV6oF+fu/6uJN/fSn0y87hD2puQr6
gJJD6fgA7zbqW/noforqt2rTqI6jILo4SlVZo9SfLge9J467Zf0yLrrL1RqVg1qe42vhgJ6OiXF7
uCQ3CsfRdtIkWZpcWsJoxmV2q2Qp0gS9GIg8dty2AnwBk4kVzKBzbMTer7oO+1eaHpdgXyVp/Sj7
fBpRaQ5bwzcv7+Dhg+AagujIGkdG1gzaHlBjTcI2WuJovE23pr6VBGmUWtfT+r4ZzWWbT6yo0HBN
EUK3h6UY9POXNFaHscykhG0TehLT81aPmzkP6Zk45+uL6pMFY+KZaulk0obhsicDQhrY0mNwNQo3
6c+DUoJ8PojAIyrogU4kv2v9bTl2c9y7lB5OJN0AIn6y6INbIYvuFOyjNU3Dx6Ri+aHyexNaeKRm
Rkg6e1kMYgyZyV9EAlFd7UQ63EloDveN8lYZFY9pms7tM8HkUOpJRyMIPIPHW6JepRPfB8GH05YL
/LJUHHe/m1iqV94aUZq8YciyaviRkehCYaefQO8i9GonFjkvmzvDE5gO81vyJkWIs28TDRMtHS9/
d3xXjjPl5QTc5/RLNg9UUT332RVxgLOqYTbBxdrb16SCeJRvYQDBMHvFha49VccPTL55O03rTvlI
HMbkOTc74PiK5l4yvbKtIDBmtUWdfY7UG6jyIwx8sSlEA8YAIixdZ7NXWKcdpwyke58CwT3pc1i3
9w07G3Z05l6gmobvTpX/QslJ8b6VsneGGE7uTwYVZdq45a6fx+ae9eFMUd3tqOawY9xb2WdPUg4K
98QY3n4pTt5PiRqa3M20IIN/SjvGnJA3uNIgWvoCfcmzuJGLX6jt5450E0fU1ypQdR7Ojgy4Jo9D
qUhIK/mLHFz8vzFN+YlB8Of2/fjO8dBIcEnZ5zcNXYsxs3AubZ0pObMNgnv5rX70gHkf0+KAhl/J
StcbC7U8sgoAfzSI/SR3gQ2YliGfqt/shTrcMCRy2jDGpM7SXVMtHHgz3S+blk3vi7OxjYur2wl2
knk2OVwvqCmmiQSFaCijQTSfleCsFYUt1wxDGZmwoUFca6qoJYZuAqefNOx0KUwEy6T7kdiLSDFc
0o9JMmppFWuJNq/3b3CL+03cpwsuoAL/GIfn4y9GhxyDDhJKjE6aDbAH7QtSrRohbpIDhRYspax0
qXkogPfHh0szrwX7QM4yiHGZIRj6ESKskXH1qNl4E4nwydPu0upM4M4xcZoMCZVCILjx1WcAYtEB
VGe4ccMWK73TiF+Had2Wup4SZFRcswBDg+zymLdJoFgIudzTaT0Wcbyp9cVpi5XclOU2oWzQB91F
EaohG+zq974TObwrT47Q+iJgKYivQSreqN8tIuxR/Ee/oAwm672darBwyfQclP/vr3KNM0XqZJY6
458/RdV6VztOdhqaznUkYiWDh1c3v6dXZaSoUkBhqZdCLSQVLxMoH+o4Cmv3q+PoC4suY8qkDdGM
FfU3sJjto4Lzyp02x9RvCcf6SSd+boaMhVztqgtZJ+l26Z3F8etO70ojNDOK5NDEVKDD5o4ggLmj
NJZPzswjD9NAsFT0i6BqEL8LSN3fw/6CAy+8EcBvEV+P1HNsfTF2WgzRXX+Uc4pfiKHtlWuO01QI
kEtel8qNSV3wscUzGfWubQOQlkxw+c4z5bF+3rWAVDgn62q+2n+u7aqdS72Hk+AnJb0PRVHrw9P6
3l9k0QWhNt7iuuF3E2M3X5oLOrNPYk/ovb/YWmoXaBfdcrzxyvxAOydFhX8nOxyYgFw2EP84Ggh7
WBl2YEH0pLm3hWDj5K5RHSmzrtn4Sf6yFr0+2AGFEvjn886pvw3hOp4mOJ7piMrjqdp4qhy2NIaU
1kp9Q1AtzPn0D0cwvCr/GzPbdegaTlb1B0QRepETGJYO3qFr0LVc6NbkQ3+M/j+qb2SVF+Fn52R0
mj6Ceg4EXnNfubh/tKW3JQmhJ9ZpW4kbq0Mh3DwrwLy7h34JuZMYUfwIprL2P0csVEyiRM3/49Kk
FLZzR7LUt4AnyJ1Yb3QExFcMrk4dwJTa6Ew0YpcFZh/1ArB1SGR0y9hZBVYsSuk7fLWdYHGbCHge
Ki7FtioXIMti3yES4bPQR34NGrzWMSfczEkaigoRtBS+EHbRj/30nVrqWLsDaq0EVS3ZY4EEsLWf
p2J+I1F0ly4jrincbByDSOPaglFBP35E9ur7KTG6nNMJpt9mTMG8KjJzeSbnfSXDRlcCBxbmXX8p
v0J/B66/MXOvRzwDF+mdMABWqR6H/T9NnBqxCs2I9yM5Z9Wm2x2kt99OoCj4nXkjymbnMAE3/HqZ
uCJJFxdxbvuEOYFxqEY6x6vq5Wwuf1BmGij7lYn6R8SHS39TW9JphSIif6YBC/ncUKQlu+cym3fl
AU4Rik35tMfbI2f0bkMYSeV1i5mX5uTE0s8qF8UZYuq7E+gcWsU2jaynt5C7jpLq5EH4+5ol190m
eIme0jLbv1eJoYdOrPeKih0eA9NDPMv92jHbwgt76cmzfErcdfopzukxFc+bWrx4xex1KBgOZq64
5J2nrygAmPEfxd/y6R76S1YylpgYY61qyeV5Xo6I/HF3ohn+YhhCEPHgERdMKOSPAwjFqOB2NtFC
bweBdgwDfBHhJ/Ch+OX0HFtYaE65izDDatNAxTE09gGl8r4yIxqPvY/3eXWFbmEQiUl/yCfzjfSb
gFPhyYsjixVY4bI1Qi1ozrBBRfd28ZjxFAaefuCpOxEI5LownaALiZWyEOTGvRLN7ShDuRJhhZH7
vGOT2zDFW6nj5Ul1lsfrwFEttrbVnY2DOG6x5KZAXoiLOAV28WKtOtnFAickmYJ/BM97fdg8SNCI
xo6EkSXsVtgRh2W/+W1VajrGcrhG8q0VzA29I0rizEkq/cgRzTt794Ay8e5LHNzig9ySnmo1QA/g
ymT9RXSmVPro7Xxe601JSpPBMu4OZtOHO61D5S3AZ8HjbQXtf1Lmu2W3IPplmdRGOfA/PWF9C/zm
tmccTnaco7Q9QjS/0ceybBPMNAVl1iEo8Asqavm/JEnAc9mCJNFFfWZdkskNnNvWNUCt9cUHwyG1
svswFFLpbnvJv6WEPAwNaw2qUb6c6As8V4FwmDTWqRJRS4xrVSsKvZqFyeUSa2575Le9zFwCwu3g
eDr9LpVHkUmNcuV/7VSTU5yII0bCppeURDI3UpiECM9OYecqa/5f43bfOusg7DjZ9B27lDCZs0Y/
jVZJCR/UQOYcrMOP7Dl2CoXV45g1c7EEFpK2pW6ZfvYKMq26qGLTLGS+BRbSJD+PThT7piFfIWtL
AknO8SY+ISAmtInUUp5HdiM1khyhlG93rhSm/xBUF7mXlYUG1WJOGBoAlUeAnmC16NVip2u6k8je
zhDbdCwIIuNtFoFWT5TA6jqoG5LGX5aQaLRbzOQ3opg+aUZhnkdtboGC+fOd3CXomuwqHc+vKCsF
hbblnygMcmtukRFQZ/fDOpu7XCRYDT9ceSV0CZPvoUurNxhfs0wJOoJCs8BuGtZCDIf6Q+BQ2Uep
HDtx41LvFULOiqZQpOXy/PgrRr7qYh6lyq1vZq2cDhFxHKHnZQXY11Ru8amwiIRjOgUv8a9NIpeu
eTx6Uqcu047WZIuaNHgycZUtMLXKzQbHaC1poX/+8OAa4vBj4M9nMiCMS3xZK9zbdPxgYw7EUqdG
pxF9Uoiy48KTKU/wehTF79V3TdCbe7xh4veEtaWNKx7zEk1L2+uHgr1szPpZwQ7FYAejvSjAtpsn
4uaxZKhOZsRcW/h94NstdiUarGWpba4fON0TkCezVie025iOnBsTm7WLeDVqkcSJg3EjrjR2BhHW
y63zi1P1R0W7S3lIpKQVGx+DE9MifIQpnPoFfqDX5TA+KP5W7BKNH7h7GnQXJYAqIAtBHZ9qtSaq
7RTgGtb6NazfbicYH3vQoeGU7F6QlZgdk6c60/6FqZy2zcgkjWbGua/kmLI6DMoet2gW3yCdhCR3
FoPtWEr3e1fd0TPtQ7FQw8D5gW4ywhibVBXRltsLCmbPve4QVXFUvenTlJ+pQcAQU3MVW2cvGA+k
um6jvN64ji5iR79PaHaDjm2VBk2UGOJNI3pLms4SW5jwUqO2u8cNY71qgdsNbpcqNzS99lwYgDoT
28/ojBkxeRiaNu1waqWUI5EWilnInnI0hbFEDZvH/twzTssmU5WJyfqlbFnHUBESgCukQgOgzH9h
dPZICX1hRNROSM9RIIU6Asgd/4jwNbQXj6V3OHQDf0utvLEAAEX44nqC6ZcD2C0tNK7GteAgM2rL
waj1dUb0I0fKdRS4H6XTNXKml5jKlppZXlQn42x4bTD1PP++HjA0Oa1V/26RsjoW+Q+QMeiJ2tn0
a+InYi0tTZJcSSNwxJ9ziRaaHY1+CQ1YqgRkY7zYhGHr/xjMPnRFa2yTs6NfgQiZxeHvev58DBWt
gOdzGyRuEXCcbTMOHwihcxAS3vKaExrT+L+8jcCQCHQwt4UuRy9LakGTP3dmDxDCP/xkrHQQYTSy
I4fVZFNH7E+OEreeOKQivZJ9tCcm/PErbPcYItlTR35RL2gOX+BjNaJ/66+sFCkKonK5nmBPjz0n
jWvelVuVC/pLiIS+n71rM1pYtzfDRBOrLX1+L9uXtaV80ZWNoJx7GDUaB0ehY8zsc+AkYSS3sMBQ
Lv3CF4YWQmq+OjU/bFooQ2pDSCjnvCU43ztCqXvCVbzoN33jkCvX6KgmTpTwzMeqUdJsgs97Mr+G
5TCfTQRESJIrrbxupGND51lSmAUIy8vsnsl7XtiFjB8WLCBwRW/XYhWabnH+3KdxwOy5W//w+eVW
GxaNH/VAQ5X+IGEzO8f+o7d6nL8LbTkFv7fzzMVheQZH2Er34MZn3KxG++xMaoFAvVoHE+A8ezz4
saLcUz4xm2pMX9Mdjt/UbhB0AlHmQu9ZBchogOUCsxVovfUOqhOyruz+KlnLurV8gXWzrzMaGDBe
/tg2sOKATWtQU51AksEvVkznk8GECI5tlLvq9yaFlVj1P+cnwB0m79Oq0Kd4GX53YalYyRfGr06F
ZVU4l7JIN7DFeEjMaxT3reOHSZQy0nEVXust3cKVzxtLW7RQNPdndZ8y49ZfFE1UaC7tE6kUEGB9
yLa97oZyQ1blxzWSNHvh7axCT+N1a3EWyWoVhBxgHTQaT2NNkfD32u6VHoGgsAntg73RFdBgi1AE
xi4x9d/XZH7raFKUc9NC15nhi7VRoKuHCPVPvJvMy+9tRUhpp+5sF0eCJ8oE49P6SxpvJyGxFTUm
tmGuvnf8lyDLnC0LHbPeIcDabN5u/zG3nIQzqnjgUiQ9gI9olGvNiA2ZxJ8XbXOccB4XwbzVH+tL
phn3KAqgWOuwqTJTAlRphNTkl8a0OymIlXZYAtJsHtnxE+fvCVPs3ssCXKQlDVA5vDvNcdJCN6eR
8H0XXQKIDIqZpmkcNYuJKjdXwjNf6Skw+cyfka4kc+bebVHYmWGtuHL1Ku1wQVuUBos0mRQ5Nii/
7WyXQaw/qqajuckK0Cy/Kxd32WVJp5pSsCJcX4BzRexLNH0le0yMpC8sNISvFNEI3vTzQ2ZyrbUN
WU1HK1yUiSnUr7Tm0emZ33G3awyAg3ftfrv0zZBAZBaddC00snqTqnOLUdW8+hBnNWgQJhDiTGov
SOk1r/UTv+/95adXVjbHv73qstnreyf9U5pf3pX4HO8Yhn6qVHLE7kq7RfLD06lkrUYSqRLqImN6
SVE0zN9V0x1suKBUW7AEJZnU06lnzpBrH+HdrVg5nFXw9bAw5T+VJg+gI6bllREfubk5bIUKffrI
nwXrFHti2+gIHLHs+Br1pFg+iJzWYR9pMgLKAtq4iI6/Bio1xYfbnMEyBAxAEobCU2N0eNsCQnBJ
736t3vzXFgfwotBKiO6cHdZ5j0+4LW7M6osPZLOcJh6PQf1+etLdiDGFiZyh6UnECo+gyRTgJ5KS
FZRbZLikIVQN2Mf5CCydEn8Mzp3iKecbuOMU06OOyFllNi9fm3GG4cFgmAu0lOJKvv7nO2QBgN8v
CnnASY4N6tg3bEHgcRrid4qK0FVicuvvP6SBFGI3K0C5UDNJtXPVFaKbKd7zQGjiupRsz4GD9YZ+
rrwu2OHbSgG28Mo8CzMoF3nQmKaXCmHr7oWiDes+o3rRIZf263oJwqvi+29g7bwOTrBoqpJMEbXP
KbuFfcwk4P9MqqP7S1CjRhX1MvE91tQ2Mam6RSl0gWICD2Hv+/w96fd16YaN97YpyRXcwhrpWdsL
N0a/mZBL7U8WMCJTiHwlwBzx/Nr7nUfPSJQUtqwJ6XxQHOIUvsufPfpKZ3PH7QgmrBNzBSwhUWI/
FEaH9WhjQRACJuLJfMWeouI/wNPyd52BIgwsWFvzu+rWr2Rumf/p0fnarj8pkUhf0epl+ySkaMKL
T9PgpgQY1069BICS7HSw/VRwlGmc8BFMh78JcujjXP1840x+ZZcWnmrs5+jibDydY6xW05xoAOlO
iqkH+qxGYpHVQpiN/EowZu/U/WqfEY/eNLX1sSYg4kxRMUPCUbBjy5IeRQVd37RmjO5THtcJs3ii
iQ3DLdYfovrfvyk4CI2TrjZ/kyE0im6StNHUg77OBITkPGcJ9e9PXJuIco/65YATVMY3IMNHmwgF
aQYt0DmEze89kLvLIxvIS12JyXslkR8vz4JTdkmhE18bwkut+entIFqPoHBOkP3qxYLs+Az4rttv
N2LGUcsVy2MStE3uAm6z9T2lCRAyBUMVHcyJNUPPupJmyJ8f48ElJ6E8/QwNd1WEMLlCzy+p2QYy
zHkcbxGx1tUkmZ8aFFkF47NeXWpz/fr5/quqQyIEVOuWf1Lb5qG3Un4hNHttIEfkhlWbtrH1NYZI
ylKsxPoEjZ/CVcU/dEOzZroD+A9CE0dnJEQUhhqTr9X1iOtf5R8f1ro+XUSOPr+JP4hez6BAve52
pg7owbpcwGeQ8FvmsAFFg25ZIVXhSlRQGki1AYpf6159jEWKBw1U+mkmapj/B4FHdaMLKujiPaQp
+pC3wfm4VL/SNWq8YIzLXVdtGc42dd3/RD5kh+/GffIQZCNTltkZ/BfMPttpddLCHBYAuwORX1aC
6kQ5Mwnqg86lUru/vquGEfTCvjnZY7SmU80nwBRPhoUR2UUevFvtUNR4EDI4KmoccAkfoFnW04Tf
d6WwnRKsQkYwN0Wt0fRlYSh43MNSCtDpxNXgtvYx5isTe/WgRF7jUYhx2rBpouaHXce52e4y6f5X
FEAGvC8A/6r0dWsAjDMxsPTe81oEYsJ/9KuyE62jSOWoT31XAmyxvPIoyvs3dbE4eKRK+dvCm1XP
s/YOfYG4iNMr2NLnL2/n1Sup57n2mUYeJYURX0nY/xkcPG9dPKQcEzwh8XLpyW5NXy2xrHbKpYrU
CDkARUt057xb6c1HiO0rcMRfQBDIGCN+EEXfYGIofIl789K0yTu/04NIeVAK3nRaNpDnxzL8ZS8w
XTpschpJH7s9O4nGxYsfBf8G7YF2BrURsr7iqQoa8AynNw1uR1JWLhOUHO93G05r+zLQjDLothSx
APkGPh0CAwIGu/bImU/3a7PrpcmBWIbHapvX0sqv3nk/4ae/XTbk/hUO02FCpNHzDkoJVM5Bfo0N
cjLMQzgKqNhEVorPv0V/4I8/iOjSZcrvpnC3oAvLsC0nmXD3xCFRefTS8uYtl5B+o20RVFu+B8RG
j+Fybo86z/RyMgj0h+5YJHxfQA1I1zV53CF+TPHJEmb90ar65Uc3O+4VmTWCsY54KvB2ot54LQP9
xN7MyJ2fPIWVI9boHVkt/VlaJM1VJTtI1eOCy6Uh0+PKj84/vIaMO4NXUUqGoXKfPYlJVyZ2FjUO
jQXJOLLS+HIxF8Gap96Gl6Iymbf0fM3BB612rhzcFwqjx+IKwMpkD/4hCmdZrE8zC5sq4MSHBusM
YgIOIN1uoAtGvmEcnWXTOyLKtBkcUlyfL3Mgrn8JqyCm26EJV4qSR98tqSZDsxjQJNbZqOCaq5Aq
9OjnIlpnUBhOtLleQ3VZ1HlcuT1Gp/KA9+4IRiMkSUXBVbdtbIBk2vrfWUqmrersGWQ43dbGeE6X
PkqwIRt3101aQ3T5FKE89WOd+rNfaVGZJSIFQhalWz9/s+JOEQ3zUCZ8t1YWB01GhQKHhJqDK+S3
f0rcsa9111UAJllNEcqCuqK7rC16m7aC8Q/CmH1PBsoD7CXC7o0IYoybNJaqXSCpz7BKiXwwIgOX
FOhZXWLG5KAYOmayCjj9nIUYZ0gCOleXWUwQPbc30/AyPK5sfm4e0gFTnv96n1IsV/ml4j1ydSaD
s5B5Qnx0Fo3saHBj6Ma6wDL1jMS/VpezOIQtJS7om+L5QQIj7Pj8ZxEXcpBHrIJz8LzdNemHaXjV
Vd6M+aGxVcvlqIGlD22OCiGqEu6e+a9n2cCn9DGdqIqZjtsRH0KIgjU0KVlQW6NMCtk6jCYHja/h
XFJuaxfpPGdem0MaDJEMoAmxZi+XGaTiS8FETKyl1rrLZrIt1KHDWDXJm0rY0qlWpb5mmKj9KEDW
LllpGoZfTWrM5pZhyvZXLW5Aid8kPyM0oUd/K6dY+ynsjbPWycz9QPFum1J9Sl3bKDUnxhD5H7hD
fGBS7Zpi7j4HHqJqdFhcIyQzLrhldFypMG5zwtAslMx+PwqeIOALkbgbgBmy3q4T/AAGRwDtLMTS
wszf86zQqwb7Bqxh0Yni/qcAL+HC64AWdxpko1awL8lXnt37zS/O10HerZ4CyZiMHslACdkOaVOB
i+2FpMBQKekk+bdJuGHgL2p11lNWNG8sd3hkpFrxRsAmfFvZ/Lk0eYnWFLZOzl8v5MfP/Oa71BBb
wwQluP5lhCo+pbW+9Yo01LPVevTzEM1pjVNBMPYUJVtgsLZltCAfseME8y3TEcpvKfGNxFQO8mfc
yqvm6b0hkERXQ2MdQdjs2t8ZxOdo/rETmBnKIUrc3pdyWDasEevy++cRvkTuWIEgomamCuvS4kM4
nwxaNeCdXriMVPuzt3oQIdXdjc1UpUOZfvwY5lY4HMYfxRuJPzKURY2HFWbLdxQnRwASy3sNxCIY
PugyJCgc4VFoz/znwAh6I8X/Y91r3WKY6rWBmFCz6E79eiYQlcyAlFeC7kip5xduQWwvWaiQQIRn
CSnEVCIzoAlaACVQ5pkavZCIfFdK8YhDWxLRbhKKIdpTTQqHBAWgRYAkn4uMOkB+eSZYzC3/USKE
wMyqJQ4y25hMVpZ5+tmMpmKSBC7ezylwqq3W6JtL7ngLTjbJqHqQCuJ9ChxjV1CWg5OcLN5+E0nR
KXHjzKvFSxa54ZySK32vRfDJWbBN2OkKrtFJxTn/6LsDRGwXWabd9v/txfc18MzX5SM+eudXvFTr
DamsrEIryVV49eSt0UDijdp8YuiEDfiP29MR3GhpMakPQhAd7RgznVxUfr/7hzMmKAZnmeEhI5i2
yMek+GVjnCyUw33mFdokFHOolU2+Kh4MioIs1X/bIx/JBZwstEKdXNW9jJ/WRaUwZaV97tQhLrRb
z1SoVFWR6PHb7KtAl1vG+bclfhidLskUYbERQ+OddeB7s48aBUpwwDxVGjKx4DUhfvvIUTz7vQUF
//R0AX+U6K0VdKSsy7bRMo/QPWNSIV8SkC/3ntHZlzVbAG13QSFBYrm2kBkFttKXN2Z+aHCHiY7+
cLpP0B/bJX+ndGj2tiBmDLgqabsTpBevXjsKiY6zP4ya4bZ5EajAEWIkpfu4mttCyublrnNY336H
bUYHAM9vrZbY0vEfAL9kI4tKEsWbFNmfrg1XWZxnwB56BHZ7C+QQkufYl4djaLXr7UkM396D79zj
/LcbxFaTvbYO+VPkx4Lg3oEayEIhdDxT4cGx2TN4xHXc+sjndubD0eBu2vxDvB9vUYpZEv6Iscmh
4MRa5rQXD9y3CF41Osef5ebRRILxH7rcmZDaV9pCrUNe8WjN76t5ZKYslyIqciCSYbAXnfqj8pwu
gg882ut7S+uOCP1MslS3x5DG3Yws1sgyaKkSg85ZQlFlsUBKB30Jx2Kcgo/Q839YEiPe7dLKrdEZ
IFAnDda2ErSogvnx0ekXBbFCJ/IHtMLqgFQmKFofsLTvOVJanaEgrIuJxlnqFPJGqoQumndt/OQX
d7V/kraVI1O9WvQI4zyZQhqxh/GuV4kWZdAJCqtCrdwWX95fvR8o35HJxiYMIoj2DwQxyslWauX4
1mPdNgEy9bM85g2ozOmw66mDZehW1XCCmLnbnOFzalSb21pIjJn5wxI/Z0dkVBoHxKjA9GLPMMto
of3mKa1N50mdz2lLkVYsvfyuueWpAhsMVqV0vzAzI8KsCBOAxIX62lnChG5ZspovbhW7/tMzgRCS
ORyR+X0uYwTF4SCldu3gQ5Daj1hfWBvcpUL0Ts/Bs6X77/ViCRi8VDW/bGMd4xIBC4kEFhgjcn9a
zCyj7i6WA6QiHpcDFy2Qi/xviaQOI84+92lkuTSi2D0VbaOS37TxJVV7cm9jNCPi4abrglDL+Rys
VGTwCOYripRehnaBwiAoqSK2BM+yNopZAsajw3cAgYKVdBY+L3YC5p3MizpHsFEwCj4FfS78sX8V
+rmkWfwAHLvtoXRBlahW8a2SFc8jZOpeO7XAZtlsQXOEs/bEvGo/Ly640FBsil/6AwK2einageqa
6W12VJ30WSsdmeDJcdI7vbT1UG0F9rnnqfenivRG1bupDJTvH+uFyDxDvQ+VBeHRm9RNtUK2qKu0
GrJRQyv61PJUIbFsI0XTa5QKyG3CVR6p814I5UXYuox8Xv9693DM5GttUZbKiddnTV9XXo1waEcF
OnVCl9u7bzfc5jkP6i3dOGb6heMSvTyNEj0fyeb6hQB02HVSwFYhGmbTvTUU57Du42676dnoVAVA
dgeESJDfjwmDnRPGzA0k+pq4J4ojTOA81pTV4Phux4AppEqVL2LAB6gLmmIsVTcOXbINZBxG4OJ9
rl/DWyvbwULNZ6JsQa30yDEzjSyUtrOw0Pzs6Kqp1TetVtfzA/stX8hEO+ix06erbGh2NSqjsBg6
CpwDNGNex0DDW667YX9wLqAM6cfHfxpZvVTI/QmwUj3lbbMxglRZ1zAyTsikQI85sfYSF38IheV4
PsY/Tm6AkFe6JDMAqG/filvtfwL3ILcZMzJ7zRI6yCaO1zy2Aivk+KQM0DWxBKrCJkbqKKkJ4lia
LvLdrIgGEuojRF3gTJFhFqCIiDu/qu+/hVc9OsTimCpsY0SxHMHoomKeEVycS0vMJncyaJx25swt
tP4Dnh796I4U0+tYTqWxW5Uz/ViN9HjdycBIMMSDcSII905r08L7l6/N2rR4y5v2dOIz/bclJv/x
6pt1XKpvjMMNZxGV4rwu8Qs9DsCSOLWRzQ0OIoQAnpLLeeve1dWnYMXprS6MB7mU8ToG25nz3fod
z6H4jHriOU/8G1jSsF3fTVIvnA3T2kh0IOz3ui+dSCtlwSBpnuDC6Dn2bdSLp3HzvTQR7FATGJpB
ToAyy9T0OgsIi3xVbijZ50ZAZk+3cH6NTPaQ7QPMT2hzVrYG+29GEb1ydTjodne9/rZeF5RMz2XY
NuKrrJoY+zEDPNwAN5yBp+7xyrcmjOZfkyC7AOEgVbKtUpzOWEFe/ZDlfJmhny0/xlJZjlmJcocw
eTInwqhNSw41PPaN37GxoQupw9YPHnN/fOMIawT0vt9lHCobR104rhIhgVw+3aaud7SWn6eH5d62
3TFxK6R028VeqTgljJIZVBu7iuSvtW9vImehcmtqBTqufjgr9qs3f3xWTE69X4J/OXggHElb0v3O
Ft10GbjXsSn2WljTY+X2Tmz1XhOz2pGSwxssOcYtFtAHpef3WgPpBzQVaZaJVmbwbgPw639kYqGv
E9rpj0zixbfDpOOa437SCBxYBz+HcCyuyDNJjk6KaOpZ3CpYPNltfuhiApYj2V9gSJcyYJ74p3x8
hDiw4CQkM9mEciFpjjo6/hmJVHDDvu1vbrChaDm2XqtYLlqr85SRHEQXWMt/owJTNSHmhRPQs0QX
FO41pHQ95otNrGbA8ZqsjIvwBUYIEgNFq1iwZ5/W+4f8LKFjsicPEEKe8EuAWI7m06iBa7oHiiow
7ptwGgXCeg8eNnV/KXjhJuuZEx60R7hcF/kIlRv6MAmYCm0XPxslJ/nqhrA2RlJZBWjWUgjX5b3S
njwsehCGdo91Z/ui0nSd++uyqkC71S4gj6pY4j2M5UIO1DKke3AutNLLLtUeuDy6P2P+di2i5p17
apyQBLf2/pDXyQs/YuHGndN8O6hfNaRSNqK6HOFFiwB5YsDBncItq086iT7E3fBRqaoUKUqjvQmm
3887av1cUKZfwolW4hAb0xOaTVFLsHQ5NW1nT54kLgwWtqOSonQIXQbyAukaYBCSLzYh8802MqM5
ykJPq9ptyZWMiLQDxISw+B9XKlz/F2u/VRUk7AGb1VyPUNvZmOA863GD6ViJ+c56r+IqVWoQJpzW
ahequmRvvF/ZSw3yKl32qavlxvSsyHC4gPOP9F/u+o5+MIT1mVokxmVgVdxtyfsnpTGiXW4tH2Qm
Hmq7oquvHVKw8Sagvi9qKSIQFBAfunovdOOwMg2dCGmQgPw43LcwZqWUH7XB75xPuc6YhVV2TORR
1w0KbFPHfGJfnm93HrmkWh31kEb8AnKJvcfZ7Y0ICA8KBU3vmLPt12Cr2qBluhfpvfsjvTaZEZeX
C+sPWNDH8ahHQVkjJ198ZJ6PiNhzl5gaqwrnhngFpYzZaXyagPL3bz/x4yLZ5vO5lywZIu+B7GQn
0m9+ZK5IjxajN854WYRtwsM95PGd6ICLryvOhWOTjOHCwbD3jL1eHFkYOGXGtjLkw5ZLkRLzCITD
yqUptP+hjCqEB9f8tY6e+JNJVmoqKSfOqq7/7p+G0SCOdAENYrw/kenH/JgwiGih5zuHCaQtop+e
9jsaFV9UVwgZDyQos34W/46v/KKuv0u4x3o5oc0IFeP9i7DL79PXye7zOzIAbPXVZfkO6uWpgcpr
MA5PeidLPdJKpIPb2oRTXslBdtf5cAZ3o7y6oVPiCQjdbVyGtkLYB9gCwUn4HrwZMHdnNEDULird
eU0i/+JTteBLCSdZgWaAkCLuDTBJjKTFHp0BBNxcEyiTtQXQxwoAQvypq3yGr383v/mBm4pAaybi
ykFFPQVW07O8ZPNzq/qgnBax4YXFUN6CkbCkXTVsaMiwx9uhDSqy7EV8ypsscRV4md4mNINSVwe6
ZJDmHwZv0Q47cYbW8KyVjf4xVM1Rz6/fdeDx3+LpSxybtt9Ysz+d2Z6PqV4Hh/H46ofdPnPu0y0T
KOU+hi0z6DEW7fg8y0JZqYxJlPFb1naIwlFOLUV6L85+zszfYtabJHcgoQuOM6NdaXBGW+n+X9Fl
pgBHvEelcmoZ7XnHTOGGj0xpTXrqgOPqcEeKvG5Oc8CUpLHJT2ar5VDdEFNVU4MGgHciljS6Erll
Cj8ZiZHcUMosuRy8DfGmn+cErTvBpNWGavYNQxQdXzdZybztB28+MaDVXkFjRKgUSafZPVdIS+v3
YC7IBvm1Wviok1qxfpsFsGVtgi3X0rULlwe65Z9C9cDclE2SZsTGBQSjplgl2K3+NKsulRTzbwD1
/Yv1vCUElZYLGuswC5T0XpPfCvzuF019uOGkT8Q3iAR1iKuiAgou/hwpoilvmNVaqy7Z/w5T20rR
c1gtTbux5addtmzT0SGZ2YTe7/udBroS4eyx7QL4Ld4MvRx6JD/qYq2JPuCswAUWSjs6GPd9El8t
r8hNrmQ/ofo4CpTpfm4v4fkrSC3qavY+grnvyksJkvIhz0K+0hRiMdAZTQB3yibq5QZKmALOGpED
/AC4lyu/XrJ32ei9Atdrdd87xzrwQ4FRBQ6FlyjqHeHqzcC9j99tYanB2b1P0mlQE5nVlIlSrdxu
sBgqBivsx6NhO92NC0f7/bVajMjIlMiiCcg9gCgYpqWge4FzJ10wl8Wk/Jwj+TcV8U/oscdjMYfO
yb5RGRGjDLlD2PVpwf60jwDaEYZPAgVlKsPiY/ZNBpoIpLYrRjnNHXmFONHL+C1jPo4I/gyLVNbF
7TKlKJSw6YRb1tedHlT57LwqxfmAFb5GxTBKmCPiUnChA1L9NioMVH5gw5k+rWtt8w4Q0f+w6f5U
Sib+8TTZ9tqCOdTdwKmRvhodKCBMTOGGEiTsMQWCqY6gjo5Xp1PSr+Qy9FUfUyAlEW9TfwFbzTDG
VZEJj9ftdqn5gkhnuM9tXOcNU6+NL6sLyPBts72vt5YjccH5WcdIy99sKWUZqipdJ4XXgSaRf3zZ
1LCWR5VUuVqn3ioZ4AASdjkN1C7ccDrrE80Te+nzfI0qKEPFpOE/1TfSb3mq9KhbKqQKCaNrHuqL
acVpxHaO2oMA1oJh7/4wAk6XL7hHp44O5496YIyAkH6XJSI5KJe94j2tL2vdA51a9PAlSt+0GtlO
egX5+zE8FBJVAfGop758vCaJg3Ep0jXrAOYdQWvitUEIPvom4OEMwOOTROhc4BF+H1NQVR4zL0my
CK4B1zrhTtYW40WWULu2zZbzoykYnKRMBE+gdfxZ+nVEAFkC2C7ZhjV48N4k1wFO9OaoDD3He21S
legOXnstEcYmEyjpC1mAu4c1JHOhPutZF08lMvSV5hCDD1WDnfrzQ4wgh6Hz5BT+9zU3pokyTXOf
ptYIHZmq0EsEKUp7nG+8P5E8hRQxNDjDUEM4uMzXo1CdcI6Z/6BWeYn7Jp3NqGSQ9u/Q8/voH5qY
UlaqwzU+X2jiBQxvmTPPzVHH2vX4lTEVGwf2VFxIaAoh++yqlgR0ooiaOvIpMVuVri0A6tO+d2Ds
AQT0hDPI55Miw+LHPIuKTvloAhEsxSrG1WiCTHgNoCLKSPnvXg2JqvIfi5i71pPpoFoKvXuureHG
8chsC9+l4Gxro/uavurUq4RLiFZk3OIjok4ZVFgwjctCalhyP6DSHIQOSrDQkJNzvx4iSNGQnURT
69Sg5xOsJxy5cyLOM3/fbpr8ADR598zZ+BvJij/ddLvlRUfVxBfi9wAd7uUhCTs/x7FhOn3a0eit
e1EcdrTpXdCXxYKIx396v7gYkn0uRRhXyByPa6FWZ3ADOkxjfaqfFkvqyBYdKgs1B7TTM0FbdMYF
5qnLWBt9YIhZQySGftUBusNKxRSzPMqQKOIRAm7LUt3tfGmpoKHNUCox5qd10aaKHBqU0qj+UVzR
r4U47+kuqUZ3BdJYh8TkzOfOx4yh/ZcH4GXocz/YXwojY+FBMhD/4SRsxkdCZPjJYMcpbe0pd//R
G4bKjD3R6O0vFxH75u2DgeWUI+NjbGl40mjkrDrOCvMHN337XeR2ZQj9BDC4FKWygGm1Iz1brnsQ
gG0HuN6bPUz8Y8uAdPTY/qL51CHvHf4BLxBq1v0oDvmfc/xv9+b/u1hbclQ4wsnJL+yNRwn7MU1w
7YL68KrGrz9d7IeKcPFju/uyiC9uBrTCan+HAv8mO1uPyL4z2J4HSaSKHPqBUKCMP7LNEeohxmYA
CD5OydqWWqIicwcSt2seuMr+JuDo3HzlD5qOa/v0Mam5uEvV267HxHbEqUkksHoXYhazjx950xQE
I6GIlqlBxZOmjtNXLjY7WwQ4SSERlU8sa1UvH1ekCpeadoSrAUpvYbGR4JeKjs8gyup1QVYxRXBR
goIP2mQBahrawuVxXICGZdGQnHcvECCWJpPqAWMIiw1cIT0BBJEvubD4RR/41XHu3RSe6pQsYwZ+
jthfi2yq/6iZw2Hx+/MttmBIytNC8kFSahLfUjTEbR8n3hBvce2tCSW7rkRNegksdm6lWntEBS2Q
yUym387K+opOoPIIS3p7OnCrjrfSGJadKjtvmM9yJXxjGbxedNvHV+ZpUhIqJIsEop54lqFcuG4y
BU6+oC708DpkzLS8mv3GCDxptmVPhvjSq/Gn10zdquFFVE+yjdbnnLZswYP2Cv7X2OAmPz+h7iNK
Dmx9wijgf36gcwdQZY3vTaWQEK1C0jO7FigfCBKg4QVSP5YT2qsQetBMQqo58PN5i/7oC7vyoKp1
uDVRhwcMqzRxTLHcsY9jckolpv+JwBQGlmyb4tkHjkvK9WsFGMeGb/9Ms06DqtFLk7X6Yq8aKkA6
dCrHk7XrdW5WedawubgfZEgQFCM60SWrDrTXQPgc28fBsrXjJa8Pp3+aE5FNVPR15sWm9tRy1c1h
X+f60XqV3gaPxa+UjoT6/a58pEM0cBVVOUG/2PgJBjieOjztkBWAU8jXx6N3fgL1c3SowCAxgSC0
DgsYjEVhR7ay9z6Qvth9wt+m73v1oDXpHuC/Kt1CT+OqjXv8kXbGtsvoNQEyxJScMeNr5UeCznXY
LgRWyo7kYgC99Hm7CuD5Yh6RZBz65jOIjASe6WBHZIkNnbXRjn7/gD8vbknEhEgJcn7ryaHf1w6j
iRUrG9imBeK2/Kfe3+x41OXXL+JFk/MsmsL8+9ihgjUl6j4FHCwMrz4vKDPEzLrkIYr/mURNA+fV
wwbEXilY3nX3srAC+ENpsPfBJyWmO+Dt6QZAU1iry8dEuV/EafyAD3Ac22ngditb8vaet8spHLTs
H37+63LjckBAO3gjrR90s5ylP/8hsViLrjLmA9hvZb0Dx/I0Hi/BVMD0dA95Zdx8zLDv3jqI6i+y
lh9wL1KXnFh7fj6w51y+DATDldu2/GDYIyqFxkZ7Qn+Xt5TgHCcBp/AM+QcQmxyasXqrq1mOYevl
ul7A+xgebVoiFQ++r6cvgIBl8kx4Mm6zLgYd1kRT6ozxXqt0ISH5NBGxNudaC5oKy5rD5PVJ4YpD
mPI0FMGBE06ystY2S0yADviHFmjkRu3ZjdH6RNboc8hxZ7DZPgBEOO6IJeOYC/XRy89yvANSCxuU
UL4ZeHurIO86IzE39M6mQeq3i1LI8YI6//iXuvokCw/WVAr8BC6OMKCezuc67YV+R88Vh92G5r7n
9/REzRgQV1H61faBvfyA35ijwkD167N10TsZ0igAQ4/rbKdy0YyvCmgJNEx97AFW5j7PU5FlFvha
lUXJ316njS8D0R71nXMimV32xYHC2GXmzRZs2qXWheXpESEPgDjpNeCMa4HZD5dOaRnTpoPfTtqh
TwfbzbkWq49+lzi7+7ICbzjy2iDJj8cuVdaKVJS6p8R6QUyasHWxNiD0ToDZ+LJliigs8WwpUX1C
veqf1QEAqh/01XeVlXxt8PGJKmJKLW7ePAXURfI/NRSY9SrSJFdUKlSxM/5HHxowpfjCZuJyXkv0
iosSodkbUNPggIPS0Azx/oGCAnJAK243pKky8EOFCQa4gRRqN3QUpl9fIHtLrUgVBEt+uKbg8APB
FREOs0Eigh91Rr74OIq0KvtcXs3LfLSoxToTHsSxsH+RN3+iz1rpTZdZFQnIuWMibYPPuY9aQU74
L72EqwKwGkPkxGw8+OLvKbV9ylfSvb9WDHSbhN6h55vxg53O7v9Gu+ODqOjYdHF/o9kFrm3DPiF0
TyusVqzQgJhfBuzQ7IU+DxmZLdRfnmuOsV215zcnasK0B2OiTrjIouzIAzMWzOyMvNZy0R1F5VHp
uAf2CoI+u+Tx3otemWbBrHZrfdthedFAC/0QSEzBVcvqrC5YNfliHcwQyea+iqBPsEirFhNCawaZ
WSJeLHVtV76KCRfv2LX0kZRGxIMDW9Ey78WkRRJv/rQnmi+u2MfNoVzbpOhoG2FXyepidRZHTqjE
L1EzFoJ6fEPS0kO5U+t4x609mFgtjRNxU1EoGUnZtrfRqitqxuTk+kW2mxPWrpwAIfEVhSqUtpOp
L+fFDw8zm6HdoN3wScq/lfb7EAzPcd8cEegIxau+02IbJt4J+7WEtl1E75+ZGqXu7Ai7tVhJzBFl
+wDFrese4Qm1BMXfWXb8p9Kexbj82ce8EEhq47ujh30lgx/oV5lnuDhURNTigVDdlFnpmXvMzebo
wee5F3dDVC4lMkRHQCiWGO8aDEYiu7RvX5EvOyRlRlxtb81UneGzQX6GmhicRrFiCyDexi5wHEZH
+RqelOrBowyPC/FuXcFoWP6wb/pWhKKNTVGo0bd/eQSZCdXw1BYSPcHxQ8m2aUkQrjCF3Qg5jofp
vC1yT+uV6huYJYEuHC259RZ8H6UShdPkfOgt+/Z+JvKPRkjOseuDvIQ+YBFiqRrLLC6g97olKDdU
CAU63+ay6D7bohYd6OFc0Oo3tTc1fkG7U2xsNA/8fMqsBoIoEajvlu5JkxWemAjQ95deT6Dp6QI2
ZWVluHQCc4uxPSsmzjO9Sn92EwVgUPrPV2Vyppgpjsq7AzSFvOuMf/HOzr9Jnz6Cj1th/+l/mtu8
aSST0GzjYAx3NrAQs0WYpryA30CoDylfELDHDtWiG6dm2sFxzj9FVRVMZzygutwhYTszU3FBfTgL
Zqxa8Wa68o5yNSV3OZdnPA5LB1yeS1nX29SY3mEZD6fOafMkz93BiTCV3iHq2KT23iwO4VhxY5Up
fKCDQh9Z3axmO84eM/QBqCIwX3RRXCru09MZ6+tQ4FjXyOquKLF2FH/CyQGdUYYJSTeoih5Wtkpz
M6BIYvGoXwqImdRGoCeoY1m6vURartbLZSaPsCbyjIMqgp002NL4cHd/mIefoC/24gnCVrG+0RIs
azodwRCz/3PU73I5R4ErYWfspwZuwvD+B6JSsYOhcRDVyafm2077Dy36yu+K509VBO5GOSO5ndr/
hXVihUOhGIdUCxfMyZOvNni0LPCbY20DRVulvzowzXIygkmJ/cAmpt30ceybCQADe4Jou71+Jdss
wzL4r25rMkly7QAsMmDCVESHM5vfqy3Vhdl0qS2+HSjH05vJGP/17Pb8xfPfkC+OMFAKhD5/3vYB
F5g5SPohejI8PuM+iD5wWhapnba05xf62ZZIMxKETM5P/ay09qjcU5djGC493X1j9RyFGPy8KZv1
02pqktLlwOwgQrT7a6HsYfnivGV89SDfc1Nyy6JM9ekv5Ik4KVr+alr/7WlNd7W2aYOQEYRlpMfA
M4DR4kTyTUwsraozjSrK2ICh0N1n55ZZYxC/VAAO/1USzvqtp2Ty+Q5fHlGS3MtGkD/VuGxYglXf
2wfFIGqS+1zpYadobr67PZT56J5fvSYtuVsHMjcQuQSzS4lDImHd83H3KiUYBATCR5IU4iOlo6CZ
YNZRT2+tNBB24rteDKav7NlW1ipF/ybnZ6PVjh52lBdzqep7Nw5N4YDt/cAkzbMuhAptP5V6KjQd
YokqciTa9L53QfOWdOyZG0EBaLpkAFeI+EQOnEXy7QjMqBkLJMq47/Z0uhPQbd9SwOW6FtnywNNj
DnPWta2+EDYglJoSWmceR1uNM/kkXYKTpFPr+dQ+IontBTsd8ty45rwQR38CaBAGTGrwrmyBREgk
u30OVFcs0rVPPizNeqU7PKPdD1mCyag44Jdjb7v1JS7j98kwg6VHjSW6EZlWSYApQlDwqFPCEPgk
QiqA0edgTrU9mtLkBVAxGPuRmsC1bKDFtqkvD/TNgbctWCRog9wxQ6gKqw+4TYp6N6BBPzRW35ko
aY4DDIm/gtMftK/KG1CnmxXq92Bj0nUyoSZFsdweVGHdkTW7itN+ga1hJnRgn8TzebxCzdjIJ3G/
HZB2eGB5NqUkP5oZ7gnTRkdM3/coaZZ0e/zqfnSWcL3O65FcuP6YQybDP8Lq4UxBJxDtaVHEMFUi
ikcgWdqwVrdNRQyhVapzB6Chydts1rstsMBQHp47MOa2p+rfW+vfCbpuEVwEIlUnb5Y4H5mg/l8t
xPerO5rLA/UJPoinykS6KmmhCuUq0uAWckrvuuiowodHdry1z3V5qrIu9ngkOXtblHj7szIUli1o
NrfN0JJxS8yb/ha5d1Prv7FDYKTuvReAZ2aE+zWAo3ljdjCq+HOGSzgy/GmE7oLtK3ab1YMRRPFC
mKEQAZnz7JUzzAjYmMex/DhsB+1+aNEYLZgSXQZeC4JvVK0SneSkiyix9KRWrRRLvtT9P+uOq+Es
pyf/n3+jjpmahcctYqT7YpxUE+djp2K25vqfEnC3TsbUfIYNOHtcty3j3uxTEVdR23nOlt0xqK3w
3zGqpn3Ruy9tiUyvyUH62/OGg0Bieym4pfYfB/kJOILGIrZW4+abbLIFO1JOb5pPnO+OVeqLQUdQ
aL9yRzDkDcRqn6t+7v1YNl3IQXfsBVLPAc1g6rRSVKR4Us254BOSvykMl3EL/IcV8EZ+rpvmkq0+
YMXRreEHhNdU6DEDAiYM1dBJVjMR5om4d4o6Gx6ezjVrRSigPDBWGNmI1rd5njkE5WxXpfz43Mz/
aaOu90J79vARslpXqYW855dkNy+l0J+jx2YyPaEAire9LyEOGf6aIPonEM3GdloK/iQMoh7jr5W4
mp/zyd+Zi04oaqVTbmjzN5BqwPAlpu1wS4Yis7fEIxf+jamXloP1oHr9UTZ1LmlrbIqSwIRvBJPp
+PI4aJRpuu9nsH1vfy/FOUvBTG7OaPEkHozY6H8c4zGr25q+cJHZ70pJOE/Lz8CvTsmzIJXlPXcj
fVeRoNiztKpb8Spx0TjK00u3Gi9RwM6pJMhE7A8w3nrA6nctvTUmzaiJp0Y1xysgWawMX4LvGKRL
4Ud/wDMNocJvIvIVVBzTmJGCOAkIylBImCHvRyaJmWm/WDlrsToX00fnhU2wSNGatZjcBHmPnT7U
QR6+THhBeEgOI028HVbuTK6SeD+iHll7VKxMwsDUiAEEdImt9hm7Z8gNQS9SspT6n2+IltK3EujN
jPU1AcnGJUH0s4n4llEJqCfPAJW6w3+GzGiBj6xyCB8pPOHvX5ybXhnnSdXQHpyToNnZxTU84cVO
jcD2maXB6LCVMbfr2AahatGcffoDg9MJ8LTOmxNvLTDBuDG+76GqLjmdMrbmijtdSVN7amYssbIe
6boGuNHaipQw51YrZA/Dw8FR0gAqrSeN63Ha3FQh5tGPAmNNUmkQVswbTl4oNnf433unko8vm4fl
ME7coFo2IqCYG3iG/wxWehyFcRpyOb7vioFZjf/t3B47tJzsc1SD8so59MySO7YAhZscBIUd2xYj
AwHYdp7mWQGtFHAFJffcE5UzFXbmiiExsbmLeHm0k8/wp+VNWdMuI1CkYYMQ7mgnxVQD9qhVy/q/
dmp8WCRZNqgh+hRAzr0ELnnH8xaH54rTim9SXRvBcTSixMLLE5qbBCJ2jJyUCKjuuONC4rWnuUn3
kLFuJ1QNTDfJI4EOjmfU3EkE1pKNFN1AbFk2VKQ5Ucic5626BikxKV8xtogKYh6erZBtD3cS7kAu
MOj0+5mZIaMK6eKmbtvqxmTDPfhIFTfAaFh9j0pD0eryqs+gMvjGpdnnPQH0g4HE88+12vzVKosm
dXlYH1+pXGYFAlheyiMhnvFrqWZXqKsEj9dx3+VhgLiluhaoP9sWqjsL5ssV2FsTtPRAMppw+NUt
NWsXhVt7Owo7h6W05sDfx6TWE2fiazBPd8KDrZ8tQYPjw/JpVapz19H8yMJpLhJ5O2jgO+RnW5cu
MHE45+2LDcpa5jQPVzMV7WmhNPp2m4YAIIBRscDd+R88cwFtKhQgTb3S35HpBEz8jEaHBdo4oPE0
xDXXEeLFd/SyQCudmOvWvbiQA2T0WOX67ptRiFHHgGOpx+mw7/dmARshN04DL6325VRLymVFWqzd
WceQKiXzFQrYcURY257T0mVlW7kF9UFJQ2/BsTOijmpjBY+KZ7K8d9ykc+K/kppPUQ4OplZI0NzC
fvB0vua09cMKH3fogItQODdigwzGCT9aOGDKUeXKOn1AITH42yqVa2hf18FxmghC2/+XjqTykyAz
+Sb+UKAa9Gzpr049//Y5hqPtH0urbI5qQdl5eWkIuFKAUQaIgJBCWRBihsTJJuhxXthkdS6IKwOu
zxuU7Shd2JonYy9QKGTgw/cbGETAMzCo1MyV3fLd0/e4Y8FysvBhshmJ1c6zhi3njgck8aFl39ES
llVW7Xs936OOec8pbo7HCug74yq8958/VejYVhmnyKNsc2e08XtZuS3hQxp9iq3e+rfPNx3x/9d5
OZbwY8Wf2e2r+c0g4C+rUJ8/gtqm2KB6m8qCoVMH4rveF5MDNMfwNc6E8M13GThd71nwmn4FqaNH
6eNMKUz0f9/wnQOi8LpJ0zzxnWTaqNPkmUq4Zbjcbn7m4h2UtUCnduECxFJRulDy2uPBd5e7RIMd
sPzx9fgoO6cON2Xrtxq27nZyzV+ttq33ueQuotrDoiw1KwFnwUGEavz907875vTh1yckoT0qPh5c
JUkzNKHPvyuRwq5C5DwCF0LvRTo8oqJL/v2rY8awFoz85mZotiKkXhVj7o1NeNwzem2IYS5knXIu
u4lCJRlXX8ABL7zs9pdsv1MBD1yLluEwA4zB+a90LbOsY+K+Ot5KXKv1GGOfkvDIwFN/B1B4Fwaf
6/+K17VWix5mG0mdHCFu/J1mQtQ8vss0HBaek60aH1u39WFXlu9vWE7oUlJjI54rfxQiazIwKt/5
SLM35jSdPzwYxOG9cyMLkFl5QEmeOKDr4SRLBxPQR5hsdUYWiYugCYEZfKsaIy4LmzSeRKx2Blx+
YSOIBFclNF+tMa94Dw3PIjkEukQt5hnB9hup3ZWSs2FO5Auo8XGGNDMa8ImFfRxmULmwOrfeywBT
5irrzCTdq0Ct95dwexR3+8PRXgNugCfnpVG1D2REkc7Fwz9MvevYA9/IQgrrl3ut7jEcT7jRevsg
qOTFlhFojlL2DM1URdfmFI+wUW2Fu7vGtoHBCq8X/57neJTY2epIzpBm9Qv302Uy71WfiQfJJI46
DF98x3xN7K0Ez+bBb08/G24KgyH1yi2t5eC3VUXEJnuR+bv3ZnoelJMXFrJMvksgEsqRYZuZlen9
Q/aITrftu5guYIBXFNNkaI/kTDvNn/Lnx7AMmtIlNG25Ufc6vbwykQlk/bkC+2RFJ//k1ZRGXfWV
4T9oEwPUNjLkJYlsqx69Oasw8GLbcjthv6igpWewH9d24Wv9QW21ojKI9u+rxtFlrOWjg+IJSiTw
rSCAb99gT3MKvvolAObHPWxrn7DHutTxpL+C1QFlm0BeCfrf7xrhYeWRutnHmEVua/54+z31ERYw
xt/GTtNmEZbkL4yxSYMML3Fn4i/KZ4KHp3hkRRPDQc443DMub/WREqpsGeOthTtA+5HYEwKYtYPn
p9NGkpDaNPWWuwnPHvmxTUK5OlOmYS7qwJpje/LJ5GV/MfgiRJ5zCzEP6CEIqgPbEKdS2sGxuLr8
ScM4s1oKpBBL07hQ0N/ZopjYHioQyph8x+HRlrtJ5332zr6sJ6TjBgRuJqT6cMxip0TMlt6RNrCU
4NIgWiIfiJzeNGf49aYNfEbOW7NyJPf/yW7kUj+d0ebL8EHh+yEEObgDUZDeGxHmbnM3+hBflNrT
ZSJy9IPQ6ruykIa7fHpxcJ8FeuGuanW+5QuPTSmmc7OPhACbfVXYdk4KLn6chFLs3gRy2wpSdNX4
uZPp79vZplsqkIBiwODbV/eo3V2O8jeisgxi5fZjIfGWiKtOhe4E3Hc0NK79UTk6MZMBqDjK5K7s
kI2U6SJ5qG8ONxQBnk5P3NsXmOCqMlffygMtnY3Jr6GMOsghuUJR2jDewTMaMtfWbBuD1CHHcZJw
ZpEEh2tbZ3KTOPXWSm+4BPlqc0hyYYWP1GBWXaV5eZow6hixovY3PntJTgMbskixFSqll39HMq/o
oEn9WYQ7DKNBtv0LuvfWsTSUWVFwv2ggNgHMFK6JxU7bwwh44sQE6XRzwgOYD7/luNg1BxJ7/Ulh
EJxc4z1nnFe/5V3iIkP4NTmm948Vx4IsYMWT8tvZp+2gTNUiZzGDzC7PmlZ9ohnsw4PuUYHS+5lo
zFTw/U1mbokLJUp6aFix4vtvq/ULK23/YuejrX7GJEEosnK+ADNtU+VzwsSSvbBuCpnZylzAvq7P
yCphB/pLM6U/sXxsPrP+fthCZrYredHrY6SPt5zBTG5CY62sap1zojqvHek+BDkEHbsLu5ySq7vf
PKFvJ14ZAGZktdIW4+sPkABU7veI0x6iLJM1XWZBzZAQovzd046nCOcx7JbMSUrZ4N3PaNmE3guT
H4V0liPXm5t3UN6KO/Uy2MkDm51S0fI7g5ixfxU2i5W4cDPCEhtbk/yV2YXiyUYVvBRfAbZWEhq+
EVOP9W6t/fsi3/7yDBp1TN0Ggmfc67Zm7KGmwKyJeHNN5OVnz5rVMv3NjY62KYwmJRit/HXuwjjv
HRwHpqpL6vRLzFX+3IO0+yNIP+W5P0UfIIaXFZYr03lSiOrf6MNoFWh1C5JKac4zZNAPAHQrDlkY
fo2pjmVAJMMi7QZArXT+UGpZ0OkOTcxLix/Hhd1QR3eJDcM7llLmL3KtS0y0WjGabCnOfOWeQCLh
93EB5/UyXBGrvYf/9yDpiVC7m4FGtKxw6EnWK0UpADdSJs6dTqTm47WWgIK0izOIgRa1XwJrbk7Y
9gsTAGynYLaOO7A2uaoRX14e5O0DreMArGB8QFe8umJBLUpLOrJTXe224Fz2Z4DRtFk21A0zako/
5CY/KwVEEkTQ0EW1rYsRyZoTFtuDLeL7CUpyNLNmJsWIJbSaJYYQiWmP2tJpd6qShq5sdS5PhAPd
uquTfl55RbPusPxCjbQq3NRsBjXSvp9UqdMTz76JQiRDKHEb4aFNJY1WoWCoRjS2JCMs/Sjo20Xz
BDo6gvWKQOpX/ZsfNKJVaowd9bflri7zdo2KJqDh113Dd5AlQAoUlooXK3RFMp1dboptcIRtJNsG
gOP+a5l7ZPhMbekHo8PyoJEGumOPsz8Cl+kLpF52f+3O4ARCskZ7TmgxIWGf2FmirnFr01V/vZz9
jIMh0II3v7pP3rEbwRQg+z4XcRxrQ58KG920Uxsl9+HEbb1M5S6P5QDIIsI+b9bSvwXjkBKqlJaT
f26uzUstxQuB0FexKNEy8z8WC4EQFQ6B/B3oj6qXGJf90A3PZ8PXp2hGecMYN4t9/yf6oXKg1C2a
kUadnHnRO0b2ns+t5+XxBtW4vmCcwC35bLcQxPkGV55tHRqcoIRwm/ejH0o5BrmdiQnIlqI0MI7b
eDG4eHYh8iDZLLP63HS4okdjYw89meyt+Cqxu7y5p0b2cEwE0ad2vuy91d9iXBinoxixa4/lZdDa
TsYjv+y/W5rmARL4TF0h3NbI2ovNZBBleXKgrlaW9fl9sFpifJ7fiYgSg6ETkzYyUhhI/q0WdQ++
hYmmDsMlYPjK2Cfvc9LDI3iUlND+FMH1NTCbwLikcxorx/ebkhDw3HbP5RaC4gAcoXYCKU22Apzn
UDzc71kIPTwViB0mzrai23OCPbvaDN0zLzXGUOYC61r4X2G6U8zoCm57Qc29O1FDisNVQIO2CuXt
p0HPIgbrTeCnhcoFCQ2ENgqpws+S3Lh35P1Nlbogd1Is6etPCJ9QAqEDzCWcFFvEFiPMu+l6u9iK
bXG97FefmvzWJXDl4fW3rg36p/wcPVTjO5drQO2XpfWU068WPfwMeePWCO6UlKyQ+StE28SQyoso
ZmPDDCXerZh1rqE9uwTFhJrsQqU0VqBQbqsEI4SFCXFpwcEAK3QG0U5hCEfWBiBepix544hWzkWh
2WiIjVwbrk+BGAH99xNT5W9VHFAK1P2OHIYgfq8rG83wEtGoO36edhv4cO1yhl8NJ6zaEQsPYMY+
ZvBvWKjXq2PyUusTPcSTJdblt/2MV8taAHRCEdxAZROZI7Rt2meuQ21u51iutT+robOvWpIy90AZ
zipSyGeZ5l5DcoZrkH1wz4ZhC1WJMZs0BTkXchoYgm0uGrpsRKhuVi1/1gjLrY92TjZmjtsPLvEo
8LLWLN6fjefSS6pdhpJui72UpCftMNH9szk3qwdWfqrkmzdpotqZ8qh3To5B2HkExh2ll6igpvch
S1nH9yDjRcOaJMbXtS6xuMW+8iH/O7U8ua5npGiBSc52Y+NWTXlvAHV6BSOCc0sdYGw0ECY1tHut
SWdZkvmamqLmWvGa9mitoAIoWednYr8iBDIpEhoHay8owVNToCY1+pjacYiQk/12ifpowtwaACam
YxeXqz9S5uYKUQF8ZHcIKttutmLNjalQEBlzIc0eNr1xbAaoh2rlr3KxCPDUkuY3Og+W4ksmfVJ4
6BfIYgjDelEeOWGzZYbArIe+gOXLqtfUVBzHLN81o+aMu9RS/me8r+lo3NLCbKgRTwvSciBWtaat
POnZec187QdvoGb5dlZPGFiLo7hVMGjCUH8LCjQ4C9iN3ODvgOUTx7CtBoB7xmH0+PQSY3fJvnaC
bhPQvfzKpksc7GUp0sAoVyzAvuUaejBLlihq97TA9gwDafXdj+I+fGQ0HiJRIdMB7KQuWYzav9T9
iDBV/Yt5LMRQNrN6zUxmHXA2wJVDd/tvFBiMzBuD4y7jdWURdD9hITP/WKsEy6PZSPpF78d3pf7/
qnOBHP0cv+OywSMLK1ZApV4ov16nBmQ1DirbZ0trdyKos5Le5TccRnQt5Tznq47ZjoAZxKTY8d0w
qCmUqamteS0F9TblhqmTnyqzLoFNqS7ZH+70qiG0feX22YUmgdE2av7oHOKuOOlBp02aBIA9+dxK
Mtg4pKiV0Abq55+J6SniafEskdvuxqkJsxINNuRk0CA0BMbCJPF0T1W0EsR+n4KL/DthSMc/Otlu
i/lEx3D5PBmUbeuxefvPga1rfKOBYfw84ON5MX32xZOgiDvo8saFy+PqnWjk41HH4k4Wrf3g12c5
BfiYgnxbCF+SXORH2iTDSvAa3oViEV4sDFoksRhoHuVbxKBRo1zZLPyetFVkYgPfvTNim6rqqJ5q
yxxXJmF69tY8E1pJreasxd2ZD9+lFyd8jL2ej18VP7pjMhnRgRiT56ZPrlaQljWdL2TTI4Dz2Pb4
cFh9Qir+Bpu8MZ8r0PdqnpBfDPI8tHg0LKda/efP62zEh73TkAo1gEdcENherqDkvvULr6RtAngS
YBsCzKqq7Cy7wDEV2uhS7fVyOh17ZtRUD2ZTnHd0ZY0mhh6LTyV58spmvkLYO2tsCQQjV1Cwu1OF
WPGrrRx8e0ZaqF2HkfI2lhGHyMbsARzodBur+xnnLkd/5b8I/brxJn8OUW4kNIVuXNGSe0kNLuTB
JvXwVYri/rEMMnK5AY1jmOiXd0NDBXgfohpyOBw55vZ5yqcN3k3QecpWmWg1+xNi3c1SHQHBYImS
W+ZBRYY4vuI5w9ObwBhPChUMGQ2wBAbatURZIa0LAIXcK0dW9SBAGJ6PKh8KfxLcevDGJHV6P2KO
xZtJRVeAwGp+B0LtIOh2eamaBGToeatgcPDscisI3epADLHU+deXH/q7g35y52apaLWl7kgvEZaK
WO0/R1yJCTC7DQu7ToqZ12dEene6+FLjy1F8LawiUHoOll9SifeRtQmYjYCg9900JqxnfBcnfJMa
pPPoGnolXo3Vru1Fn7uf2AvCWl7Alk705rGSfMvQkbuS/KiTRzAFDg2GqUJKviOtV4zV8cfbTM4Q
PdFZ4Pwguf9D/MuOBLMYrE7gUcO990iMpXIK7MetAmNGf6+7wx2iyQ/nI6+EhqpTymm+qQ+08/NJ
N30a/opNtjl2DvwhKZR+r5K2MzlN7yzxZovduKp/0UMAFVHzlmYFjOPv7FG3Qbiz4lHr6166rE9Q
ahyIE4uQYUdMxRPtjQT+2Ye2aZxrdgpujKhCzA3jk8bO1ojM3dsZgpV2hNe1fPyFJi2Jg9N7iB3y
7JG5g2RTRVwNBFgXH0gCy+vLfdNI8NIS90sa3XS/yaiT/kM8boNV+6gMdJx6TOi/70vVb3fivFzr
FDgcKv3yJr/wCM04S6TbC7qeO3f+Jjfis/bm2jD5CUmbP921QSnpM8E7L1+2oMUmnsIL+/XcxKtj
julzXvjQVD2DDoO7wvVdR2o1zU1GiYrALtAZ27H0j1ZiQVtqeTsHJl85L17QZ9Op6sq2AjsQzG/5
tV8jrn1eHxMgW3mdM+sDWEl5cOeNhya9Oh8BhFRugbzvSX/jdqd0Os6Jllx7oEWzlEmlr5s3Ic9d
YyrSnVpeGSSNMcnoh8i+L1FPIMX9sJaOrXd1fwEiKVHt5gr6F5F4Z+phRsdruKkcETJ2Q8jTCsIE
g2TomUFRwuE3AIApPNxxYLb0F76Mx5quly5ZsJbFdmRJbmfhprXVcf//Y24IhJlfUp4SBr1w9SRK
D77faCIxMCquCSPArNlPUlSoMAKjG5fDYY9o2Cwb8T94c7bh9Jp36noSzX3nStsLHQGtMXfgVQ0s
R/TWt0Tgk5+0Qs99mVx6umKoOevHEnRIsJjWsa3c+pbM88tpNPcH+Zamlb/q1c7jktrLg9BIoizC
kzDDlm8DtPrzz7w3TkeWV1I7I9IKeo39HuL+RQQnHwD7VaqbHqTiwc9e8BoxOpjmBm0Ymv90ITbi
+ntjoLdkMXzd5CDQ3r6QvYN+EFBJDsdtrlI0mYvUR/GAwUJiQms9K4re+5i22N/JEGEgZqbADYiM
HIshdoEpKXN6IVsUKAfttRcubNtEQbYCIYm1Glz9geXr70wOYNcfXPklVfvjFrmNXxw08zLAzK04
Z507NciyohQhRwd6tgBc1rWiO7JIYOG+8QqgTUnkXk2QMFML6+aX+eTjHMisZd6HaGxsJZDnIqO2
HFTPRW5xMzCYcvC9Ft1c3wlvB6dYNqbAV36LOtY4LknaH3RqhuzG1HllqEAMrrin8+NHPGDZhjL8
uiZGsHP1ioo4KYhiYukI51gGtvDhEt7d19gMr/o0TCgjbtmaOaqo6T7jHoSF8YBt/wp4+Zd9YYI0
g7q2miCI4NfvgyQYgvGoxaAa0yJ7d/dbCE6aZdqLbUHsSdsdxtFZaV4P4n+A9p1WTAKHn97lTKIr
TOdAaYcOK8cUeb0YRUMECoiNUaEimGtw1ZIoh4l6je6lwbhDAU7UinZ3ZFCjQUH0TpWGNV/bmEYj
TLpq4SUL+ZDuLnVE3U3x/hKgFYQxgPrqarcPKp5HrGrTyFzaKFni2hrUh8Uivje5rcRjxH02/uJg
Nbtjd6X1NaMwRgsQ+Wko7d4wRPjy6QKiGwyMR140R/3587D+bqosPAuR0bd9fh7FW//B/NtwMXW1
2/5xV3qXOPSP+xygbJRuZ4CMx0v9IKht+OOzsSawnaGGnqpdrcN2Nhp3CYu63QsB4EuVvZcTpf0O
zbdnRlVhrMx37Rn0Ap0lavHHxXnUrLkVeBq8I/tU3To+A5vECIkzphAVGHRlJfpJNH0ov7z9ArE+
tpDN8FYzh1COHOjcdNRvLtDZ5Q5DbqdXIuUh9gNIj2zoNI9fRNTN8HM0ja9pdCiSuqcr5E8Vcr9N
w2RATVeXOIGC4aujp/CQ0mJT9pGBtHdrrM8yVhn8H++BLbioCVgkySPDfu+429+zPmQwJPcQyAmT
phHdxrbOm4oVCQ7hlpIqePvIMYJzYzL7v7dbgw9qawXQQA9cEnIU96SkZiclaV5zL4rbecnSgvEh
MAaFbUHR/vRScEtXxwdb3UQa5XCxYSf7wWTzUW9N6f4BVGQCtsZQzZkcJu3UVCcnIggJlGSskSRc
NOElhApROJk+37keq0rgUsFWyMA7S2TwKI7ZkLR0pRuh2GsyMlfYVlPlWBKqZeipPAGvIq9RPQLc
efDwDM/rUy3ZtYMMRbKlCjJdl2vi1Lc54SYh4a0d2kBoeDHKlzBOtZ+2YE3p0juF2shNrrnnE7nf
Xz7bUgIDBGb3T7RHVEU/tH2byW28Ihw0Im1Tqm4onXLWg+RwMuUAlmKXai9NxJtL5HiogpzRuh63
ERsroDKofSzsX7dKRmY7EnE0LF5299h9RX/RRqnuS7pm9amPW41MUznqyHLphXHC/cLejD/N+ADM
XoxIUmpNRh/+RjxdTQIH1YlXw7JqlCjk7aLH1+/CmfuZYVWIixsylZ4JfTgKWf4U7ggOzCODvLVh
HUn2HsD5yflNFc4sjH3E8nBjXtEFw510ltXG83HWT4XVLq+Q5e0QACNfFYaxUZJiBRAgUXENndNT
qViLMYGypY6DH1/Qi50sWvAn9CFEyDOpzIiIKKoxItHc2LyxrxFwOM5NE0XPwqQ9B8ojG6ZCA+ZH
pUXcr62iKB+dSngqPti67tWnKqH6sp7XF5QxHdS5kOjDglke8k9ItzVKNAgoQD+AnIf2pZBuTNK9
gJfZrl609wTw2ZDDx6dnCIN5cbdm6lNuyYhrwEy2OEIJ6QAiLS3ONmRsJZv50ogNdvM5ZXElSAVg
+ecWcNy7MRYvwAvsxYEEVsuGDwbVVj3l02BVdkhoxGc539AKW3tdbUTpZQ54oHjYHG3n5WrkHSp7
ynMssYaiCkz/uHCkelE2PhFM30RhihKaFsuGqVTMpCZqG4OUKYBvOWLU2HsnEL13DiAg//Z8xpgn
Lloo4MKoYqyopyqFozRdMrGfUUYQ3kCD2NQSxYTlNkeaRIWXpNYwlAk9wZNOR75JCkoLo4FgKKdq
dBQa030GL+Bd4/2gV3ONPUPWxZRQc/Fr3kC4FO3Ml7hG/uUEFczY0gZ6/6zu0uM5n+QL/F9x33Rw
It0ZpUFxoX+kBb7l/cVVhh7rnPcywVLoZlvLImT2AB3B2yJiMUY122SPkrH2SNGbwzUkprCwvmg4
o/uKLpt1qekFpmH1uyBwI26cjVhGZZFMyS8YP3YRQFuKceUyRqS+xq/zS/cfGdqoFa3r88vIe7kg
KG8IxogZhv0PYzDxtsFOH2OdzEDb/ijfFTrpELaEUe3eDEFu62FCK0JIpwHbgu0rzNoba6U0JnLb
nRUNLCmx0l2da39wvQy1LjSUj1T1a6omtdfWal2QgoJLtnmsZwy0N9/tJAiXUzwXISQwN40ALjIG
TbaFXnjD6C8/xBkUoHo6rLcxFbbGfnRM0NDEDQmVdoQ4XpuS6SHRDQCxtqECKDIYo5TSDhlrmWTa
PeA9m/rqs+lPtbXr2oPJHGLE2zWgBtS5tHzWyGOSYCcfZMyttAvQowerIwcmnQ5sYdZFl1fHTgkz
aWvRTEXLlBKUcSlcMVbWn1hdO917IrNwj7wcxN/M+IGmfNfEXBnHiw7DA6CRyFGuLvauZ+zFKUAQ
PB1vi7tHJvRlFGpHJv/svSLzyiLRhJpBJ+UL3Kv1bUNbaljZE6kYRv08cfWR/rT5EVKMDtLkHdRU
F1oxJJ2qn/V6Z+z/TNhVrXr9Xvrxxp7DsdrnowSibnMJtiUFpM4KXqAMN+A2BoNS51ee5vWBYwW3
asKhok0ixAae3bE9DCVcl7TgUGQf4psgBwn+9xTO6kEYH7rq8MA14yMte7cOP1reG7LnjzXSwf0A
9blJ2oVeOr6ILVrKn/4ohWWKjkbLfOnm3CLLaT2uST91haz5FoogDDuUdKvT2XULCiWpMaJAAU+h
C9HH48MaiAN24Rcs2XAFCmUSvLlRT+cV4YC+ygeeTsQG6/XzU96p8jNbwqB1+7HuxLxfx8fH/CRF
Gzne2LonQ41Hty29hQ6paZtCrAGPRzTQ8nqPTjFeeTaZvUL9/gHwG5pGL1D/qKk1n3kA/bMPs5UT
y1/2IZ0+IKn5fSj+YbnHDedyICnmrT1RVd/XxWqyYi6hlnbzZMzOAny1aGD4+k6gxhOZLrQ77JAD
VnGeYqsMcELIkiNhybuPZXWmvVkfavpo9Wadi5W8XJMlT/nq+z0fz5AySjD7l071mszMVjH7f51E
l1iJ9ZygznSgMzLnPQFyI7hDZdosmCeQCljv9EXPjBQVeGEch+A3zkyPBlnEjvI3LWcrwEZ3Nn4d
NRSXxF+a1i4k9ygSUltup13Avfa340mZJN7yHJ5PQYyzRxx2Cb1JNj0PXGZauerixGeEcyYiYXsH
0sx1Ydkf61uO97idaxisahq8ENckv/OFbH2Cku2j5a9aaZdxMQjMe8lCzi662jymj67JMG1gmLan
zULAyEnjrIYXeQ3jvj2P4KeL4vGThpZVmvvFTj5BDuM4ayVqY0hJgE4ruqEGQ3aCwsHPV+4uT+jp
fwQhcjmB0p7FyiPkHw125VJekpc9XgVf+nnElLt9JZpQhCVGW23C/MjeR0xOfkFblmbcefpDIdmb
I31wwbSJGNZIApdnPYzpKb+/JbhwL0+E74aO57UvM1KUu69UczpWqy+N+qTlT3+Bhu+xq5y8Hisj
qtQPKhShnmqLeTCV3CePBSIpKXo2SEyYD37NJZP2W6w9l8m4HxAdyPGHfxpDvfnjakCVrG8g3AtC
OZUshGptxHPq0YpYb75cjiRI9C0COJ63LnIAvNOznsjkn2tir7dcEiTeeCyaFJehTc8TAYoQ2Gx6
f3WCmttYzpVK5OUxiK8INfrl+AAjzeBYA8JHMxLDpnoFuPbEWr1aMBXgG5n/uHXFRkRBzfDjl/ys
/OIc4ErkbJybOAmE6CbYrNzXgEgvCLi7rozcEongvly0uJAZaHDfYsIc3moDzqMaLIiBOGPCO/UK
UPnFeJh373J+goJzl7vKqmr4IKc88C1Mk940ou+gqz1OvjZkfChWA1lD2e+bFVh1wrLfiv6oFoey
ygy/WPHQ+5TjrDM431Z89cPXmHTM5fVGuaSyqI1isIYTYYELqnJvlnninBpzdCXGlQbiJnD/NMd+
J6Su1y2FnczV5AHfYi5HAEC9o4Fabns4vZZ6zwCSho+vExuEz/7nIGnCkvPUnOd+c99ygQyaEh2C
AmRqEEEnTXYU/DIHrhkGtCtxhRyA+50C8/HIkVW8diBQiYgEBSHasBki+FsfAz8WZul64t0RIkUe
nOcju+CcgoBOROoBB01N+KTUrnDUHwbwzCkWt+cRvDjgThlprEsEH3VbjiKHykkZABiAn++EvaaC
6gLpyG0ILmpnJwNt1iQxSoN0rT8Iz72Rvj0doEd1JfqcI3F+0fF0Lr/6IWtw5g/Gqf1j+oMqzA/V
0IqtJSvHhNmdOnnDh6EGdhbEPyKgFtEZ6AwgySKQ7HvC7SrqcwsOf+qDplAcWsYHfYX+vQQVF9RA
NKzcjW8ql0rpcSzlwiPjlyR/TlN8UtAuLJfkLilNEJeM47EWJJAu80+Tb21ZASzMNlGeGnHsX8H5
DrwNiRuUD/BQJoVdatbXU/IYlOoswb14m7Ga4rBXkXFV8YFWxevlHbgqhjRcQYSJyh9Hl18tLOGr
Q4pNLqjONS3wrC8+tdvXAMPRb/Wobfw9F+GYoXST8y2dpeAJHERJg04bGsjH0G4RzSj7+ntqBDw+
7lAk/N1osHEwnUYvBa0nivD0ZjGll02ZKeVPB+we78nWjR90BabdZHb0lUsO5hRA5q63jcmP/J2g
MqExNIUGsUnirxgBixlVCwxk8gu0vY6YDuP/c7S1YhOgq5tmkYOobBOh99a0nwMmPk2UkEeA/vni
nhmE61tZa4gF2pU99qQEUYT6n/arb8cvhPgVBBlrrTb2YKHlgRtPC77UjantiU6rnKFPWajxHlXz
w2vjb9dVCTX7oWGuDMFIXCdVIf9HYFVxF55BE3kIRzrNTWULFKomLAKyrpXW1hH1eILRV2nnldTu
fcVDz7Zn6I6hBb/gIReaGfactZDVxQby8AhMQSB21znNkkpqqXRRtICVtCzDibb8DAKigtU97zeH
Cb9/XBHkU5u2HDq/sX2gNWi3t0xPS9Ro9XB7qd99SgYU6NO9RAmm0ieszyWLHsUGRZQevN96iOoC
vwh+4/jQNuAFoniu9omoUN3eGIfJG0X+CmXhEkickJBS5uJUwrSfuYkWMwbAkSMLD/B1bfmMYCtd
l0XtvkP/xX893IDT/UKvXoAeJTfPTe/gxrcEdQP5uPLXTwe3EiCXK2cbmuF5LPnQ4f/bd2M0YLov
wPlR1bg3TVpKSq5lHJw+m41+vfelUxEzPZgONhvuNzzEnvenT0pq9GnFcTS5GkwvsXGX8WbzPAEO
JrdRJeQeU8iJrPH614nN6EKnU/3DNFb1pPn/GjgzWv2u6vh13v9BfwiTyAhqCjmYImnOsaDjmyNW
oWW/HlrYw1IE5mwvDobQmSeOqwzqfCntd21mKy5ZOAKTNvMyGSbf6o5otiXxBdpgE1gSixvJjPYt
CY4vrEGM4pMtPrdzExE1r/UbKK/BiGvrMoo5te9okfaKMzNaC5BL2Br5l2f14G5QTMeJAKMED1/8
IVkhwZXgI4aiYM5ZD4kyTwJ6hfW6bvg3B2elGjeusjR13JlCh3hBH7jEpozip1ItTyFJ1P0e+4vL
Xa2bmRCVV8zqQ4+tEM2LCHH9BWnWYWTIqIwd3lhvlrMCnUDS56lL4zWVnzMbICHGq9XtB7dNsgHq
2DW0xifY79vxF05ZFi9lzFsMdYhAW8HQXVRSvb49HJ5C3pQqrOQYV2JSTc5nWLTHRBCWRrZRYiB3
ty31A930CsUnfuDonrGkrLSzJmBAsvx/vAxNt8jh8WfG+iGh1eEjnRoLMDAGtmXoyx+KoGc+eo17
5kjSGvPzlgDeS/p3+skoRQ9F9j5kmf9l/z4/acquZ9YWqZbBwd8LOdASt3JIDoLyayCNFxHCGWYv
H2qN7uaMHHXjfqALweWQUSMtFQyTf2I7mjwJSeD7/+P/r4sLrV2AD8Hi48wJbFXnFTFiZqal149b
5/LWD/5Uf0XpeUXGkeDGJ6nKR9T5z/VT5aL2PLrbs8LLzyyeh+/MSxHgTPGtP6QpUN+OCS1pvtk2
Q2t2wmUqOr6b+H3MJ4CK25vEpD7fiUp3izPbYlJ6P2LKGVXumbORZdhfF6L8eKaKgDYXW6idmgaV
zPMwmQOkHj0EEXxOuuGjVDAlpmzsFyrwJYXkSnA3zc9yw0nKZ5Z70i8r+M5Kl04Jqrh5QmuFu3aq
IzUl0Txq2+i8YimBmM5hiHGmfTaP/xdp9RijnIGFb2l9LvGKwguCOX+WJoD9DI4H2gXHl4kObyWt
ZNvC39kCOji2oJQ4IwV2bkXMw07peQWYaH5aLmFaXLhP4zDXMdwhjsxWFeBY+um554pWpZvwyBvY
FJcCV3Teru5tZBjcs8LQbNyNpp5cBT/HGRL6T+dvyRFHGvytD6yBmeg3VJLPV9NYYxWX1ulDf2Lr
i8NjmyP55jHo4CI1RKFkdOKx5u2sGTc0K1M4txnVmOFw8N1OWGy+fSfgcDYBOc0alJr3diCu+HNq
WNAyOSHPXvtAbwjKNc0XTFEjGQzJL57J2daZ0TSz+GL73ZJWUxlWvF++TP2XXnpU1lpoHf7XSxcZ
9OpXjhPrBa0PFQbXPVxxpdH45XxwKPg2xaW1kI49hutWDUinTYCFtmZ3T3W/ISgGK3x1YjZCVtS4
6wPaMMQcccbks1GYhCpCL1FbTs+2G8Umh/PVCklIZuVxwjqH7AKWdoRCShPrs65qYVGT/SGwKinJ
CNyedM4r1YZ/ZeghAzizO3qrpBHA53w2xzDhrOf/JQ+w2lCMkvIf5KUowMNKt4uvhdLY9/w7EbCq
9Kio1ulQekkpH0/61cFgosf5WeJiBtAByI5C2CgwLG/YaRUaoejg7ijNJDorvYkONXcJ4bvXkq1h
9YqBAJp4B85LPEU63dqreqgJC0rMrqfCl6GOTfTEW97jrntKwIE4hzXJ5HQ0aNeTVWvJ3J5YZoF5
pmM7afLLrvzYsCn1DIAarqUmDiXsHWznP12XAhewXiBf3ZC9AqhGUBD+6PNFFj56EfkjJEuBDKPA
Ke4DQjxVtIgrtMqfVhLZhhqkHUrebchZ+fQWlahNrgXQUr1AreStXdDvskGOSVy/4mDybjjkxvJ4
aPx7Weqno98+BYi5DL76kZassPsX5PZqeuEgHTbxDeeS6SW5QoE2gabSbvQRgErcvmjgc/jVQQ9y
VqXAhVpsVEudw/U+E5PbMBWU5nv2ycF+dpG0ASD8GlJtwrC4osfY9LAIv9zHfK2CGou9C/B/NzNJ
GfMxQlH+uBSfD0CFgcPBHze53oJztEkKPvhj87nmitORoz4iFYx2w/KMOoIEKjZe2CTXUInTvebV
9MlNINDARFvFalBjqmdl4QGHVYGosEM+RPSFBhAcsXRAsgPeM0XNSq8wwq3Rnyu1owz0vmbjZ9aa
em/VmR2fq1bEkPWe5Is89xw1E7KHHPBCDCpnC8BnaECTYmW09KlQqDLZ8pEITHBmeJ1GuVGSXYW6
9L77F24WWGeoL7qzzxs3UN+hLZAOvnyRFsZuejPHo3a4yMI/OFeToMGYAAbUWuhyN25zN6pWHrGm
jH44sdEZZT6lpwKdZS0Wkhrsg1OQH8ZiC2Nwq+PByYVCR4CnCE1OGHMsZBwwpexaMjRwU+WZS2b+
O8m7GU+WJi1R8KRHg/98+XDluoPu0VCHGjx6DyxRZHe42Q3px2qmAlxZ3UgSot7uOWL8t71CcNjp
9o1Xp082Y+rT48/r/SkYWVzSyfgvkeq6cjGwNXpL1mTjT/dD/pUxhxm1HRAEwkSzZnyUxZTLerRp
1cod9Gop2qVj5yQnvXwrlCP/lXAiD0ZV7UWUVbtjoDbFc8pf99hV+ucZ0miiGpX4wBpj1A0g9Ads
RagwRK/DLy9k8UoD9FyrlK2bh811mxuqQms7pHAFI1nhgoMoMsVpni4Hsp40ePAGzqa66Eo3th5n
ZLusDbIJc2uFOj2OsIT2hEt8SeNKDgrqyRzJe9ZKQzgovMgO09kZO5zfCDUMjTI13VWscvQBFx73
84t+9LGqVuYKi4tcE06eRGQzyakkioH/zjRFcpBccx560gC4X4b08bjJllB+ByoWoabsOH6A6GEg
fulm7dzMYjWHRm14D89Z3YSqH10aLiUrJ+ZRcUibNh1mJp758gqSFs7FIkvO24BPT70c6V9QrGCK
uvIU4WugNR1f7LuWTdavKL5meRW17lM9NQuYVA7a3m68qu3BiNUfhZRajjbKxfnkPcp9qRG/sKBz
5oxPbJwmTXRIbAJH0gtqje+v5izh4QRnEQ2SONMJlU4+yrNZYEV3BIiy1jPa+OYQA+E5ijFXA2sb
hU9FFMX2S1LxnFdlb+/A0Q8AWSx32wwggWyBWJXNzhdqW9f265BRptCz50KBOpXgHwEYddzJ/Chi
kHncZPKk3RuN63mwsVymla81Y7PipIAxdta7WWcjxENNlVgBpA9Hbx1LExzswg82HjIvq8gDbug/
dfSkxyvJHM/NHjPx/ZqWliCspGvjVPY1zdqqEvK6KfAT6DixyBO615B2ZBRodAgqgEpJ1NOsDMSe
lgg6tm3A3CEX2WA9UxKwTV/cheWHuFJ78LlYCnry8rJT3i50DcVXw38SM3lpBwbzut+j8AusaSSO
mbzJpvPsZHbUAxzQqiaVwr3RzwwnF1VuncAHf0pt6Go47RIYPP7k4Zkmf+gs/1gd4DS6+MkmhdpH
v1ve+1wI5iykWYSxIdQYdxtgnTjr57AHSJiprXNF12Z6gLaRazSoZHBeJFarEmu6lUSmnDYbg2T1
SsIaL8lB7bImICqujKECmCAvA32b2Eqyw9QAvLRxiwQ8HhSznKQRVwrZV94a8kuN0TEHoYNeST/T
q9yG8Xdaj5veVf3tM+aQoxPYi6OSPgtvQh3m9dUSBwiiAnXKLAa0+lqYZJXEuD11dqACRCtKJU0d
7viQeOOF3omo2BoYBzcgPjsrdHj0VCY2W6YnFV+CTo7s9yAabNQVSFQdFuuQUXztMAp3GPv3D+xs
7wQOuYNgJ4DKgGd1uFK3kIB2hTp7fvibg5yI2diGiZOR8MKm8PiLdN9Qjz2xKF9xv06rD+oWmkp1
6xKk3F162GcJtDwdrYn9dYf1pINOCvw4JfpvHYoCX3+UlJRq9cEQt6HqNdXiMA25SHU6WaYD+AVl
Tz8ud5FK1+4y5j2FfAVrd6GEQ6q7TLwigLKjiaOyRYit7uGpyUxLQIdMBxIYXdhaeAljTFyt3CK5
6aIywQLwJAv0rFbKYWyRrJTFuTYgalVNr99FHjyuJmo7e3V4z0oXQqVSumbfhq25+CUwS3WnbX4R
rzadqZeJaBxPaDVEN4UdIYJBBApI3u8ki+RMltouNVMpsmlQ7/EiNsAnwisbg0euXVuaXwEGSzV9
Z4V6C4xWU1BZ7vbic5HcnwExn5P0jVmd+5jfWgO500ghNRbhX4GXd7r+cRroF9O8VWJUm32BJ8Pw
uJqJTbd+KrVTfCClroS+BaeiAZ6XDGduvbnv96H0ndS42Bol4SAmiF92+dT98dTsceLVEEeziyVm
z4487eVvT2s8fR84BXmndFFcftOitA7J7qfRofyr4hwL7vbQShR9gm9YuZKnqluAWTeqsi3LYQwS
wn6jPfyZ5l26dYzEs+cJAnRFOzJovFuS2OUUj6MPzFy7SA1fmm6IQB5JLtwWfh1QAd+3S3T5ziF9
ITmmESRD/FmPGwcSadlymgzBCY4Wmhg4jHExiY8LfPktLvwWPpkUHeLjrfcS1IQCW5X/+HtkE3MB
TL1jzu6I02LmhRQGS2Oy/OO4uh+hTZM4Z6vbsTZIMIMn1XfyDgSkYcovZHhRY+zg4GX37+KaCiQK
ncQMTDNPsXA98KQUC8+Cawc8L9+XL0y6RmNjUxV9gVQybf6yGlXCEtxvTbOslemb/Q0t9piBhpNU
BOIiN4c5ynxK5xnFCBwHs43q6xB3l5rhQl1rfQONuI/8mDhr2xOwgoMEojW5ofE/m8Bg6O8WLULb
/N1xOrMIvXOGOIm48uyE/5qHf9EfuvLEbZi3374YLdVn4+fYXeY8k9XZyY/+6JbBgSmIc5hRGgBY
fPFmiOFEfCsTMs6r00x9361hgtriIYpayZbP0ZeGjV2W5GyGtpT4juMURfqaxGK1ra6f8RwRcQF8
6vcBM6nx8uU5hz1go58gh7DGDBMLinnzOC+VDkKZB/ydua8t9IwIknXlyCI2ReR90dEOYNeEjoN/
EFUeJDT2HA55UTv10BetWcF+6KNfeCuZqt/iimo2cNcjKI5HDogYlKmHduUOy4EX2ua+uIaH1tL7
T5kLvOxBJMzFF2lXrT+l1NAM6lSHK0tC9MCyMqfKurMfPOjoNW76GgxxE99RkEZxgbE/9hfTZYLA
whUB0g9akaPvZxU9/LwLURDap2MXfhHLMFDnAFcRec/P7y09sAusZPPgl1auVtKlGwNXIACQsDAo
idRWUSj+fmR9upKXvkxyc4hsLjdCsKoy0foOLa242iTgsph86yO1i2/8AndIMHlej62Cp06RvTyP
VWOZrSaKve+KGatE7HKoodLw2CH2OCRI6tGnNl2b3Teq59goW7fdHhbS5ZMqzzG00k9gf+e2Qo7F
D+Mn1YZLgrneOIYNLqrM4Sm5p3RqRBylnfFIRjO2mZ0bY820ZAT1eyMyzSJFaSO5nK50c0kt9o/5
1P+jTrTyuE+jwmfQBXARgoRqRPT3DNBBnqSR3oxsyQQtMkqfGdy7ATVoHE+ILX1B+wP7IRasTpzy
4/4kGAk/GaZ3l1vlR+38HvX0AsnoB2Je5S8Moe9SxE+RavW/YMFEqzl2nrePx4f0fjtflWMJtu6T
yIObiufKDOM4vgMMz5cmmapANa577nTKncaWqvbdlmNBoj4PvVJysdPXtBkscSH6UQn3Kv8awxeg
lI/zo6iGOYEgjOtu/KRlDDZSrfA3Zbg0NG57QA1glyPo49L8YqJKIq3QY83L9m9JI8HRuXtiqWcR
R121Up4aI472/r3eU6jFDPcLUubgnn8ZvpUpgQllBdhEvQ7e702KwmXWOruKEKXgBWXu6yGjDaWq
CPm9fVVMUORviUthSci5E65AsmYVrrH/n9amw2i5MpBPyROF/hl9yMe7Owt1ZGe9cQ4Ehtv5q6RH
Re8DlhOf2U8J01jBdhM8SbPz1jXOwWH6k7wW+WD3fPfTx3S/Bztn4mbtKqOZj0/EjEJea1lz2Ddu
JbxMEbOCpczC3Kh9CHXvWhMiWpeRdGhPfIlC/b/RrwZVwGmEIeFJWiTkVC/GgHrUbtg2lhVroV3F
RzeOWtdA4eTXh40k2aVlRVzkHDjL/dxwAvZ2haUvRosufBe+1ydW/WI59INLoxTjxOFe6IfUrHIr
7U9vauNOe/AEHUg3ePyWqs0yvpTjDquyBfAGm8wbfEuYtQQJSE6ovahHH7KA7vgb3b1x2D8wW9+I
qg9nMZDvqau8/LyMhW0pVZunQcGE2aQLCXP8BbZTHrU8k40lkKKhnKrsHJ+ipGK76mCaReMCrEVK
GezKGJxSwivM1vZITBmHRRxJ6xkK6qhw2snKBWY/U8+aFoOfwOKIZHNewwRQRLaqChenhBRbjkfS
fPIjrcsTSnJxYxdY/6yvMI4h+Rugtfl2LbognNab7meZBErzpFSOQL9/LLTfdJ0x3dzQUmj7dOnG
3bEr62v0BN9PXt5MDTI0tEcmQQCT3SUfSmCNEYFgXT1nwzNA6gPPA7GphvGm973xP8aTZTqcJmMB
OGl87A8fDmTwdESAGaWwHsu300Drpz/Lkc+8QH7JlQTHfPv3dI551+jC4bg6XOcBRVuPEal9BBn1
snIQFrKeM2aoBJLDEoEYLNjw0g87OwQo6OImnQhWrYzc7xxBJ7vHYp+6qM+/UH0sTcbYOosw2YY3
B679GfDeks8w2Sm259SRzKw0Jq1uEsyvgjyTAqVWo6fQny5FCLmyFJCy8lZ99eOkQe58Q7dp13Er
FhT7uhBqwRDQjq+6wGIqxvCbR/2END1Nsdo7EXND5y7/pKpeyBxKNaK12R1xyPEwMOph7OBMv7iJ
I10NeKdzCi86zGgJEn/94Fh+hxy/SSxtEjLpGQx1gjeZCY16sUv38TFO71Dwdh4L9UnUaOSpkvwm
oDERZn6B4crzTJ0e6HxoCZ0lkPrtvbHxlhNtieU8/TtBjKTv/9kT64Pb38wxH1yXahAwtzOC+j0v
2er9K6H0bGPFMccMP2DUqIbUejWnZEIoh2pRykOJt4ttCfZYSWrCYRiiXCdYtnSIJhVQNwH5aOOh
L1nlGuHsEfFfnFpBV/djjuw7eR8sXoaStkLfJy6r9Q180ENgg5GstMWpFbh4eI436VNt8YBfsm8V
r5AITgmaptcpEPN16w4nrGoFd/lGl8nwqdx2qeLAr7/xEiI26MPO775sJ/stsSWgeVBZibdpXY2y
K3aJ1FWbz09lb/bWSYsO5h3Hle8kPXz5nbYk87UQhZ8GOpDCcXEzwXK2pJqLJNY/WjfUj23KzzM8
IyIe7PkZINJKGysQwbo2FxBZGSh17CcLDGpSZx0DrhmckvCYUz9t2bvtgg+Lp/KrUYRkzVX+sqfm
olaXjxQncj4+S7ZHQPPN0Y2R8Ske3ED1gc4M1UZVw4kY9e3rPUi5vHVdRtA3bb5ydJFLj4KiYMpJ
kWZvRt71qc/0xaCwnsZ389yW01oWcmRQL46gcLE5fmBu5Xv4gBTv9+7nxNvVNQI3nUfsr1YzXj7H
i16rX+SgLd0K4OhEMMLzfLKvyArQ7Sz7BmFYCWzkPfYAyaQsQTD4aE4BWphyX3OwLmpQSSMV9ffJ
Im4odZ9iW1SQDBITu/U4WyQBoir6OT0NhLWBLPWgfGJmLChNc04ZkuUHxt1XsQR6asQQYI97Q6o6
hLCwCKQ4bWuLllRy5KcA/aRwjfQmikBtEi9jSriGAfyyGAQvHzeeG7ljSp1qr9e5joorea86icuL
7EWLsGyMyMDfNCLxmQoKzSqCoqq8lgNxU1e/xC0zb23x64uCG5nEhI062hwamkCm6hWZNFtQIRSv
LfLAMsDJSWXv1KJTfZEw8jsZL+jYdYk/pA/AAaZ3uA0BFHWu8GNF/FHCWSLOaTFHvphRt+ioS750
5vHJoEM+Q5qCKIALnOiQr6sA3ZKYj9sqgj1cosEkwUJ9Oy1yQIm7a8/MgovZx3/tRu2xYZ6Z9Kqi
PtgS9nb3Gpcb1ZTJaYT9Nnp9Ceo7rwUdTwSYrnMBC2/ROTMyxwnnQjvhxZ1VfXdemiHZyWeb9xTf
f3Psmkm6JduV0zayCgG4+Iv5glU/PiHNmauQvyd6A44lr4Pst3dDyvDzxxkVa3qtQcvj6PwdRphg
0zAGB3cv5s3kZCZy/8AmePfz4qDDVIyk4A0Bd3Ysnv1uUIxADBRnlsJnrBvecBwZ9dMko/1ToPnM
o78oN0jgTEPI9ag6aII1DvJnCDTy88reppifelMXcWWmSsCLRGFb31Xtl6PIU/6+j5aWfBODoxx4
3lnDbCZ2kGxoHfRBX4OKHYiL/EunDZFlE1jwROgO8Gwa0J+PuELcNrPpPRlsCQ9vFCBJghwrdsUh
5tHXgaXovBthJ5mSnFtDINh3xbi+pkDh64RcivYzXmKwCfcGPmYeicaIgykbFcaX4oDzZwKxpl1h
hLlXyvyXzmmN/GZXkxhhfODUKrd4wgqxyoAfT/GUnlkfCfXC2nLlI6GIQTumBB50dpOluDybNAN3
Ie/H59UfD1Z9CLdHuNXGhIKAeVEtGbaTRnBjPxO44MIUfCf6s7jwjwEO8zAIBYW3tCchqZOzsV7E
WwNXchzNFyQXQ2tiR2JZpfLl6caV4gBLzpeG6pkFv4yw2RY3WsPlcBdwuZUAYyx/UgF9erTz++up
uGhxQw5oV2fJpajP0hIeVDD+G2dTbc357PD3HUnkYIUYKps/zrF81r6rpGa1DKGvTDfSmx6yyv1J
ou+aJWjAzRVkXn9rb5Ux7TwqIYqP2DuZzHyTvwW4FEPvNsTCOAUcJKbISbicDNuKMyFnOQbJITiJ
McRyj0MO1F/AfKO+djQ4NCzxRf3rwWNAmDdBr+wChWuZraKK+nbg8OD5B9hrZn5bSdiZMZRLiYdp
8kXsEAQ94UNZ0Lm8660eW+b6EpTtqJp3XjL7x2qLKFSjaoPREKXfX7PXA+p5zkyjgm5OKpGkk9lQ
KaepPdL/b8fsI76trdPpBjFrLtR5sdO+0Xr55/ZSa5iXuF37SRP5YiAzz1kJRuAcgLFW1mJ7UEIU
IcmzamUgZv5neTdVMXEBxFJxnQWugHtJJCqi/ZXyRaSDotbbxTfB5Yo28NhyhUgedsWGjTsNAHoT
z54CSq7YvLqsEbUELm9y/eAgtnhtDkarENWy2jsmGxiatpzTwrstwmN5B+RTq1JbkEQko+obpPFW
iW7ilaROX3MMYu3pUJ7irlrJ37m1O2yPOk/aZo60V3BpXz6wt2FxxWL3Wtt+ltHW9GoAxdubE2uO
QJN424u2VvLOk34xc6fmffbBD98UG24G6D2yaYtPJxgimeIAOnkz/CVI0ajHmVeJZeEd926NzoeS
m3xw1JZfi20svZyc8yVar+dFD8f9EzTP/YhV7IdICMcNRG/I3nY9bkK7QGW0aBec6kRO3uzrn8Cn
gDiorusff4Bm7VOuFGt9WDS/PBTA1EzQv42Pk6y+veOn/jqOQkXUX3IvogZJiShkbCvzPrR+CVjf
izIe8/z4Z50lyTiBf9hNK2UhtdfC/z1wkINzr1Z4FLfHrBCQJv3FMj7RIlLtph+yyMvDk/X2ePKW
d1AWwGQ49jyu+B4cN/+aDN8sC94H5Ak+mNi21i0bc5mtNLYkHDMk7AILu8WwqtqThsvX3Jo29l7X
6B5r3lSdtQ+2OAsd4A9pdGUI7zUwXwKAU8UvSpa8/GQJsu4hpyAvYn67NzvRwmgvGVm5P87/fXLt
tHleq3HYmxVNDGPKDveiYGziaNB4+2YcPxlvcsB/Ih5WqRgHNjj0zRxxGoJGzRMYVYP7eTQL1Y8R
k5/IKw8wQL8jgdb8BQIui4cUFN57ISGuUQo8F1ZocEN408tJhKjQRDE0PDzneJl/AhJHgH09J6oR
HJFuhrFvCKIWiKA5rvwph+W2wgkar0P9jQVgXRtz6zcy7t+Odaa7HH6j9Dk0VGuHlGFYI90OW8CE
GvhRwkTOUavEBmM7k50BUfHOK3ctQ3ezMyC72dE4k6CXJUhQP1Fe0Hdo7gu2fLA7BlMsJjceMzZy
VrAVtOoiTL9ycYYdxZ8X/bwmiv5kOd6XCd+TiLYQuLLPAFLSAPTNtOqNGsnNJzP4D4Ep7+Aqf4vc
1z9RB6KkJ57KiZStWH8ml1NdSOEwDDEriUfT+Y9FMWSYnQUgB2uLjQpuNNSkUwFheQYZsimyipXJ
cpxjtdfrhhLi3vt5iMtWGEubcb9jD4lZFtZtJfnC9HJs4YF+GtuGRq6AhFG2PvC9sfK/1m/Cp9dD
RkRmlDq8k1QpCDaSEkFEBzJBmUfW+/87JuQzJFGlFRS2DxiA6pC9hQjPfKcchyAGQQkVDLtuWQtx
Y8XM6nwvZWkuA+bhbqCE2V+OVqZIfVoPyS4qjiUIrj7GDCclNHuD+nK8QaL30MCIVwAErcJVU1CV
DOeKxLjr0AcufxZg7eAu+23L1MQiNyBcpWjkxSQm0+PVXq5Ss9N7GjelSaBkiMLDEkcD9RE1weD4
dLSWif9UMkaaaix0qZZmU7cfa0W64koihBs+oXv0WPKrD93W0Jm1hc/kFIW2loThJpmS5KvOSDjB
OzH1MKUD+EWX6I8Ut1U95zud73usXLr9pA65lxGmdPlSeBoUi+IVUajC5DzwgQPFg+aUr1AXD0/u
AASnW05uTabTspPcggUBXHImJtZnhSw8wur9GqVv4GfOOh8jN5D1wKXWhhZQ+m0AHqcIWKTGaPl4
TXRCjb/nJbf0Nv2lLAATHlwNl2vxIM3sc4E+n7LSXPxtlEhUfndMZD4hv00OT6rk7LR+m6dXxFvl
NWlOMNDjHTlfJyGTTJHwvrWGyH2U30ihz101v5jF7FCxMrXnSVrjnD2oAwBmSgKfzsYFWtKbDYDi
DOLCJvAQrHu21/rZGnBhW8Kt1eGO4Jo7hgKGU0M34YKTRLWoNil8aLhi0q2+DHkAxDorQw30QaSz
BqL1beZrXYTKBdL8kl3uuG7yniM3vXznyop4F+I7CCmSFOpM4AJPGgZ9M0+o+4pstmryJy+gf7+4
U/nIJQ+1ycsv0wE3H0Mmlx2x/yE/GkgxGiF9rNkAvfim9gOMsqHRWYygxCKMUXnjYupWTthK7KwY
BHxJDx3tLyWrTmYxEsEOFfqzog3wb25SSr8nXfysqBHICuUnMgAb8xfRHrivGYudI15ikwboDN/W
evUlcUTE0ICb+1uRTqUPkiMYYRbLgORrTDLJvtTjcmU870K7msuPLywBxQNTSXBj0OWJyS8Gbsa9
/KqpqnixvOeXtMNu2hSur8DFSWH7imwpsIIQAkRrLEvDF2eWkblBJJawCft+dSO7J7J7mrspNcOM
qSyu8g3ORtieLeL/ckaWAk1+X9zbprw6zLIOpVUt4/ecAgINt29V3jetQ58o5pGplkHBUcD2RWv3
cE382FThta66gyuoGSp5x0fhhnO26ZeXS2JYU0yUKuoBZVNrvV3M2+Iz0ZxeVw1xLKcU9ivQsYY6
4DClUsRzQMkTI9M1F6w1hK6ck5VFgnYNtM6kkmw6mMobS3s60+867OnNFjNYuY7pyWx+01OYjhop
kodpJ/vAwZgiQjOT2NxOGoHhMi7unEgfZzPOPrf3HuqOEgDLeQ5WW2+tcZLK9Akvh3EQ8KeZI2UI
dmstB5xNDGeyukqnwzfUsfc+yKvpQb2TT+1e+AW80DVt5aACB3qXAQjHgAjx1ylnpXzBbTBld+5u
d6sJkWmjzBaa5wZLtov5Wa02mptrsRGbD50aWzQdkjm5iVPqE2a9ZCpnve2vESblQnM+snhqGdeb
/rUy5sFX7U57593zQLt9C0mr2sCuCAEBlvN87MyoNG06/oj7Av04J4OhBuw0m0lJBmr7ZlZKHo4R
JOLUKhAuAjdmf1rwAngAUeXCrVSkdC278ab4j222Nz0gr4u6PmRRUhx9pmooZtBUaSEwY8+76Mvk
q3JBUrTg50J0RDrGfK6OKhFRfObWfeQD4bs/sW1M3C5rUP+Tyg+CEQNUvp9PklKf8cFn5HXFSTi+
+ippZQ3CV0x6VFc3Y/oWB0LtLNdmedTjT01ZQE/MWuQslj3Jvd12TfTXJzKoZEdZrhbAhMZYN+cR
/cKsVzZTA/lhKMUtBb/KOHGcFbm1yoYiODI4QYuYUB7uvJinxJjlPArC9Up4R7r3HbwBdQYOYrhM
n8CDpETaVIKchVuwZMedvnLznRGzG8sZB7pxdeAKn3CRofkZr2f109cGlN1wrFbELwPkn1TJ/LAN
fQ/rItsgSwyjx+qyWPtSQgq2cfjSZ1yGJrm/xl2uYVeu5LFHgn8Q8fR0WJ1SJWIvz4uxsBXvhtEz
Sf0GOn8bu6jfk53xu7Rf06LqTAwA5RjBl4w2hmiP3KuG6+h9ZpLRILCQN3C52XXeiHySJiCy4K+W
Syi7cqMWmF1SkeOw11wSTAcpfpMHWcsZ1vr7HHvr8tyKrKrXF1VU+EtkE5WeIa2m+0mrh5URyN+d
oJ8BrOJcFydeAVUa4DNLLgT4EzIXZGyMpSP8ydNGhF1Lff9Wh8e5Tn8MpCx2kzwlcbxY8fHoNVbb
8EaXVNfpBl4T1/XeEyDbdrCwSpNor8Wv+3f1dFhmXF5gMt0EwIiDhaibSpGCcEMGUaDfckc3QFmy
qg/NjAyDc0H5j+Zrg2lFEDiBQHnAVhbIlh69Jhew0JzP/en4TUpim6+quEPD6A4L55BwmuvbpodW
3s1DFu/ht63k6Fqu+mT7bmDzPEDygEDtv3Gn1utR8EPn6L6mX69Vc88WFlsnJkzeZtshO59b2hRY
Sv0DHbdTiU3Uz24Pjla20sOKp1ZL0BaxfX/QjcW91Xa0eJHB3SZ0k9mNhMQ9VUWC2/mAkGF9/mQ7
74s0yWFsTRnplGAosYULCcfa81iHmdzHLUqX0TYiYYaFxlouNoisZGToZGxDHQjZNNi7XHRuycTV
+Dyj81W9ROsm1onesG9OFnnpw/L3RxwkfTPCvEBsYoxdTJ+HDW50c8/KMinemzVt97PZ4n1Sr+rt
1FqiFC9vYsfc/+ExYq4VfM6d5PUdACALdaYWNBcCEajZ/l88i13Ns4MBU3FCtc7fsx8TdxY6Wv3U
+oxP3iwTzMHn/z854LRIIZx59rymrMa8qHb0MY5XhMP4VjaCuMNUJBFebIIhCZmEw7K3idlHVg3i
Nq4amwxL4Y2HyDtLnGefdutLIJ6+Upc5JiEjTzRruuLojr/w8tav1W6VoQPTcWpRaqkK119X14a5
ODs71fHLUX8G8TJbXBb81ZW+L7Zxi5WDPd42VCprVDQPsns+UfDjDlDVPRYQAmmuAGxCudrap0ML
t5Suix/rFyxqo8SPGcHP6N+ImsLqdW4Hw/8/C/fp1PPyJx01NQzieL/4VpOpCsw29TvudoBa/FAl
z6ZpBwS6lyJa48Wt43p9vQ+thzhhYjMpUPVhs6qtJjvCUvh80FRuO89PgYO1EXgnfie5uxh2Yzt+
zJcxdL2ADcXJP981U1q8pvNdrA4J+dI67JtzgJagtdfYqtkjhQh9dVix1+KocxzNbf8CuKugC/f2
p5sQxc7cdUfzObSv7OeHlIPYeXH/rQQ7IpuV6DaujOJPclfSsI2NcU/tK7FHJVaX5THBwYvu4e2y
UllkMFEKYHx7yHWJF7ScgLGMyFER6cB5mHlYutoG6dNNSvKqZqBQnRdOetm+kwK9p1y5ulJ/VhfL
58JymRVcOuBYXqtCEWEb9ONyme41xmVLXaVqXLmmhV30Q374j1vBaB8nB97U6/T49paRorGOIZnk
cgmjVgUM+t4mOjAJkieRp9svhFPYRDuJyqRYnDT0zNV+LfKZDClp94lK/3sSlN5H5sMtvjWA1OUN
Zmq7oVTJgQ8prCx13t31GuAUWuOV6tjddxHei49JBAi1JrKUi1LF/cMhBEv9e52VHG8JeaITABm9
iG3THp+afd10DjIgzOB68dbLU9zfydO4YY38phlcz4Xw3ttAJcBru2Qguivp2r5Ns4pYavdnArVG
ZS4E60HhaYUbhCBgvxqaK0YX8LJgBY5FyLs/RyUksRm2tY42Cfgs7YO+nOtA3YGEBIEjXKq+mQC+
5WQEYBrDKHQxTg4B/b1bsEAk408GFFo0hCYUBNERS5E0wf4OWdcfd4xYWH2yWSm3xp3tjzJdBRiB
bs/YEXJSocTK3++xtkkY5mjcwbPu+S77NUUdNugiulB+R4DXPPWJCKqhn1bFiW1pdxIXozPvz4eD
jrfbY1h/DDAS61L9VkOPT+RDCZB2f/E215FuI9fpLBjJAklXHnFXiXgAQvCn0ziVNuO8Wpk5hIyR
JPTJYXGMJ2WUlzQMwIJPZXIxciaXzRaahp6PrUz6fERedha+TBv1SWva2n8SadxiWxl8MmVkxy+5
YNRp7mdBQsC8pei2LvzSblT40NWozsaXhdUsAv3ogwt8q13x5ESE2HyXcnuJpunYCmp463IyXdZ3
4CV3u5n+0LiQCB4kuwXlSBG1Pimgdis1tgkx8Itn17NA+AP2jo0lDX0J9RD5sro/aodGcQkwK44h
w9KNRzBOmeEKQQbjtz0tT4xGrqoiXI/pMZeYg5ffn4JDdEh85K9nN8v8ue2tNnXJ3LKgvXzcuR1a
niqe1lBWmRn2XjxYDS/QJmhHpwglSq534RKf5tFcB4myGN/Peuo93QuH0jCG1M/JnhYt82kzX38W
G2arqxwEm7PU1fBHpHc71DFfKDCDk21/8+tdEx+ZS9FcnYuMsflYqZB2wJu0Q6Z5xPULwA7uG55q
Z+s5fxqbptQdIZOkJ51m409GjWekj3XE3eWV9YZ4rdBGY+RZFmDkvPE0TvXqyInzE1Fxfu45QYG7
dHX7dgTwkiIGeIJ/QMkb0EOflCYtuOtK1277uiPcQoeyfUHQEiLnEq2kYiC8TJNpiO3kleaMWTOR
5XReBIRUwHEOpuDlyRDrcdu7yUOHZWjrK9NbXT2T1e5P86QOz0P76cDV/XYshVt1yhUR78QQMBRp
IGOZj9Ti2sAPTHai+S2xSEajFl5sYM6MErcx55qYjBJeEig0jte8/tbWgl1+1xwUNh21Fv8nH0yL
1AHrYk20TkufZTyBZxyPZJr5LjSQZnuK5tj8yCMdE3sOnepiuSn5Ivk6bapRA/43QzlEiCN2R8Dk
jPlxpxnXr0HxJodQbyUJXhZKj0tsQvPu1jdUVBv9O0UwvZLbhBoxTL4Sdd3OCD5Lekf6Sn8BTWI4
rioF1MTyfEs68X8BRdbO9msxUPgYl+7AEuUIywaqBoAn4jFixDbrhj8hp5KEG2jQsEwFbIVhXsiR
10flQF1j4XRA+Io+pwr+fP+hzj1lbEiJ6ipoi9AmvKq4QAmmr7fkjTq/9b2q3EtJHsl/g6bNG9Kp
47S1f9G8j09A7bEkzjb9YdE2OgtrzCtNR/Ec3/syYtQhGHhCvGcOLdLoBWLdoStgm0Ij/GVDA9h8
YDEub62qOWuR+FXL7X6oRIZ9FQ9r3jdWyjV7UBcC2iwe7I5NfJuwg++qbKy42I1HXBp5GtvLG1gz
8mnkM6ENfpfnH3CuMJB6pJMiIwZGxkZWXuqur8s9CIpoU8bba9YHZop8uhVWr4pxCluUuPegNkBB
m59Dy0u7YGW98XyPmtQzb7tdD4JThaGJM/nfMaJ/h8IrZVwRswq+pNuk6Wmhmrg5mc9GwiyE3qPG
7qJXV/e23p0Rg31xkV09KnTV69/klZMvknWOeJoZTHTxayJmhxUSQBJFFNrq3eogfTS7WK/0sS7o
LGaA9meCXGwik0ddl9qLrhPDDbGrYNUoMLlv8/rzR0a+CpDUO9flY3z6UoufgWluU0QrfXfNcAsR
tas77Nl73ULrwlP9b1UkwW0eMDq/ofWnBB3ri06dlehFkOd82MtdENJb5/kWfSrtB69Sbt1GF12p
bsyBtBXsRWDrDJ7z76EtnSqMngIdkGXtJNWy+H071GUSC0+N1Z/pO3FmodLs0XLEXGssRwmLfPHr
5tEQfKL4rJXCJDFjI1Bie9WVuQIEtKzQaZp8x3gN5a3fxoqCzXsPjpT/zArwNKm46VOC8ZIBgyWp
Gh0ituEdWSdUtlQvptXFhzepXHQOzx73DVk3zeaTUJZLne7YveCUqY7NXTbNHq240i6iELOsVE7e
impJ/I3d8NGbXJtLvdV3Y6PBnh1TlGRSts9IlT8SGOveWv7eEyXtbwCm//dX1TzhWUEPkbMsbenA
kissB54XabcuebnJEvAtX/BYpXQygMCz0uvWlpPRFJl3WFXXVK3TwI5vxhVByOxPV+iSbCawepD9
Tn2uxFaqDwrcFv04Qbo62d0GWhjPS6Xrmcwtn9Lny+9EIjpu/H1Lh7AQdkSd8v/5ZfuWmR6eJs47
wnZbtOClE0HNCItuzx+npjbiaOsS6Y1r86nI0TV+95fnRzrWIuKx7VZMyHnUb0v6YHLqvRXL0Bmo
t9+XHRbKctoRMTJhR3duVOO4tIfbyh+1lqE33NWqdSMSyJR/SR2UBgW02tsjY5zR60/UBz67WTHf
2j8rHi7H/s6cfE8Vx9IHczrkIJAOKIpTNS+L31ejn2HveOXUTxh4ycKsUfM8G2fLKyglIVJD55DK
HJDQV3JcKcTbo9u/kJaoQKTVHck/45p0HD18Mz+HUIKGDRZwm7RijRsDDpfn8XKHsWnbU2OpgjE5
MgT+kwhTVA/9uTN0P1Et1D2iqbg86dbPNhh04i3qN3P10La/YaYzwwj6li6QiThJFx3FKeLFiRWs
kk7ERu5BX3L5J0wXXWC4JuBWRfmvDf0xMjs7nzQW62Ven+ARKdVFehrhm3QUj93t9X73gVI8GM3V
+a6YGNRNmhSKktd6M3YEx+rGM26t/gwjm8ivn6awU31SP5SkvPHkH8CFSS+qTY7PGnZpPKCNh8Kd
v+kmLWp87XAIY/Oq7+eBGrf+OHgUhsXbZa5bGqQCOzpAcIdY1dzuMz5c7/huoy3Je6qET1sBBqgs
9fwaY7zi13gSiA/SA7JzCODCwOeUS9D2ZgPSQsho4mfqf798jCduEtSoIwIvqlsWJIZ/ox9/bfR3
WQgVXxL1CaoWHlrezTo54PWayAIaP+S1dZca8Wz32MfE/9CapXcD2tlD8MMHZ1Kfyc0w2igIQTnR
IL6yxkOn2kahkK5JlLFiMzXEYcI224KH7tQbULDoBGT3rDu6sNT60qLLKbuCQaFw5ShdjzZwAN77
x//qDgixdcz1k2BfTtggtspudSKELW69FOqUsoUeBZLh2mJncGdHBcDpze441LeNuSXBA24tm6bc
0gFmvSUpLxmLPsKxKSBWn0egrL9ybq4M71Q9az4WCAi3lhcnBHKVv6OyghOrzjr9R1zejblnE2nc
HP/p7DTlHZ/rN6/CyeIxeYKEQ5cF7i65K58k69kOIs9R5/+vBnNQgR5v7losqEZ3frdlZfrK+Dtm
7MXJs0gQc73QL/u3a+BaxqQcSwmbipCi302I7ys6XwIVQ1QCJPtvQgRarUeQZC7buFrOk4YllwAt
J2x5vgNa8GpgfqR7lAYgR6WBux2hX0k7c1IGBhcgutTIsKlFRPpWeVPCxWXxo+cWcu2V6UfFvifz
RHt1zTWc7MbJexaod0v/LsMLnl85bS8+RbEElSY5GYsPvk/i1/mAjAQME97piU+F/tjiEhupqZHP
RHICLQGUF0gX681FEDBIztXeszANHD3CP6nPT3tAfowUFoH1bykEUybrG4zFCX/+NLefa4P4gSPx
qCZAfTbGVyQ7QOomSswT7E9xQQzjszdu7y65erbDvfFToHU7xZxxEQK+dbXIfCpjBJVJMkVkg08J
/dUMvVpfv6Jy4gZ2jd3nagjmjI0stHo8TKm7jRrmdTTgtLNGu31AdAQrI4JfRLO+Sh7JQJHUbEPu
lMGUEw54Ezb40KKg5pYGaOfPs3btvnKKF6njveym+PDnGdb8UyqfHT3IT6rpuE+usQCd9weIbcYw
FFOFuIjNKBACYgoLuG7dLHqAsBTZIWMtTTS3riJxVdUpaplq2/0Y+nC53pFbT8AdvaONn6aRupJ5
pZ/dN/92nQySAU/hXZ5Wx0+OGMwZyjy6jubaOBXZCjc1cSiE9BOK2NlKxZ4EzoH6uY4AxR6C8mhI
eHVTQdCiL8XxhEUdX3pA5q2LXygL6vhxVxWuZsOObjpiGqrTBZQ9jvko9Jx08bpirzRoT4md8/ak
5MW3eBsoa+omavpNKw2QKmNFMegmBkglRyjg9Dbbb51juoNiPGB/0fKLP/EWNbEGimfDiUDof3bt
Fw2vtCpYwzODDeAh14J9Xj3jruOnL3CUSTR9m0O4+0otp6GcLCr8B/LhdyN78Z5hAwnqDummjwjM
lxcOP+vu+As1SNPj/UqZYK+fJpDqT5uvsR9xUkvCQ6lDNjRkQL2wvuJAwFA6IOB9rjmYJrkg1Hay
f/5yT8QRPbk+GFDMv9TvMsZhR39/a2K2Exiy3DkX/3ilAkiSmQlxgINZd2RWNEixH6zy4lPcjaLQ
Lj0goFTDZ17qe+zV7ygerCak/+XfzXnZinOe+rtjie/Xa06nO3Bct2gyJveVUCyx0/AD5GpJ99Kl
FAIYhS0+2o3U3GK8Pg443P6SUA6YlkYzpS+kCumYoKn8p6JUPuYfBjiTlDSkmUh9t3pzRp6cEF5N
pYhrZsiVGk1zve99KYeVWq0FInsqcbeY06sw129S/c5f0FYmZEREqqh1jnJ1txQljGz1LKfeIjOl
egSR9oNvu/O3H14ngQfpWbExFKIukf2T6j08CQ3t97GjibAd7p2B0GlWAs5TaAmxFS1WNI8vyY/Z
+9hOmosWdpGScWtlkbtRhLtk4h3eSNGMXxy53TEkLUCPkJFAXoWTlXn2aEpgqA07oBkaRc49HweC
PfZY9oPja56M2qiJZ6y95RxK9N4rtTOBoqJvrksx4Ci+tJZVtBLjuh31F/9mS5Qu3dIU4oGddp5r
AXjUDQcIhsxRC6O4VEyLCwFTsLvqH0NxMhhHNBmVwhIa7p9pr3Vey8mR1ahN3YfdvYnE2EawLzZ5
GYJjOp9Ts4Tz6uxqeHX+p3VqcsdU5mbFFEmv7P+pEDY8pBz0DSvkuJJGSMPa/cg8JawGcX8y3pNr
FPy4z7xECwoLCTMDNbWQdOavJj3SdMeXUsdagYW4MivdP/dM0aAWyf61iVK3N8bd6ZVxysRtA7Ib
kDI2A0z3Ul4gjVhDWcYYHeW8JHpE0iZgspQVexrPrVWmpV6CB/C8TYAPTIuUQlYejLaw/DclG9JE
JEPQRCFqOeh3kNyHOPx0t+OJ3ljNMHyD/EzoZYVIcbcnresfunG43PPS1Kb8YWRRhDcaXn8sL2TJ
DS6/kBvvuSgeR6syC1S0BdWlhKDAEsCEl7H4FqPAquTdYB5rzRp0T6vniREGY2lNcOKBvQSeBE/z
itl5gcA2LKTN/DYxKTRvKSBHr1sBysPFp2+A+SDWAjMJBU3Wte3hq29Vp5hbXkvGGSB5eHQPdZb5
FGUU7mBL51Y3Mg8V6Us5ZMIccv3eHY5YhHUDUFxa7QkvyavlEpHftvyP4Rik6ibPBrLHPQg2y7Xp
FhiqlOsMbxA1oU9iUVDpaSlEZY0zCnVIBUnGP4nEyATu68d2ouavbV64tLC+c7anrkxrY5w4/k4T
CydJkRmivrY8x2Jmi6IU8c3mA8s2cMDMnfN7ia05AmvVDKqeOUfHxLwR516RhhgBPAoSNLMdMOFT
z8n+tZgXzsutpxWpT6iQ/EP1xQKR6QfUQn9wAT1ud23VxCHAOVZDcaVIBfclftorw/mFNStMy/fH
QQhfzI/FeWqqUfpJneoOo6bthsAbtQiq9Y16vsU8nf2kxtGtvxpCHaBluX+LrzsbLe5XdrVPXOqi
3W43Aa7v3jrnaHTBHSTbd4zRxDaL6KHfj6QS1UTXTyI4WGp+SwVMV3h12WuY+9vE+FM+eolmPs8U
JjPoNLWA5tqjTro/gmR/d+CMdMUra/IaWJ7R76m0oKhMuJ7i0jissemNHhgjVYnumBbLDC8xijYn
7dvv53A98emEIfH8803ZMz0k4Bgodax41N4Jj5m3DVv7QvQkMYkmmw3tMzoe7mbwPbOfYASFnm8J
rEkyTB3fFbd4Vxi0gib0a8TIK0T3q8sClZw20rkfQlYDCEsvvfJnI9cUCeBslmPUoyvIT88RLXaL
TK8Yc8K+KE5eSRTFQ3eQjOJ4Y+b9797B9Cm5gXs6KGhR03LYHKr/TcFM91WpqNYqCjUqzLA0IB1e
xv6vGKQYXk7M40bns3UE1PYj0WI83tl/xoSjbdFblCuyiyqCiLpIPTmJsQ0SITPAzusR+d7UUFqw
4bTt8gcndX2gUULQPDTBnTCHcWV4tm3G3iMJbWeoFuk5ClXP6E/b1VvCGG1FhHKyY+NjyIy63PD8
f2weksjGx1u540382flwABwUCC/Jn+pSt5P5RfKdZDx4025tXtAwDeM4FUGUz1N3oZXwOI4bfJ/N
SyxFqIVgD0JPTTjDVDKV6Zl7tOhbqlI5dAu2h+iunluYwd4BgAQaeEWHlVxy41QJSs+N/Uykr1QP
iEX7x8imOnnsyX+Wgw57SkrBiCyU2DmSvlJ0arMec72hI4ZKcyNKgyyQsceSzhLNUJs25jaJtZJo
6qqpvFLzxsXAPjVlV/J152TV6JeYIzIkKkT2QMmnjOX3843v9sRVXPhm9CMpYm9nrQ7a8IKMfac8
znt//qHRh7F4Uyk+JgHQt/m7cJyHG83Te2xURwtclBzj+dLvARBqDCC5rZ7VOhqTNoU39qjzh3oi
n+JhmvuCP23dwQuHZgbB4Hr6WS7i3eGiwl1FnZyCh8Wh3xyy6dMAizcBxyAKM3/XGhrE2WAPE291
dVMpBtIG+CIEHlzS1IwIyH5v7bPSezb06vYZ9PyvcBsk0cCctxJtYYzevZV6mz9oj6qL8FBMM5mA
4S5NvmQV0B+ani3pUX7heyVByW3A7oR+DXitYGfOtK3hiNumouuqgTse8wTRfgd/48Uf7++htrPw
udd69gcVnLc1S0lIdbrvnEsNEqDXa+6u43S+eJ7U1YYYih7KeNXbVs2oTXE4vLo/2jrjB8twOuPJ
R5BAVZq6hnIZo6I9A18XRDiiZriixXoTZ6sAVQCJT5zYawMv14rK0h0k5zFCyYVtw6YdPP9M2Hq3
WbyIky6IwFEQFQZBxQZov4LCweYU9cBqBlNqJm8QfWRALeoqNdAEBAi3Tp2JeC7/asVIGr9P2pYv
j+NEflXhYmDM0uf04PUEdO9piHbuwhHRIIHJRe2kd1ulhxJzW29C9wocXP0BC2pgShdjs5gMyk7O
flbdReQi5NUFXs7nbnqdz2cH5Qb0IMvjnw5DHLPV7d6Fn9OByM+LS0sX8XOQUChBq7BuOeqSu409
WmcgB7r9FZoHH3xABw8a2f6Hl31hz9DNPkJ2+HmQBxT7ndf1Lg+7aEGb8QCeCxyFeJMHEY5kKj0w
V4Ki23icnecpBhOcC+YcXMj4LeF568D4AsT5kNdslCTm0ISXX/orMvW34ht4H6dm6ToKpKJxAO+P
bPO6e3DsRApc4URxS6CG7Y8ImuocZYHD9Bsg2m+Ee0rB/gn6Dob+8zO/MP+XBd76BHosPazV1NKn
qh+CSdgTJCFFNf9itzJvTSxKjKf7ysDJiaAdNF0LxLx0Dj1sSh0+Cysp1po4wp+3UOrOdWEQW6nf
cNjFuMpljkb20vJIjBNuC8lEWKsOziAGdgzOiFovgFl4vD/LRF9Lzn6dv/pWiU5v8PWMsZXmZDfg
OwiikYNwrYkFsMEcQevw1OEekvnXuRpjYjkjTGgR3Wfmk486/xvsc2WYiiYyWTqaTXW/X6QUzpYD
0F4ANiVWN73Byxz6U06+pYMcsAAZ31IjB6dsYLgSqF4yOEWIqpFQHshf21q9auqvsqHHrP5xDUdY
5DcboniefkWhFe/hFawya+I0j7ScSeFEdc4uN38CNYYFjKdOyuKJXTaGpWy2EeI4Wm8sP0NUXSQk
2RBVy62MdTRyM1ApIym+Fv+iOboOVQVfRUszic5E7yfEpaYRtaRecO2I4KlYVanxNmyVsE11v9t4
qGDTkNpGXsoA8+5Ero9RbYXDROlFEQwVowOV0lociVzB4DqF7oTqZkI3Bb9OJ3qyGzX6Qyryn2Mt
vp9WweDZ9vccgtikAEtkD3mMPQ3GeJh+h2LiOoh4z6EKccmIL51bNPvkpCuiuIxYnMpTpoP5Traq
CEq8bB+z44XCGnnQB1hlmSXHUmAP50L/MQw3Qu85UShuyYf9Go36JyXlUOLZlzjw23fG2WuzkcfT
2QfPojpSpCeVPd7TB7z9xGVnjhruOHd9en+L5s2AKIsuiXNNmrNbjTV3DBxipUKS/vCqoqSusZPW
pPSb1heQQf1rA+TZa48t5wTBbeZlmS+QjQGgQCCGlJfWPmj+4sHKR7fqPoFgfym8EinPi/XQQxR8
oiA5oyFlfsSK1jP4MGYD9JP5tvmR8lrS+Kl67Gi3LclvpZNe7QuwKtDMFifUyeei0JK8vgJVsSVS
2i4Vo9pIIMvMUFiaYGjkz3i+pUUfKOYnHzNyGU1ofU7xrpHVzsbfsdDhWaFh6TEY/gLgJoNoaaX2
HAqFTrHIhH4j9f21TqjQ+RLs3EQq3CtLb/ftMIiyQAEg8/yGpd8FAYG8oAY0k95fDOODZVRrkZ6T
zJRuqF1bD0NCgDWFH0pqRyLeMZMPGQyeix1XxLEuPSIp+RTY/A7dVvsbtDmHKPyxZtsJPtxiXFLk
0WZEOXa4NU+2mhP/HSaTvFsoFxN3qWDzE1UaO+j9x8ypXsAXbYSn4rJrv/kDrZUbdHq8DFWXwmU/
ButY9+zqJWfBl7Q7oi3E+tzdgPbwNmfOv67PnXzkXansg4Ani2iR3oGBCIDJrqcylVDc3OIqpN9M
vPQ+n8rFnT8d67W+EA59aKTARgwjXhN+qOBX1KrxwJSfEZnRd2S8EWZKjH0P+9bMXRR2F6xgNQc0
4fyOwdjNI/GJa2x3FVvY2ZjlFScHaaQ2z28z+rj2XJER4SP0DM5xVUslrg7QCpnIZAeWnuEdX1M4
gbcZwgfAZfhtbIP29v8tX9Y9fwxGZFUsaUYFEJEY0Ycl8WNIKJrjUXbcm3oXp6tKCLUtSwNL1TO8
JGQgAbUgk38qSm+fmQ1tOJN33Cfpmi1EmWznRD/NU3oB9/Nv+UCcfMLVM2ABD9zNBKMWkgVUiW41
gIKJqeBezs/4rVj4lAVT0GECFbbzKyZ4ZPlmvZGcpdDyemngt/wh65BVWl6qBlFUVReNl1kfKnGj
U+T3ewmEul+ikDVUkAGqD4t8pEGqGGrdVTPA6qMktLTCKEWFJzQy2oUVtOygKUXoWmifc9RB2+c5
+P+Ss+hdk3vF5EptijdkFegT309fhTrIbjkkUeKgTNAvysVe0EL4IIf7HR0zUF1P+FCJDTuCSJ8d
fLkaYXsBSizXxHO6Dm6kKkDHZWV6o4e3n5dhmtWkf7uZPLfdHWZMXpL6v/q5GWWHiRmITCDZROTA
XB8jc1etYFYiUawZUNPvHNfr3uloZGSeHVG4+IXPGRgClQ0ZZvF7oMO6M+o35f7FYzW4ZxUX0OJD
Ab+B/wkBwV3YChi6Hqr/2/X7Xi5AaB4rsRiJlJfEKRaVRPijd5nC8k/TJNdIIs2s7Wkft8F9gqD/
gIu8nvXk7TEoGwwvQV4EaBqOS+S1gsOKXZxynCKHOhIxlcxEScg8C3J4wQf7/0yw95epjoeYAkr9
fpfaqsQ223fE/kX8d0usJhS+0poKnzJxzBX8qn1g+y/Bdy+S9lNpkVnmFCuUwYWuS2UKhMPupnzl
LX2n75nzyNMA56KN/TUST2kpl4QPe3FKxqDLT04QsANs6k0jx3gr4ONju+GSF5mh0pmMHGJP26r4
BK5eVLqPVq6CSZM3BAEm4qMZCGH+X+FyPLvl4XZU3o+IszYj7ADdJc6qNDw7Tboq4UdBHsCnF1kj
RrOj3BRkc3W/q+wSsxzM2eiL+fWdpkyE12YPlZO4/FYV+0L4Gd65pKpEBkAtI0K2CKbD0XGsGMPw
fKZJyaP3svXsNFA931nyPp9XdNYTDtYQOrMPHZ2gEV6qg37IXxkEALtr4OgW/eqbNLhaH7UjUABQ
OAo7hr9p29/HNrT8bdQ8v7c1JFzbCYms6uXrfimVTySidrcUKS6ZpfB+OBcihI2opjbBQna7qxGH
10LlN35ivajZfD/AMInNtKq8I5+nxQY9cHBWSP8sAIM89EHNMkpUKjk7izQsaF7+rNFYL1wue/lr
XbWUT2S3DycOVsw8KyDqEC2MSc7Wed2pw1WUBf6IQ8+h5AcpNLIuVYrVRW/+ixwUblrkzkqIgrgu
ljbX+7tn4O1qigw3FrJ2N0LlsZe433Smzz1zmAu13m8fceX9fhSxDfdcKVsV15jlHR7rHTs7WQqS
gGuHUtXteBuJQ0tISi6BJnbzVW63rJFVTNyjzPeeL8PS0qUWrzNF4wF74xElO2Ag/X0g/8DrZDZZ
M2jBIQeCAKSpRTZOXtwvqFtnMxLr3XEhSfgzILShwcSMbUP/YU2jEwKnukVfA0SsZgQtgvtYkzFX
Dbw2M4kvvUXnFnVOUei3WZjEovnrq3/NjtIKP6PmICrYHB39++6RVyIuDvuRt+Cab4pAUV5vLhnN
pgBdpAmxfYme7+GkJ7OjzKBHHMWqT9QEqQKcpCi5PngjrMIpBYfWKtFfzHF60uZXESDT8Xr0WNUe
2W9vBnTYt2YO2mTR4iS5KwKxmgIotVxKDQVZZ6laOd23tbPsiBKVcG5VBwfv5uF7r7HoEJgshxkt
hiq/9K0NJR+d4L98dwwspjRfaRHfUVbtsx2HA4d1xq1OKeWK34V6zS0D2zf9ds06CGEwZvRGsq+1
Oh/3cLMoKqhsvAdhPRY28u+iBUYlyiwPxxCPV/qdbCj4Eyd7tzpAfT1LyaBOMgyCI2R7v/AYy6lz
PsInmKlMT8N3Ra/9L5jNAoPGo9waEh1LVkWjH5MBvxq/Yz22zsow2TVUZJX3QX/JGsPl3QrTBx98
qzuzrJ4IG8EEJ0mr3hexcCBvzge2FLDctJMyTQxA+nrvCo9yOF5tW43lAPVVBuJUE91E4aiQ2Y61
CRiuRF7LI+zGdNNm8dbXGEaCFW/CbNSdXuFjgmpQ7pyqH81VEFanHQ8iSnguQq0AZ7fyFTEgzGUN
/CVjWna7PXR8Mg6W0LVcK4rHXlN+rQAGkFtwhCftGFM+rwaYKwVuQrE19YjORVTVKnHVNWI3gBMK
z7K08ak06pHtj4is1GewYewINv3IrHgEusIXSeEdjJMF5wim1HzwRlbNPERXe0s/ZFAJLSK7S/Os
sqINSS4UTBXNRCw7G0rkQlP7OMlcTp/5E/7AWTWMtv/DK51fRC3dR1FBasoOTx9T0fOKvkuOwg/u
t9qElKThBPSXRgajTOZop+cDl6g2rqp6lMlg8G/uEjUxsg1z6t5V9ibuXfXRBE9TKEJQbdoen1dy
9d8XArkyEWH0EASxxjfxDfdRlgwCvwHT5H51TsWtxYD7Ni8u3lMBNRnBNDZHXzq5mwml9AABhuF9
yMVzK8li73VcIC9Fd/Ef2iQXenOKUY1/Z8E6Ac6BeahQT0CfW6GbI0x4aER+pghw086RiT9T8OuH
3ageZoDB5qCsDHzat7rjM0Y1Bx+hEDcKTpniaiUhGGzKbFatbcZyd5XjH/s//jOVz7hukDgcnoCs
n/gPrihWwAj5bRpM8D2zY6Py2ucIWjs5fnk9qWu4DNa8zN7jkpbGRUTOW/WMy7724S67gDUB4wva
rCdJ1mcoRAT1vXBSuou2SKY7ACIDBnASi93jAsYb2I/zVzN+C1LhDAq3yq1cv9jAdUK/4AHKO+xp
CQMWnrvFowRRCvmRfAxMXleAFeJO83PI4oiYhWu7schRD5oIZfuZ7bqY5hf651cg4XUQ1v09z2YT
mwNBrpSNyfaZWRQNqE7UFaUB2wZZsYIdM/YuS5gj7hjaC9d/TiqO3s/Te7X8+rN2Lc1iGUq0CECS
gDb7NBMG2auqJPN8L64SrjQhwpJahc/RpG+UEmlBB1wmKfsrr2ujZsIIjBcbqQJK+y+pONy55ihk
DK4gTjG7ECeKyaB+bzvzmeeK9NsPqu7FrcVkVsHIGe71vB/J+nVM9de15ELVb8q6RuvjukZw6pHs
+jUdDVdmywL+49y8ajamXpKIDgR2Y4JZPDaShJKKt+NS2WGGKF6KVasN4tKjb84fSrtOZ+5Lj8kL
0f1iSpQWligsExB59vs7cDYFOL4HyQfL+evdD4xPQZNNWkjliGpM+vTawpQPSOnqU6yHGZZLrfBM
LdwI52r2Bc9ZMQmfs2m4YMXh4Stmg5EYQCyR0ueKYWqA/Zh+m5fxvv/xgVZJXGb6y+B4B1iHsYxw
AWwAH+XlcSjsMNnUpP+wJKLGVTkIG64Wkt32NO686YfkTxH4pYwS3VFLHfrBR8hMu822bR3xldYL
HLdRXsgJNXPl2ue71DOCx+a1K4+b34Zf8c87/0/5dqgkkVeL5tRVUXuH34u825LFKWPch5eJUI4U
7YOKwNvKrivDjR9N9sTW3+TI3re4pKqXXR+dwHYbdTrtUxwI4VpTDcS2JcNv4WMYxfZIoR7mvZrN
G/PUJL8TsAXwn61haEGZJe/lf1WVeWAa7hrLj6Vp0XXP2DwjE538lX60y03aNcOGj2B1Vt9fWZam
r7Mfr72ZgHeuxPxKuB0HEFyFNLgbp/nU3ZeTg3drm7jZHtUndc3Cqyz9F/OwKcnILeJ36BrfxXLd
MZ3qAH6zFGh9znHxowkAxJRhkj/wT2HPZV66VFa2NwKHCrCYYhq9ebBw9vqSmueb0GG8qIT0iihN
2M1BrURW2OcoOc5MjrZenGsI4iYEzVRigX4sQCvD0Gc2ArQrt8jzLO/nkBSWt33gtpKlfdNWXJSl
os7/PhiD49tOxmtVphknIzkdpKyBkM5sxCMlp3etHWlzjAatwxDLOC6Za9OC5eKMCU2WhB5e59jA
jho1mlVSqoI38oJBtPuIh1hQszQEfzpHZSXpuoMgszlYG8ne5nhI2z1dvvbGdg/tQyZZjZhgOov7
EcYNtga8dzIGWjV/w+QlT+Gae+kNeVgNzrvUJwrxLKVLK06FGpwV29RieM/xY3DTlHbZ/2A1f8pX
jiz2QLwDc45VE9KQP6s+6S4pflXX/oEshuUEjUpIeDONmVeUx7wsZJ9/Wj9k1IjlA/63Bhv6CslE
wlQM5YiOQYXAUeKBUj8TkWBeGBEXPbfYktbnvl8P+no1lCsKoPO3Q3b9n8DFP8WMRjKT4qvRNi13
Tg3eWE19VGCp5ThEaof1dTOFQ8LWUBcigJ/lJ86dm6oxEpjk8lVtmiSg6jIh6/Xt1K4J09AXqv8U
L5zTmBUBXUqntnm9WK6TxgJspJMhrQM0/pVkrFlCsxQdqElFZfikGDswQ24PVo41adiFGlSjGgV/
LoJNwOKEYqqvtimj1AUNDMlIMFP/cJ3Z3bbtvPMBCqNmj5T6qdN0ck7gAUqjAc6O6TOad9AHMmX/
rCjZuKSK+BOpvqYXNUFBWs4CeqpGNt7/WCSHcfD69zVl31UKnIq5U9x3B1Yqg3D3D47wa8JyNDQw
gbp6bGcGRSZQOuQP4Q+77Js3CZu5P+0HWg7o1vNjMh9sft+B0aiD6syszKj0tgMZUr+vrB50OeG6
SqRetmsPyIqIxARu1gSp5TtcWDjLYQbBBcTusFbnomWsccqpvf2SK3P5TEZh0JT8ZNlrG4vw1myn
yIgq7f2o0bMOP/oZgzOGjCkA2bxQPYqQ6TH8Z2d5OPLvH3hE2LtvOCZ1z9dzYjzs0JjDb0N8jNpq
p8XiRf9WFwd5pEgeHpmj/fSqV6sIKx6U6HzhOXJVa2+04VXhMcZj40jwUQ6KUghUJkeL/P3LZclP
MObc8S1zlMrd8xYO+puSSQjcrHmPzBnlEGI0utsZoIqO/aTH7TxJsOUnybvg7Of/+gQj6zLyhJzR
iFsLm8HFrVWjG7TDAr4nFWRhnqlv24HvNyuvqWKDf1/EPB27OPNLk8X7VSkld8Ne8qzQy3p92gTF
eYuPr7brjCtJkEOnEaQrZKzT4ElVeBul25KCeYcXBt+YI/Jm52UQqtC9fTQNytHBgHhDwBz+nYn2
dtsIQd3hQuNWPfOsxhJUmH8bcaN7bjN2DGzAOLTfZ3nF5vaJOurjsyU/n8NVuMZyix2lx8t70JKh
LjUNueJ9dw3BRZUQIp/+PbsgJl5BGgjOhVpMgNWg5yYXEM/djeSClboIloCh3IxZh88ITm2fmFdr
WA50i8gOdKKx684cIJZPocgJDSvx/W8MgOTj6i8RD9uLU6LoVm1VpR63EwyJqYGUREMawx0p7xVU
RsKGI9X++HbwuIIJRRaarr0g5pkt84d8q7fSq4Si7dDYLnBmlj9EUcArI9wefA5k8+TSSYGX6Slz
L7DMN+gIUKBD9cn9Jrd3DhZApJNSV86OiT6ltfcRaborYaNVZ6832mV7fYuRMjjyo+OuDM1QhHNi
sWrD4HD/fTSZzv09+s9SEOFBo3jU3fSU2voelobp6sGQgGoplyv/SpwKuFUXq3mTeHdzBgbmpeDm
bWhw0X0k8hLPaB89Kr9iXrOFTukBMno/qsqz+7FbgOuS4pNOw/BifVQUiGE0zLKH7JmDCph52eJN
pdONH6oiURig+EO8FfDZe+GNhmDqwqU3rMZUCIMRI0G8qrcrv1FPgAr4qonELvUXwn2Ph5/cfZzu
nKR6lLNAvy6HKgkoVXvgImbiWAe5X4tl6d4BuIowf/xuRlFKWsDZZeV3N/jFDTeBzppuM/On+5Uu
WZkOQl9RuOJjCtxSSUL0PQ5gWXsHC3YtBAVuiuDn2YKTZ0EjUVTy/lHplTkn78RwmF4+bOJbRKko
qBm5QXUTUGiPxoJ5Dq5SfefiFxFNuCmvwjrdwtsGYCmpTgyMODxGNC4tMVSgad+VMPRtiviLp5bl
/3y9bSGGh7FRdOmQ6mcj5V+f/KMOYbIRldsDIzPfbmLq9OMfHDxDkIH64+wmYHwRnG/IAEYhfLOD
tBuooxh/zZe9lf/Fxtwh0XHyg3qqgY5dwE+g/gdxkW41OdRUU8/xsQc4P8PFJz/Z0BYBbHNUAjOG
ZbmzBHfUg0pPxdXS6i8SjkRuVFjPQVKq8WSAE8Ly4L0JZz4hq7m4/XIDQ0FrNCDXWX3sEL81ABEX
26v/WEMOxrP+KKIZoFY+BUMNaITHDs8jnpWciyf+OkjhFV0fW5LySMyWGp3ud94u4ef/K/5EfSEC
pySuA1TrY84KBgpWHGn+r/Ua+jszEE/lNRXeiiZPsUiqEs4G87nRpmjPQPj8E8IR6SDcFsxX4flB
JrH4yFtJFTBL3cBvlywXz8iE48zxGLsNOplmnBswWyb+M3xRSOnOV2ruNd7VdpJu5EnXeUwwB0VA
mlNnwk2t9m+70CZPxaH0IOZplFI5CgvIifDXNUt0CqYIvAixTsjmUlpoYcnVuZIqqQxV4ExL7+fJ
rbv1V7XMDFeb4ThUG37jcDvC9VNr8CmtwwpkDNoVQy7342KSpLWmbR0a9vju74Wt8dNvCh2Bbew9
RtemwKqIys7pCDWLTAzhZCsNPqN09PNy7n10ZKzHGKPnOW2tdipOKJv7z1vZ6rQrqGXIl3bWJckt
mP0KdIZb0kfAbqyiyVpOBo3Y6zFGmx8kj7k/jJVjYy2jgGoAj/uVsFZeMWm03n21R7cOYsFgj/n0
Oshjl0+QTfSCiIe2bf0NhjIN3WCCSq3uOEx8h06ri35JGfCyMiQVgbJqhXJAkg082vBCOK4rV99s
kaGWtmAcseRdCrnAjIPM0/c8UxzWA0wWqj8/f6Mqg2xpX8+z/nm4HURynzFqmoDw1TuzdAPfaVqF
07G6Bog/1LN7lbxK4LLsxdBBjGr/wEwdOGqY5NSI6KMKj/gN5JrLEhHYXSEUX8jQChBude1GLF7h
8PbLHMsYjippKKAutvIZ5rDPiAMNbj+NPdlTqBDl7PweeMzlJCBQiEd37Wmh75su3KJFYHY2b6KT
j+4FyW2MIF4LRhhJDfKhqqXSkdJMInZQEwXL8zddOVgvYF7/7goFuUT/YkFWjZpYg30WLuXHiqoy
hAVf+gM1gh59yNJsmHtSMRPKyI0sw2Sx0kc0wmA7xa7uIkqsZp1J2NZXbNl2SCEwppolAyC/AUpQ
n0JzJ3T5qqlL5gulr/2tlpHUD3TbIm/5E3xxrT4RWrLNLcaFojFNxZDxcMvAf8s0Mm1gOJ6xBBbr
MHCBlrq1UVuOCcE1nQJBXdcqHlLoe+30nFet/c1C2XPS9dArmEeW7imh0ZRCBcvWbwOzT/HQ5QcQ
U/1KPY0ZXZOgemVUYN77Tmo8mIxXv0DIz+dDH1QMU9i63+0kRl5yhY8fG2mwTaVVkQakkX57EqL/
Nfv0aospG8Dq9vaXk6jkMC58E6lkC8I35ioCh2BK0pqdIaorS1BUK7kgeOsJ2UVSrAWAUIiroGDk
YkKAR0NWAiAzhhtU93V9fgeQMLp/rwrO6V9//+NncQSIgXLM8AEykEJfSl+W/WGL7AxpJhADhyeh
12jKvLeAOuZreejM7M2P/u5fGQykRy79DsFNAxyer/TCRK6uL94nb5F68WWMx5fe/9NPQVyrFJrE
2PQ1bAvF3S/JK+uYX5U/FzJPcOhvlfxXFcWuWyf/uaJ5CZXtZFL17MavDd3rHQVSMi2I6efZpJrL
mzEC70u3ky+KYdyz7GflSqAyBC+cCdvV7lFaYoP/F/iDImgz31ek9u02N00y9Vfirnn0GtOqCy82
Cn6FlJAxT5uHyQm2CXuWL+PkqyPm9Db4tL0CK6/saVtEdoym+41hXaJuDR1GIIE7dqPZze60b/qk
IFTma6qaRvYW2q/SaU1fOCFEDJGyrVKBZbnzR9fWkeAL+1v5y80qmtBFodE3yidcJmchyy8XRE70
01GRDlxz64xP7z61hTqV4kYZ5P4BdtqMW0Of9JuzXSrtCJRsjjnBIRRbN7GWYo49zVR5XvsZyov2
bs88HpBxk78EDaCEUU3UqREckSQELTUu2iFMGmc/5mynXjEv1Z4kFfA21zqEEyq04qLTdscMUc/C
+2gjZAvb7NvxWNiG7Q8NK115kWXC3dzTPSDZWFlokpYMQD/zfLVj6GZ3bdvvUlnfReIyZMPYF1Jo
jfSI8H33FJlq/b1XHHFc+UEQAxolx4NL5d1lHzls8x1rPTPt9417dXEV5DkMfIrxS1tHGvZizYfA
OMNeh73dKzYi4BZjk8mNQktYeeEpYzPw3AW/IFKAieBbxGSnpeSr26h1U4HyIF/DbLeF3igcJEme
qKpCyQjTzZhoxYZP2URNMW4N1alz04aIhOu+VD3c+6nv9uS9wS0S4ir+XYghDrQWSkxY1uju5ZV7
iAOPtHxNi1Yd31UIrU+ocaHw9Ajwqn8utU5m94LUVyo1BbkgvzjQooXfzR+fLv92CAKIyiGK6Bg9
EoxlSR3I5UWwsEDnheSceSy8AQbtrqFxEn3PDUB2OvT9lNItBs7maiuRlAFzDLTa6wBn8k9TQcc5
6jzPk+qxM+0jDp+EK3R7nLsGGgFpZHW+IPblISf5u5f97vgLPrPU6muDO726sXMlewqHY0f57ndy
LnrDlnUAOsUsf4MmvFeVmW4vKD7bSsQazf4eOO+uhrW5FuFbfq2NLcBYWalNcUvcDL44DwcG2Jgw
Gxi7Os/jJcCPqKQ7A0LnkaJ35WMmtPbHm0BRKVgjXLZ6iwm2q4FhWDQqVNDdbNNNpYFV6Q7LtwOg
UKekTNHW946IJuHtBeqjRriMB5l671Vzkt8hqQ30s+8nktOP9m3I2auws8drFAI3KuPDdtSTkt09
DW5/jg0THGwYbxnrkpXTGPY+/OwH8Q2i3qt8ORlyLF0w0BjuKxWL5v0eJqjxnuDO8C7AxyeOdwWv
GXngvRv2jjOYNwHOLM1IgQoUjYidcHZ4jSkb9Wcztb+gHj2HMDgbsjdEHoP/ytSOqvxVLR7D/IUU
Sa/A4GFZA2FSGWNhhL9XwD9vqk/01PNvXJRA460T/PEv540s0PXzW5alZnqppSVYv9ld6h5ek+ll
JUNnKxGILsSlPfH/7jNe6N39SkUrTSaWiXQxSwAFMbZXZM80zMJte5Znib6qWwohkgGlTx1U4fpm
v/hx3WkHe8Yky3cRHDjgcm4J3RGXSuIPCa2W5TEQegq02gO9wLKRDkklCo2Xb176E9PyRUGvcKPA
0wY9+mv6PgRSN3Ad3Cb/9Y5EGJquzndv8n25GdmwRd/oosO5yS7RsyBSDWy9/nR6BEWkICLZF2Sm
/blHAiHfGMNrbRRLd2e2Rr6h6dKvn0tpyei/O2ZQgiMtHwbdUt5PIoAlr0pm0VefZS/Z1Yk74ET9
6g4sx9EUtGhyqAe+mmOVyaMQQnNipF4yw/ShtWxgT2pLXRAwIInJvop35c5yZ/vMmkAvo4RcQaq2
1tJvKkWeybHkTra/DUjIq0WdquaaX2M6eUOPjDTxuGBV7wxRWgYurJznh6kRT53u08SW3TNKQAlF
KbQG+uC9vGEnwapeznZdD2GUb+6mw9hhYLS8z/wj96SrHj/cEZJQYNvRhTbU5zZvDfwVoY6tfb1p
0NZEa9oWfVI3SwBvl82A3w4O/CwJh9kpRRE9m7Vpw1/9rRx4lnwJULbcJQ2RRZ4LG5IEfULIIGZ3
EFAD/YO6CKZjLT4ZvCJc9k1P+QQt2H8ao5mjebXhjvg5QHV2kBuwUzcFCzICLzXq6KMa6neqPUW+
gUveMJLdrdfvYHhfZBkaWYmrz+swY0t9Eb6tLjQ09pgrDJVd8VXHGLb0iE+42Aru1SN0u/UxtQLq
FagEGTFek8CrPkwdfBYKEH4s9uTAxuHzXAXuiJnjQ0zNkeoYJLSf+XHxdh7Ebybhexkid/1gyE7v
KOxlpilizLRz9qYKv9WYsyEhKHOgaMGpekCho0LAezByz55xX6FolsT/Mm5VRgTeCZpsbggFeLKW
yfSjFzQ96URsNjS6QvXnx27A0JNnIP7klTNkWvYOc73y5lJQyyYNB1UqAUS9tEm+ZQdNecFflgN3
cpYP+7pEyqrRXRnkYnFlgSqecNUI91r5uYj/O99okc42mLYpZhwdQNJFEFnC2516lx051+LO7sJA
lGpH7aFJ8c60CbB+Q7kzD7ew/YIdyJSSPfEe+KUv6n4ws9aIoDE2r7pOvG8X5SYl25wepLjgI7jI
7IuFUL73lE2/+WvOB0b6nzsMw4r9PmmHj47GsaEZyIzNMTDPJt8QBFgT/9uThDqy7F7ZaDP4cf5M
HRMVuY+WQ8fONq1ZF1NSOcu2fRawK3Kw/Thy86dILL6B1FWdwovkOOeGkrbteEUKJJE3A5GR/XMZ
Xc+V+LM7dVoyKjtkO6mSnH8L7UMZDvhOmf6xwRbvmupwVCcCrPqBs3cQ4wnRWEmRaqdp3x2lchKo
sray8a6ZXFpp0irI20EOe9Mn80muavuWg12M+N+su7/xZa8OhNmKN5sZmSjDCpEEKxLzBmQx3q9r
cXuOG4QkX9N/zpmdjSCMEYy0p2uLhSvkkGUmAcO2hhN+BRjmDST/FZf6ALYjCKdmpGjeAkwI0l7U
dSIKaIyPIt8WWJbgbrs4P7YL07bqJYJ/i46rf6Cj2QzK/+cZ6JmhshOq062Bgg0SYZz2Sxle/ORl
dBVHUOhvCFN3tDYgED8cY+30bNB0xGdJI4MsgENWx8xu+xAAIUbm94nKEB+so8SsmjyQh2qjgI9z
iRXiBDFf6xbkhtRhpRJdjpqxR2JNQxNwA8kR+/ky+nRR3vKDoJbK9T31kwv4OjZZOZAIfjeJkkpg
9w4Lhp40X8n5fmV2eE65+8Cto4hrX0Cf3CUgcAn0xsLp6hzfX00mM6LDLNiv4C3xZykiTucqaIQ1
zYennDZFuogbbBY1pe2MD9iEHq88VTUrnzFJngdQoMDe7ZwxEs3EBbwJlmrALCbfpuD2h5sQSvln
kyT6f8IiMb42/27xqYiMYkSXa6uLPEtbNwIYHlmu3axZsIuwkq/R+rqVvK+3IX/RqQzsA/f9I5mO
ChfqlUqZlE6UYjQo6uE1NjPaMCvI46Hvjiz2CnPjmh9Q/h/9Imx1WJ20Y3Bax7r6htzjZi950QKA
2/29d2XSus6dH8D54QawfYLLDlPixhc83xx25lfnTATgd+jal1mnUM9hQpXtBRANj3rUcKUX3nnW
T6KoaMnYQgZ08QL1NiKtaEDBeys3wJLCs/TP8p6HXcjixia7d4xXH/VsbIkA6rbK7EvBG6yJTXin
f3CX+oGmmpu6yyCA3ceK7fw/DYRiumB7QMZGXlI/VnNKXsJyCfMUdFGmKEEAdn1+xpDn0g1xYpTB
iKNaMzu/URqLYCN2toBk+WaPh7EXrHI54cO2d9kUQT3Y72Rc9GDTRooJdanymgKgUOHWLNAm/aad
xLy4yrP6pcY9GF1hx1cCZnJr2ffy7IsgFtbLzh/8PAddU/EFwXt6NMAleDLrUUc3WLA320QOWQlB
Hp9uBPgHnCIMFeswTDmAQVZthQXXUck4LaNlMGwug+c/45mIjU8p5ctvz3kqQL40BBFjKENJiTU3
W3NMZAi7+gpnn4+wju7BC/TaikKOEsgcxW+VNJGleO/zSMlRp23FwHWKbEzzfA4lVxQjQRYegtak
08UYxdO1p2gDVLDjU4JoejxSk0NqUgLJpZX3JWMsDw/WaY0nb+bBWs0bd6GmA9vBoIpY9z860T+R
cyOywSMoyh9aLmz1ZWbl6jgQS+QMbl8jYE2frMCGh54dtbVhQmMt2ayOPsrfmW8mQ6ZPXdtl6gdZ
CsWM8QIyQT1CqRV39NY/KrB5C05Lrm6OGBEdGjklFXCXupQXI73HMdS9xo98YjEDFzbdnJ5aTGT0
7kAxu+TZZ2kWDgaaIFRRB6BXGtzYJt+MdQBfKb5LumF5juZbZe68Lg4j1Mv9SOsskxoH8dWauJ3J
yauqubsMB8yaH0XKfY9EC0RCnwEoxTpkxBB+Li2WlPECn72EwQ9J/EK/DYyGFT1QJWPvxrxlEAUb
evCdfnNVzOiFdk/ihkM+9JHZiMQVpSrLZGp4GeQABCMsJEPH23uYxdOu0Ax/fD62ZFesW7OZKRCc
atK2BuVJ8ktHjEPYXEIv1Ps6eaf67WaGV+jdegLy8iFBp+eJ7GJ4IYE5+uTyHmtHRE+vJUekLb9W
ptbPBxPNqYPEsYsdn2O5Lkj/0PEZjQj0Wdb1yMMxNjshL3WeVqqtNSr/4p6zFDX4FK/3mkwLg0DZ
g3yLquC5rws+0HVYnGULQXMPmY0uomqYCNIE34Rc3Vsq71ppta7ai6r0cLu1r+j0FqkVQ/flMpt6
k3Qj7cHY15/gOR2ZS2RxHSvdsK+XIrCgsUFr6JSdEpA1JHoMDXJJrf//uv4UlsnEwv/zHOULVp2Y
LQi4zaytLiQ1Bj4vsAjV9yzmEv7FR+DagHvACyBRTbogEYarbAFk9zq2ADrZbWwhrkqT3TIpqVUT
/TkJ88zLJW77JaI7NwGMewL7tdqnqwpZ7+NW09MNHR3KSLE546jNO9H/ZjZeql7QnkglqxPx45cZ
DqK1l717fDhHHTYuygdyLWWv9/2aPtwXTV1zEkHd2/Cx2lgha5PgRNFG/AwFZyvEXKycj5BN9qQ2
jmiIsoBLFSoAXIvN+7Mq2gNuLqnOfhLTxDTvlVC15vr+pNKgLEZk0w1u/2E/Z+q9SqP/wzjJZvIS
Du2Yc+ZZFcTFvFQhmkKQc2hGbHqhWprJ+pSP6wMQ3NizRfXi/p57zfrebp3VWQcXSZgs3PtrQhc2
CydGlG8uGrq66+qmkAIV86y5e0U+gaBANO5hS5izXCZ3YFrhv755VP/z39vnHbPmfSQxXBAYjHMp
2bBBiMz6tzu0wJCYy+Autiz7AWjTI41PW9fF4v3SC8xZK9U/cydlbet48EHzgu3vkFtf2dr2QJOA
pLrM//J8vbbkDf6+xPdw+jp7Ym59/+Hs8VzWRBktwoDbPh+pxEvWKlWerQDGk1tiyG477hT0YVyQ
+SI9msmwpA2mA+uxcd+bUhUpQndPo/8iCblPyGAITaYxj5cs/ueCl/ZMLlZO9c/tLP0P9hEcm3qH
lXDAU3ESPbVbi48VujuRnS5umKCSt4UkOW9uNNcc1NSXAdHJU0vcr0CAQXhgIAb/3wR+3kYJMfQC
SwVO5xPJUJcZ6IU6o+uiHL+j0MKkPdOHdc4uCcvzMKCqNDyRrWqspjy8CdBwZ9lwcqdwXw4ZDAE1
t+vxhdV0BFWJxdDvcpT0HVTyC4RMNekTbcMx7c8r/HifHq2IvL8URlV6P18/dK535GnC0nZ9uG6n
EAFp4FN04B/BwBljancRxvMkaCKHD/qhfwQRjY4fTJogRDVfzVUVVJpSjzuAWphzY0Xl/efxYOz4
IuU73NkR0imwaXTIZFmuxc2YYojU6X2k0dclh+vtFz1AomU3nDplWIRdeCT9IEFoQq0+bSA1z6mi
8ceSf0qXbaLNo2l7xp20/4Yk7RJt9+SaxR4CYJseW3X826P8sA8tTykWU8zVREACIuaW4rWaiLSU
WcocRtUy+4HcLvwgsAjGQpw/tYDJt1UKV6z7JCi/KNe8cRBX4aQJbyCP090TEv7/JZjoGUM5fvwA
/DOo2ZWGrku0NArXlByDDYvPU2qo8ABK2bw4sGD+nUJKI5+7gbSe80YvPgE+Dz+dicsjvgjd9rIL
JeHewsiv9zYMoX+sLHl1Zm+6/tYnm4/V8HSr/rMbFjvAC10fynzFBH7OhnRuB07x66hY84Z7D68L
SpSop1Epo3qlQrVEIT84ysQTXJpvmNf4Gs4C86nvhh5mQigXof7KCYGns/5FklSR9jC7rAA54JNu
lxdWydXhw275rKEDKKJvWd6viCKJfXpy1qKsZJ+oi4HtjYjl0luHYci0N+5onuPpnqiA+R5oGNDS
1pBbkQuSEU3GjiosXKXI8kDZLb4GxiT9tJDLdhhq7RwxvvKXRDp5eATL2l//kUrN9Qll0IS0nGh7
u0+QkjROj9EcdSXIMW8X/aMs2rYhGO4zYDWqsqJmoRhwNm3RFYNpF4NqCD9fQwKgHAqxpAqen0K3
9Q7bo6Vhn1J38z44Wntgg69SgMEk9LqHXFC17X7KQCLxTNnjZn+m70sSuCAgnJz7N7JPAVMK+JDU
kAaN/wkH7qk6gB23Up6IA2x1quQ4zcnyyLgSOTqhbnHZ+Hqx1JbBQ4ROApWoi6sDSAH3p7IIp7z4
58UouFs2u8mSkXgp6KkBpkW4ztS/2NZ6DFksybiWyR5xKuhf41YZjZNwbbEWmGi5TMsksK4Z308E
xFm997q8sJ873AkuUOwVG8n/JI3VW513eW/rYe4nFjZmLZ0wOpyUl3c8hEGRe5KLwL/R0Ud6o/Cm
Xsp3YrusIGUU+ZiHEwZWhoZ2XWVYT3AyfOE8T/Ed7KPj5avHLG8OEO2+VXl2axhXL/241pdmG4bL
36Vebi9yIPevrq9pu8XDcCmb1S4/7YGub3VMzhewc1YXf+ccnLUFY1QfiDXXbpMA/LoAzXbTcj8y
8dIBX2F98JImoSpKk8y09cNiurxiijpoqj5RDVeguTD/XNWiSXHFTYf/s1KY319rEPvJPnMm84cp
Usrnav1JqolyhparOiAGXkh01uDEPS/OqHtGlL8/H+kQDqYHFhQVJXnyK9kkwORGaBErZ/Jmf60d
AECLsmUwpznY1lpeqHe5lmsc09T/l9CmfjWuhf5BZMKpEd1Cj2/MXprxsQ5r7cZb10WyvCKRCRx3
q/SY6PqI0lppzdM9MHigi/vSzRmKkDXxrfP42o3YPB4hx3IKLbInsEXCrT8AoR9FaxgzgnWMVAHz
tpX0TEvK3CMA2Gnf+vaZLbrWODxKXApqwhlSGzK8wPQbzHOFrZQLuTfZ3/r9JrWX5U0fYB1N2IZB
mUUBLi5zExRWB70J5HiV3G/3+wZF9X1+4+ysCGMHbpKCVSfMZFNu4OYdlviqa+xhPAW9EAeF53uW
7Ffl4Kzi5eFvzq5z6Zm/TXWq5UshLeuuIuzVkIpyivHbwPdqBrb0pf1TXFkpgWI59PEjBMs8ld1L
03AAqCwFCz6k4YGcQtYkTvqqBs/t9AaaYEt1Vyje0PtRHXw7d+2cV1HEMp7GrDeA22v7u9AMCHFs
FdqGR5CAKUP7NDo2RBtWZVuj3SnXAUdRHJDYbS3cHZeRycV/Bk8IhEbV2p62Sc0P82ugbcKq68WP
DBSNLWvuAso7mkh8LEnsxLpNCeovxmMisaJL+TQRSHbIqXItW+4Y5/5mLKf1pb71UwPZabZvJsGk
Rll6Xngpj0kc24JFsfYL1GN9RbqO2a3imO+u4LyZq/qFGbLoAWzr7SMcm85zSldFnwvphq+jmnpC
QKxl4i2Qh0JiGKFMyYxCo0pG804i1UjZLQVLyhV3VdttAtprPoSk7xodanrE0MIsJuWbNUdjWvr/
kIBOJzkznk/VDKdd81ScGtqt9tuOmaZxOiXY+BBpyd2whZv7DIjA7NtBGox8udCVmdXG8GbLHKZd
2chZr6P9XpaGPhG7OcfD6jZWTRe9U17aO87zq8aJIDqiBMjJ/g7WZ00B/RMVIhTRlLN8caTgFS/Z
UvtULqmdZGrKMqkvzMb4yDpvrZohruA2jE3mMC0Oq/O3Yn0dAWwpB3yjRpVGLqNn0zKqsVDRXYcL
xUXo62WlefczUDEG2djA4pjDwiW/mLnk/PskHyp9m0ppwujxCwITmbCA8WUk+sUsWPOJMZAaD+rS
ogILaLYJuvZ5vnalcdhfQEbBAYlqJ4trc5K7y23YAND2R4+Id0sRI3+Nx6ZASaO3SKhPdthwDgtB
S0/VsduDQqPZLtL+YKd9hLNwgwmMIJJHuaJ1814uSEjuPj6xnulqQ073qNyQEEFIongwznWEyAVe
qTDvxL03kSrXQ18url/yPEGiZiBudez+fl1Fbfb6x7xdrwyL+N1eXeeNxW8kaAs4vm6n3IFNYPub
vxIV4fUbdxglJ3WcdpYF8PrpawMeGDX/43/iD91oGum81IDwW4fs3wXAgr45UfBDfwwDQHU8sZL+
Jgi6zFri6krpR3VoyU5hOHMRCTdu128iVP/J5ThzDpdRaeMuOj5YuL0LONov5n6EsWxP6Tp206/Y
O0xcO13rmmX2LiBjfzQeWtgNV6FXq6Ndx/3C1tQbqbpoaXZQkNlJoBQoOW9SZArXac/N10FfyWy4
3QsKuxTAxpiqfv8gMgxoEZY5HfqN1S80bdZed4w0+hw/kwzQEBQUMyXRRUBj8BeK6cesYQ91j2FO
SaQFR9IQJRyOoK/meYQ3kQvq5NIzT8sFUeoQM53AQ0raJ6++czpdZspeCsCgSJkJfVsU3umfhxMC
JQr90TW7t1ca/jiE83FpoTFD9smbknkLH/LLle3kdJqMCTF9lMfe+ohANFJsjxHOsd+oFJssogoP
wuzuf71VqbSClPdi9mDnPDAxj6Zk7QffLu3ljyp5oFTaYbpgeDfI7CbzZcf6xRplCecdl5d7xw8D
AhKNPiPTYKchb1B0JDwWT9zbEZuzl9BiFQjaig5+RHLn2vho7hG/jGNsKfV7VSOI0GcPM5953UTS
VUvxqpvac4j1bKuPSf0aQWXY1WZaehDiFbkRdGRDUg2id+17kP+LWDgafmu5jrEQ3W61fm48tp0Z
ITEQ42MCk+z0y2b9aOtSbgb0Id+ePba0LZtOk6Zhw3jSBHDjk8IEArLItYVpL/gWH/LSWoDpbUQj
cVq2sAaGzr6arkv5Is4ic6QtAVFpzOSxtuZYe/OKmaBcirn1IxMuCs6G415aPSqqIbCMUbN++9Zp
vgAWg89/oZCSGWVN2HSjgFEAYWWwXw6JQtKsRFaXVYbH031LEtJPNBAadFxMGP0uQLP3reWXxwRn
c+jurZuHCGYEQjjec1yOEDvqgRqquXrcOyTrEwnmL5z2hjpG8fB7e2gQT3ZoKWfQbxYiMbW9yvb5
bk9z3V4d+ZDvR9FNLCE9OOFNqFB5VPWT4ZSpzaddwvr20moX5hAJ7fah0JXqP4Dy7L512qZJvpx3
UwRpWAHqR3jGQf6ujeBFB+B4CHEAWwbzsyn0CSPZSLUWeDZyyduaq3DGvbHbqEC77M5VRosghfuF
EAIybCwQPZAqX97Tw8zaueWFVIpR0PGrafxSkpKGkM+7rprVdMmDP/ePVuHDqyTEibuNAISTNmjn
GnWc4nKAVkQEAxtW/T6oOKeakHi2ZF83JFRNfwMLoSlMHJidFoB9HxdflV43UapRepOxlXJTwhY0
tvLukz1khxOlwMQOMlWj4PAHq4QEahc6xz91E/4SJWjrfXnqsge67J7m+uW3XAZIj3wOKiOrvWl5
di7EPDIgdAh3De3wNJWijQTtgsz1fnZMWmafzHtqfNzWAqEnhv5YVSnKkEbVn0ExSEo4BhXodJ69
h8vUDx+AVIBbi/D4ufI8H7fkZq50Zo7hzqh4P8UpXOKvNqW3E2JbMtHl0CGYUiplXX3rvcyQqrne
/jSuEaNjj+pgFrari8/8JPxzTTdiazf7BSAyGXAue2qR2DkPAcWG7rLOSa8y3txcIdcxqbtpF5Qi
qmZrhoqr7iCQPt+7AutClF0zX15tA+pHcXdCj6NDVhFhMc2rNwN1ySKFKcA3lXtd+eWCwUe3AF2U
chDEb3BftIyu/QPt3YaqMhzUTKmAfQBCl6nQTVUl/kqGlNrP7gFuuGFbUtKveuQhvwbuhq5sInGx
WVXWfR+/F02/xqYd+a/3oGb9/pcuJhADUCybky63PTt5I4DEe4LaNXb5sg2JdAxvtE5THWHgWyQg
YvFisO/45mYFRWfLFGiovRHrnIYgz246sa79NmaM/69liGxo8dWoPrg+3xwfyccOFajm4SuUoTC6
wfZj/jzzt8JLQVyq957Zg/E8Du6XjEpnMPw52pf7hk8YtUNqXsfSl9oWfs1gGOg7uxTFwQlBLFib
UTRKfMhcqiShusnZMkOXRm24jaxpr4RhzkZbvnoYiUWua2hGILQCnMxtq+jheQe8nwdBb5uepWFC
oZmVafv0bsm/TZdZk/hVFfqdN+JwEC3AWOntv96ulKiH60ph3nu8D5Bd7UAH2EhP2+jvkkc3ZiJJ
lKtOllNmPl573qNBlJQLFc8mctbnMSzjIt0lcqeEuxDsTUWvLkn5VxJxGuTTW1PsRZFbwsUsgFfD
/0/zEaTi59WM33wbaZps6PXX39kjSojYK8Moh1w2GFW9occopjROAsAZvl3sGlz5TIJuYEAxb+6E
2qA7OjH5t3fmIXFJ0SVD4RGhorx9j+Zb0xNvihySUJ1eeWT2F6O3xLnQL4LevFwJlaxXx8ZGqdxB
LfPeUYIYpJvdcDc/QgqRp9B7WHRXb0PDRVpGwqWrXLv2vCYSkslGyULjXBDYMdfFI4tnaXMJygOA
sIcXF7S6/lzMbGIbZaismpDwKe+mhZWajXAwmupueOJQVNSnbl0cmlcaF2OcdPTVIrOp8+onDPXa
9W+lXj+rl48+tisP4+Py9LwfMV6neZnRA4WIVKoOe2Hi5AFwHJhf5EZW58VbyH2NDOYoJbxN/6C/
KFDZshv/Otm/bbi+MWRrv3DOJqH1cN+j6xwpFYdjlhGgja0SmOSiw/KzjnnjlT+FsAdDKBJCSv2q
DlIdaJjKRFDvosMV76RfIIxm+mEIUsx7wQF2aJDDjHYJT+8eMVx67ZvKXywdvBqylMpwSyJRhnmY
ZegyvX0HmbhBiS6HLtD29mPliqXR9TsPbGDN2xn7x6y8RjNlcfVZKnRENJfvXS1UV5Gfe8xLVQlg
dbbdE4781aTB+YmovrSM+nVNuNPVvSP3DYp+Khaur9azER/avwD/i9Ak2WCILRK+CEk/1RHTfzod
xGCOXVYSXK6R8OZqISAxpfAROTRsUADrfc0zxOrJSVXidSVGnx7r0yxce5xjW/5077jYzfdgAcFJ
bUGLmrto/6y/HxGVENUtIBXUrq585mb4L4xNV7hdWFUpHYXqTlzczsNC5Wtb3RXif1V/R13KU2Wd
fy4/hLMjcEjyoaC+GmEbFTr4CTsc2+Ge5Dtk1PJl+XaRhXnhJQFf8kkJMlmkLg0QxsY3BCmW4G2O
zTHsYGaVImelx4OK4DpXLCd3ScvOWUeGCdt2LhxXybDwpTXof60BYNRqEIsr2wwA2A1v+YF5Ulrx
TDDNgEHuz2fyGj7TGrpZIAL1FiYdSOa+5CGzUe90VxbvknOVI/UIWMC7WFEUd5d9g+YxrcexXVQ0
9U0z38YqkDlYncOX9T4hgmglamZ8GGNI0wpmkdyV8AokdPmefLnv/cqOqDxarHtT+5Xn+lftK7Gn
0g8aIaBW/VUoFLlksdk8pWZrCwgFX7gu3ApPLz5zZ/f/XisVQkcyXlBBxMe0xzN7nU1DJ30clxYJ
2jmyUvJjdaheAQucBKU/YzBFHGu6gIul6mw+LUKxZ7h9ipcA/R01HaywjRm5K+Dnk54N2azPDkDJ
qs5yZyEgQz//TGH8ZOprk49okyhvNmj/W4gK8Kk+MNk6BLoPwAXRtikNPo0xJ4G6scZ3wzabinJB
2+Gx7ryfzR9y/LTbs3kYH5sphFMu9hYTaMm8cr0vwBTg/B8rV7f+2Pof3n6+NYOcKhhn9AmDZ1vc
WkUYbsnyrpXuHwSkLqyE1p6brVMf0fekXy9zjIalO6yMOngSBka6Z5Q41lJDKXhPoEafNCDmMKkP
bxi4PpR0zqW5geKUu1PTs0jjv87KaDwZQYdtfLkIPI9UrpPmM1r1t21Dre8GB1YaucfdXJlLM0tZ
hSgDA4AGX8U4nPtPjkJowjupu36qyKYpt30/Gm9d7tH61xPaoiyfJFo2mJYRZD92hfuufBo7iWpb
kip0hUJRe6VoeavEetlsDNOoe7YWY/q23ake72HiYn7XoO4WBE93wt4951jVMQ0KDk2LmpQYyXnh
e8wVOygkWqFiuO+TYOd+UjQRJPB7iFuHnkj9qqDq2pAKkweOpni02jIOFQ2dfUn7XTtwhTLZjwsz
M2nw4d74IVYGsnd7Oame35c9+UC/XEz39/hFUcTm77UCl6qpkZAu3qN3PTGLQlqx/XsPjKealRbM
XPKxwO13gYn/VOls3C4cGGVdmKkZRu2W+RcYbCqqOfn8IQJcPr01vcFtnGrvPETtANkiqNOMTZ8w
gAts6IaBo8HoSq3ayQtfg5Jc9UzV5dDYsv/9712YUQSqUMxwFNbB39Vy19J87eQq5UbeBqwAQ4DR
17118cM54qIhSjM4WGO0ledeKg1kLDCuBtsjZgvoYYuFSVJfcTdgpV79LjHVlB5FvcP0RjMMQj4F
H5PK50zjztbu2A1nxPdnbx8WcCX0Z7k3TAMzn4IejiWTv37SKKTyy1o30UzTLSnz5Px0VAcVe0xm
9zKot7DfC98I1/Q9+Ex0EaM3cFqbVUEGf4T2C+Ph5lLuFh/mTsijeGuGnCVeGUIkz8mKMIj5kXAh
XkUJza9xRfpUQQzpnKEZiFLqTFRbZywnZ0OEWJ4+4gdGd+hPKL18C3yg9EvdWFcftTIhWwV303/V
LeKZZmvuncByTQXfTSn12gbwkvEVceuZxC6Eb7Y5tbCI3YHnv9w991tWqe3axbTuAJ3ukoDE1aK0
XcttzgFUQG/3tMrk10pYpmj9u4wrm6WhjOXlPHiKlcGjCJ934jc0+YDh89h7Hv4WJbw68bay7Rfn
bMo7Aj4wYRx9RROKftMldokxDW6Ffoe6GXew6ViLyUvCZITkfW7EYaAzDIQcTRVw58m2B/7L244i
ZTlX4VXUaI4qYBo0NeFtRmEp2EMOFZ4z3RvjKh1Qz2tRM0RQ2lQ2honMaEJy9cA2W0fu+NvUOWmV
fYVzijoqLUKTSGSD2X5CNebGzSbVHcQ4DKyUg/MYOqeeCmLfIKhddGoymWWOz+6okZaogWfdRvMN
HdQx6WJ0H1GgJq0KBwBJuGvDImu0UvNXqbYGtxqIUvrEg6I0OiaJWndce+0fO34syrJdfXmIcjkI
KgseD2dHElHtl0NC0ZLU89ubwjexxZE+AXR9wVrHo1vV6H/vrBpH8te+XfEpEUE/seEXdT9l9lW6
LT/1BygU1WgJsxs07gxNfKw/nh4BaHDANbekLRfws13n2G44eN0xnaEL46ov2bSh2cOdNsdYEJ+x
pUre6ilakmB9OfpjKnsv4ndLZ5swkwRwMCeGAA03iOPvhod93qM5bzMloZYMRUEJp8YjAMYTnk8h
1u2nQJF9fUenMz2KkghHlmzle6ASUIxubZ44GwYNwexLxlWKM24wbVIkNthzrq0JnE83wuijI4h8
L/iJ3I8T38GkE1FrQ10BSiyea5Fgb6hKql6PgrXhW2eTpUx/ssM/9+eB4eYMKHZm7arQT1KOsaOb
v88b44NyRq5KTqd3333NrThqb1qD3r0PswVqwGy4XMoq2L63OmmvWbb3E82AUBqvPLKu9b1Pexul
32bcQbqXF2tgh24Rxqy6daGX7yqMhGhZ1BM411f9drvYwjDYHPodiVYRwz357KoqNsiX1ePHgyYF
lyBO3liTEDthKtrC7mhTov5H5ogTm/G49efAPLfONTOiwPPLH+g9TpabDrfhYn1tnUo8atovXTjA
uhgBE/kBki0PCzAPkfXm2dPpyh7WGMOXV54XSTxIzsfHZyW2nRF8Qh9WjXlssSI/AQ4iGTd/kxF7
Q0ncerNGtXVK6wSjblpcoy7ZLC5NCn4b0Eh+8nCgtjhGsuy3sNsEMtII2Qtd3DRJWSeyIN4LA+8M
eTHpqD4YHtTM9slePf4Yd96/iqpsWdUnzypnmc2LyB9Mj2CmSKTcNVn2IBGsakAxFQMtI3UBb8Pf
yZSaAn/dv4FJm1qF7I2/oDW2DzDZXBMLolSYEx+3TNXR0rjkIkx2hk9bpYPOivCgY/kQ+mPyoule
7fBJWqRr1pG4i49qPWp+Wx/9kucBpFzLvUhQSAO499cV/nkwMq+iJFNd7DNecC3vVdH/HW7jNh1h
PVhuOnyC1QDGRQs+lqW2BlSG/REaTlrljKIlNuVlGlLLBoc9fLX5xrkrMaP2Z/Jdzvbx1fQl5GIY
ewVmIE5Dskp58RQRHjODjrv7X2w/wbh+c1bRZ3CuDlQclgBKPJW718fg/A2PZAcBhPK+xBO0MllW
MObns2NySraHwAPd9u0rVkgonkQbbvTufQjlMQ4wQUfEluhvU0pPeKl0iE/5OxEgaZVfDYUr3CMk
JmmKlk+eoCp4r4aR893gANSfOEUyo2aIrVU2tAvoN5kkge70ZVe0SyMXkt69nU2Gr3adQchXqoRy
SvR8PM+2KmwZ+5fA2b4UOP9gYdVWGj/3gw3FWqI/zCKzep22czFQkOm5zwI/5SkaajkQ+T4sFkhD
YfD/R4om1XHla2MYpGabz17EXChCs1dwx3KbB8ZvPGYjGcBUeNQjp7QCGPHAdLnHlyPXPETK/MeS
ZGA6tDQb+xDtnql43szXV7Z8pUVYwqy2SEXse9uvDu1xVTEOegscKsHcH6GSVOd1GBw4PIPv+g+5
24dM7JiuqzrOAqfMUe7EMrNasCxPsgXuHyDLpxRGVV6RA9nA+Ouj4NGTk/rL6SorlHuvhtsoVB/+
mfhfTqZPCs1r4hwTILrq85JBUf7GAmTixlVw9yvqy6r8yErvxvLNhZkoos111c5/CGEGU0BU3MN1
4RM6BWX+8Pi0WDTGjFjW2mTOwjg+dHIg5ql5CIzjPV5Di9pkJ3S7zjBH9mVxA6ps6uuZuBP3Q+ab
/JwobgUPo6YyX3LFn3cIVstK/zoIUiOHB+hNBi4iwNueSMfnbuqa82jcwIye4Dj7Xsv1iS4wWMVF
LwrYh6lUvVV/SbN+FRlsDGVXPqemU7RL35LjkacNfkIrbzgwm/AzwelDdNxC9REaPsqPmyqvzfzV
zCFMqAMQvwoC+U5xKSqpvMv/0YWbNu4t4vhnZLhbdUDlqzoejkx+D0R16T+96zwl2VKMyt1+xUW3
jfNabBfx74fBL/sibA4qOzDGhbj9Tyi500ZyQoqMCkpLh7oT/vfNcCfkoIPH26SfhuMmZEMGxbss
XH4kZ5usHGBcjgfHW16SrDN0Ud3QZFgizsYLj5kFb4R54qNivBB1Ei7R65Bi9MrclWECoQFLWVK1
pg0nWvIwiJqPYA96HnTw6VC/dnn1wBMesHW8SV8BNPmvu6klkYWqSBLHL+6FCj5M6OMqGd2qKy/e
I9/pFRdrlDTapjj4tuApUKbjhiMkzB9ppqMmfpphdtJssCTMB83X3hjm07ADUqRRgjfCxCem+Do4
Bd8FGqQ3j0/ts6lnie1byU/AvPtuCx9kJATrvSD8GBcxp5iJyD51Q2Q8XlGNa0UxYejhOu3Ht7Lg
K8tayP8obJhzuS97QMmRuJiKZlwSDdhnUOzTvJknbnXXJytzeHkSmzZAruEW5AFG22K6jKeVT/NZ
ueQejBo1Hr787o8BBunvOyxxYGz9VTTpqmDyrQIGqNxVTkHhXJVMJKuoXVHDr3bVxg5wyGdT54U5
5UOMLyhMA7uJtwPBoU5G5V4DpslmZDNE8NJwIn2kEXliDuX0ht7atHIsgGnS1XC1emyuxIlB2sYY
FUf2GXD2Q8TBl3sf/BSJrxQVmo2Y4WMBOdF/z6qIhlbsDoFESzFE110mXY9TsYldO3q+BJ5binaK
PMa9XkuJfBCvxNz1ZybVdEUKVCx7iCw2WNMIiDRNH1EnTwUu6bnoDDVr+8nhS/43Jwi1iQ68VMTV
h1xf8iSy3PxWjFNO1LgyajMr5Zja2lKDvCWdvFauH+ZEjac5d/JwR1lYY/SQEe6xrJUfjS2dF5Zl
2tDgBfVMMD2WGP9GHxAXAHWPfttHsfaWF+kEBgk9ElzssL5SVAxFKkBzwYaXdWH93ViVTvzDduGk
QnxB06TZI1sa8ynu0CMBfxFKYatGNTLQYfM0Zg+4wxnCF/BbKfsO6zIx7F4vlrgt8drjPb6cAO+t
8gGMZKa5MDGGa9C5ILpxlEZtGxO0k4/7pQZojc/rW9ymVNxSt2dUV3dYmPuL38aPlIyZlrDFdyT4
PKb7G8huKFK0oK4UIkK27mLO+JWb3OD2tK77LoNxOnDbfxmhw7b3LSQyKRDP1d9IHbeCE+a3WnLm
xq/De76MV3trDMRxkf1rdfNyLTAyCr7IOwSEbR/V5cggIINI4H1oWh1WNO/uBTXgxCqVQ3/+wRhQ
psop3cFEHbM8Tfp3f+8XLxwLpKc6MfOJjOQjx0+tKXKVnM03VApFSfq6MQUueqPfP4W/VrzrUJDu
ZYBhYeoFwBpiBgUSAwqXucYXppIPnoC6WiF/ui553sNsetAOtW5Gaz2UQE+yp9f7f+gzt37ZefCU
wCXnJj5feLWvITpcs/PVNVWxuTqaoo08ZwznPRclZ4pULziXL1F9dLp6o/cZZWyHHwTb+0ZQ5t6W
I+llhz6dFjZ9V1v4rAY9pxEUH9RNYjdixhQ3MbATvWao+Wkr39O2w45Azg+V9dzpWBRRIGMamjCD
RJg3jKtXGfSWQrnrraBkVCiW91x0tLcI2tRh8+bgNEmS4MlzMG+eSI0MWZpvFAG32OiCXS8dRNtt
NNbHYfBm9qbyiNwC8x858u2GH29QfK8d5XVxEa4/QssPc+OsYj+zKmy8slBnS2DsQfg8yanTRx9o
72dZZ/k7ALWbZadQMaPqL8rYxmMTi8qIGV9WNmkulk4pbwRQQm6GGFJuMlHs6W0BZnQX5mRXSDvN
LnxVRuxQ//W5Bq5nmBSpHwK+MuTGl2kPW3GIt3W5KfCrQUhgUkJ4ouSK1zIp91PUd9dTFishHjE6
cHhz6pR4FcolgZgPlcMnm214AKIftwvYgN7TE3sd+b6Jp376AKjRH2dqrTNRLqJrc9vrtR+/As9r
xgadtNFv1Mbr3REa8XgO7Madt6zXorXHZL0igR+KNbDHZnXYaheOLWYXBfQhXM2CK/j915nKigMi
XrNgtey/AT8Y6iItWMSvyHRNhX7Ti7MPUWjNrD/R97h5q/Ni8JwB8alO5sR0Y12hwM4awS6KJ9HH
sW2iwxyUF6jDOfOJLt4gtG6rWq9KrkuZOJJFmqs607G3p+fdMqlDHnYY6xiTiLbi8dC3oyqBvSg4
F81FfR7Z/hHln0QC7j/4q5DDNC41aGszQgKLjvCWcJ376XaLythi3KxCRKnqhRK5jCK3sKk8i8So
NaTkx3KdjEVGkm0AUjnL8HgXmQphGexwoHj6oCyH8Mlyazwksjy+/PkATdbpX3AtHvKmV/MNci1G
4oaD4zwsuEGGtNiZ2iyRlOpp0F/qQ0Yt6soYXw6LzYztdrTFDvOiU604QEvo7+sKhLKPh9zCwOUw
bqet7zoTeWon42f/N+iMY88DypjotxD60PQKK2XFIp7TBiM2InOPoFlMbuu6DKTHvdFPVOCXh/xh
GVimnlSKobLiu9gENipjtskHXVjwpS2omVK3pd2oTmo5N6b7Djl/Zfy7aV37cd64xeLnvUEAAcia
MISZxurRdyY/dTO9ImkZXGCqBaKJsNW0LGZ8rWvRkbwNXFvZeo8KCWZ2VIAKLSQMum8wu4Ybe+aA
Gt50G+BOxx2UPHZSuAl/5Pd8e2aMqTJGD3HO/Ua3yxNUPtd08c5/ikT1J0N0nkOpN4qPPzbYfUDq
Vqtwnhbg6VB5KiY+Q6z/LpHnL7DmWb2sNnr9Y2vwVrrBy1mXabFPJTCX7Wl6uEe+4K2whWpAZB54
L/ht6miqYSfQ0iparHtDgzkANAnP/rvkzBQDyChJf/jTIDJ1bGU0phH8/zltlvtNmLKgTmp636bR
7csIqyepINzJpEKuZnYk6f1zyMohCyWVeDCvjn3pOTIP4HulP0J1qTRW42PRoi8SD3SulANKR8vi
ktVWJQCTpFAw5End/SZ7h6OQGjHQKESLsTSz/eQaDiOOt90EZbH8duJBl4A4Zefglob06g3zUODF
n2thwN8l1Kddp5eYyJ1hVBK1rBuT43HhrheKY3XwexcV4mDyFqLsVfp6aheVVnZ2iJMrvBJGrgcD
IJYxEBfoO3kmSZxmN5lVEjrbhXlt/ppUaprGOY580q0vGzLM7UzhRfeU6nUvIaRi8ChgUJuM8ff3
XC/pqTn9zK+aPlBnGm2FHcF/A/DE1rVphdea9dNvJ+zho3+Y14TB6Hxj/bBv9pE8Yz6aEIgpRRVT
SRtRxISS9IRds9S6HG1rx+HLiYgD/exsvKrbkZK7bQ7pc1L99g8rdvaBmXer/MVgWr0hHgBVQmq5
yqglsoWQrfrTVrDSVVsUbv9SG7rcIRAOBdcIF5CnmdAQ+/ctRffrw7+dYYNHgCQMXhjp6nMaojIl
hhdeIM0sTR9GKogCcWJotQXQfkp5wa70v4tgGTiZz62sn5WshF4cmh5l2fRoQ3SGMpT6yv2QKXU1
UoPw3ymVZ/ZWBfqJf0/+qHHxXEgIjhOmP2kKIc6h5XrqnGYKem2do6LLgVK0KfnlPPrfsonjUmnk
AoQIJQdD9Zpj73saRCwkGsuBF4d69sf1NDlk4dkFyhIgc592Sgz5yxwj5yKf9Bk9DTQ8TXYxKc+A
rVZNKPpYnEdcQBxREuDn6P0DeHTt/P9L8lEEBLaYnwdfsA/qXQPlmKNyix02s1e0d7gQur3F8ffV
3DuvIzmdkSuDZB991oNZvYamy3rPlQrDY6tPxFtYp5EksM4KYXyXq4mVCjQ6PH5RqMlgLRNCh4Rw
NPzjLeMdsH8qTCo/DAokcBsr/LycQpDUXMZyiKgbDM1yKJifMNjNqnKQbqaAtHcPzBNO+0C3fZ/X
P1wWWQA5Ch4ETuF2iDVZgDuVSfSrHCn0z2Ias1RZp+/NJsyEFk4CNvEwErAkaJqxvMM8UO+9Qvkb
s7dsrQB7kcqCsIFVMAH7tPH8z/JR4Fz5jOausH3NDz/siAsyz7ySIViKyiiO0up+O+zVBzJtDXW+
F6Cc55+rVxU1mCdA7ocO7Hx/cy95jJlWBgCdBMxRd3XYLwzQy9Or242qOfA7I/3MAX9F3oG7xotG
nKZ2sMfKgocrqC3mnGW49VTp/rMFcRzdINMdUNAsTOVZYSjp3AvETszF1F3+GDdyaKn15wRcHqKu
rA/mqwffgXthNmmpmokJBzlFjG0h32FscbZVg9IoE4sZrQ4DvGC0qKT4RbRIyMtRqP2UMsv03vmo
c2ZTVF4NpO5ITkNcrGCPu9mU/tQcvHjK/9iwtXec8xnd3Tn2FP8dZtbgrq3n1ERT6+/KBL8+QsKf
BIBOz4IXjR+8RQW+9Nzz6CMqnO006Io4yakisfWBMETnum8fx1EvUmfcoxUSLtPZVKtKWmpYNPxE
aiA3IR8B0Fke+TRQ3Moen2cj0s15akSQ6yXRq5n6ZFYPy6MWWERTQvXjmh3FwlSQyy5YYwrtkc71
8e5ChY2WqLFLlZUXoHnl8nig9rjPwqCAQsQqf5Dn0kIucqRDELlU2Ma+g16pMEWGx62uLLs2UM6H
eng5OopRaKCX0ORq1vte/B/LkPOkrVRmbGTY9QPzknEk00wls+JmX1KnmHBEzdQxE5Gceto9GJFS
kI7/Yt5cGAuwWTN4eGUEqrWodBorB4T85nDeuyqdHGUJe0TbyL8jqsnSGKY6LNPuFpmFHXey7+So
FaLqWsVu6koEyYXxF4MS+X09uSWc+Slt7TAXsw6pzR9AcBxUI95UteGNpJ0IXibwt3cvnmzdcPhs
z6mC7XUbKIAkdBh0BT+x59tSBfczF5q/+O1Nd8f+TukXTaEXYU8ef+q8YyRvuB7LO56t83sfcOwV
6tulUT/lnLVX6Z+IYqcz+lysIXdhmt16BdU2l04gxkmH+cSpC1dAlDL+7VKgF/r9cYhQ3yVykRf1
rTeXBMLWSvcrWiZfF14k00ReZR+O/08Lm5ctXxobmYTw2H9eIRpIxzviuWUj/VXnxVGW7zCmjJKx
2Yy3f2MCqYWV7m+yCBxnR0bFUmJjxOy6OezKuBsyh6d18YHkg6ow6+J9dr+hgHPHQ/N+yDEKXIlx
6aHeyS1/XKyyHx8BLsipwU80qhPitep9dgUVD7bN/0kErD7PKcLdx00NTescjOnE3dawrV79PbjL
+YlhfurWGvkHQwlofDzDE+ymKKemnEnuY8ks+p3YDNlNt3pWczVRBVRfQOSbKcpfNxPpR2brp9oy
gykz0QXkiAOldAGdJ0jnBLUXcUbQB7YLn7rWwHPIdyG0wAOBQ/2ExFFD/Uh1vrhz5UaDiAVskdYP
LgTWc8WN2qUJaI5otnUhkHX7QT+VXABAbYPFNsSo37e1vjcYCcHy5IsaGoVGW/5wU0HWTldOEAjL
RObYVF7RWdIRLZ+2xe2kJSnmMT7ri0TvHyDbB30/CVZilDfUqr5PWgNDTe+dm9n3VRdZ2cUcFQR9
DF5icW9kZaRHj3fytiTKNTNit9Hw62qobOyieTjBD/Hl0S2cNVjTc34aosl25RD5XFZ1ounNDUob
VQtheXSkpSTQbivE8BDg3gVj1OcJktNyjzwq02rO2+K+TFTbStrQRiNY6KjExtQ8SnHuIpiUVTmX
/7qGRRS+1kFFURu99YrpS812prUg4FSXZI04R9KhJ1+lV7kjC/vHGS8ZNxM9a4WSiK3bkyXl4ZLm
2xZwNqsfJFfc9jmUxipMYDMMhfbSEdaSwtBFvWrGRvWO4Bbp7soi2ttbI/ivIpnCyHDBewDPmqD4
I7YafK4vdcqimpY9+7xGWqhYDT/n7yPkJcUHc52JYYMKucXOpgKB7JfZoPt3sDMb061wDtbfzIqE
PWWMY1G3Zbv+WXHe8LLrkm+u+QMrUWzaqbWPENZq680M56g0XSw08RKN1YmG1jl029m+QiSfsYKk
UuiDWVjxke2m0kljPEPW7GlFoAO5w+kWjWQLJTAgUz4TWboyChm5aT5x1MSVxAtoRNgelqVPVLcG
R1dAG5C9w4o7nXpAVNOt1/+Rt4iPJJeAFI3Z+eto6TxkT23LsxLoUdZ2ZECId791Rvg3GKnOgzL6
idbNuqU4rLC8b54DtoDBEGwT3XhLPjLKw+N1+HOjrUA3ngd6a5SSB9kq42ooJzNcwv7dqSYHK5oX
ztpdgVCW9mRWDf/6KRmu0iTfJ6uF+jFtfI9L2OE+de3Xkj/zurGFEWz9242Or2xxJiFef+xjSQzp
vULqwc5oMKcEa7KB58sw40abIge7FFXepoS8WDo8Fxm8M29S8pNR9VJ7hNWZrL8EC4MhP9qhppiT
62gKRbo8lDHLKZ/OTZ97ddtQYKWMU/RblgmVIPFulR+N0LUOaES1bwvzJLzzM9h0qYjfCdIOZ9da
kol+AXbSX5Sx2/882O8QJrHukFlkNpWvfnA2/ZH/hZR4hjmpk6IRYgSLIuEKaI02mLYHq4w6ZBLf
V6ejwAB6fihPQmPx19APIueZA90XGc/Vu4c7rrWu+9adZ58o2KmtLuc7mIh1UULQ2AUkFSWJvcjz
aEGJpQMhPlqT+xWJDId0e7pZGIcgVXJz0nL5C5bYxBHFKyO3zoDt3j8ojP8Exjtv/Rbx6sQp3qD3
Exjk56uKnunEnxBOrCIc7E+z2gkfPx29ipIcPY0BmVJPVF9SmWmb+XmueXGqNDeCGxaQzwYK65ol
Eqx6Rv9SOFE/D/tDGQsbH3spKpp5kWJqNcR03ZBeztP4Pl+9PAtH29g+mbghLc/6Dfs5CPE0vWVx
67gwxGXZMWnrh8bt/mloOGLavgJtWbqCCsW9ozmNBdRrFmARYQfxmZZJvb0dEWsCZ2vYJd/Qcjrf
+TRWeXO1UlxKbZ+dRN4HxBDj1t6SbwMubAD8mrXXq7LKEX5+WVeE3L+Mt6EFDOXO+cYO4j18ZI6+
EPHTSYqdd0va3gk5hCqCFjTsjCVETgfqLQw9iAwWcQQGcD9oRUqlzZ5/D0SdsijZE7Ni6oWF0fXt
f0hdmAoq2luMigYJR6ys5caJJjIdZrgfx6VU5nxc/bvaBlYRZ+x4i9M//CfPZnPpwfvuqw6oLJtv
SIUPtbJuEqKM+zHI/53t2mVBGq1x/r2HR1VkPZC5RNf2ovL+yv7ECmtbCqiahQCmp4os1DxGC+Yr
IGLiJGE0VhrFNA9PCs/IHs0JgY38yqCdRGxwJeadhMbueSLbQemQJqnvLUV7PjqpsK64QLeO4VVt
JOC8sNbp4tkMr/rAo2P5GNzNL3dF6pt3zfY7egp/HiWJuJo6fF3gMGTvOGy93yBJUqtM3DdgcT4T
pc1c1XMwx7l9EIXscLOE/lf/OtUfnRbEmt9rVQUmM7woMNy3HAiSIgznRVTcJYI4faIma+xk3V6r
1QP7rSYGWTu1ZnF0S4AUcFAOzVcwfJjYmuWZLAmYU2qxRH3DU3MPkz1tNGXgWvYIxIvsATsg1CkX
ENbaKjsiHt4sD6lblkNvyvp5NqKYhRHUqRIy5LCl1S7WW+LK7CR195VcC1aBQLfqlolzY2NMqvM9
BXr+68F0Zj9/nEg2uxux1ZDbLZzaE6sdxTRm+VBphqLfI1co3/FLHZrGTJEWoP0wKYpWPdm/aB5d
PH+ljxGcYzJ+Ppow12yj3u+5FCP8wMjShH7svRdj6cBqQXRmGYKBuQqPXGYRAJVZLBl7xox9irif
Q9guoYsNoIYhhLcryk7nsxIccMB16kA2IEH1Ed7OtDhRK1jjL2eu239y/DCOJpQUEGAM8ZYUk/DL
RoKdoW3XWDlR6B4LFGGZvu47aO6oHwQBjWic5Oq3gvppcsEIOEKJssPJbMX43xuHg3oNwdmqIo5C
dAV+zUbL2Gry9I0H+nR2vwVhDyqz4OHLzv0B7NBOTmh/BIENaLAR7QXmcsBq+ZJTQDy2bDMx5KBM
gFbSYbiso3oc9WHw+NRI34523cFR3pTRfCPpcBTGrLRbz2TP13ZUxmT7qEF3N8iwDHz9aGv+U/0T
AgwS5vNMYravynPOLq/pi8H0BSfWVidjqLDIkVquR6GF3sbkhZwTaXdppgLqTDYP0IdSEJE15LQv
ZOhw0EhMrrqlrtGMdOPUeKJIyGnzmnEL2APfgpdIWJ6NKhtj1+jDgqNonAeQdrJcw+aUC3txQqGZ
6ZF7rucjiEa6FxAgaFt4TxoyUTXDGNVQ6m9Wn0MXMiX0Xl589psoGCl92AUGBWvPx4NfERRHIo7E
dLKFX9JRg7ds8kqSfpjqDDdnLDD8qSD98zp0T3auI2SZMbXqLC8ulVlMinE4abjMwDEYWrbbxJk2
LJc7TkHAXdxF8F9UdktUYaenIKpAbt/pf9rec/5KwkxGuyqJITVj5hE48ahsmztK68bU/23+pnM1
J7zLqJeksbcUA0UIGlix0hDfU23e8Plw2J9/sbH7YE/bmprLWPpbVYTpRUwSStOI5GbE/uh2kYtW
qB5mwwGs5WHOYmBciSXpOxk3LtdKy0RFQbqJN/wOENk0u6AbfZh19a0RmyaUcdZT1xTCpwb1bvJR
ClQd/x32ysQKXeG2HiFjt3CKhek91eIOhbRDnBsw5NBsRDD7Fxhqsp86pRxLTC2vPGwhUR/mbonM
U3DeoLjLaq7pY019a3bRVCXGSIuOgJP/BXt769nG1CaLNmsrmmcwKGiLHR21/yk/EiAQjBv3ewEZ
vRe0G9mZbyuS6biANii7ebwqQL3OubNGViNs3dKmC5fPDPKxtDBNggJC/Wb8sQJtGnRw4Tyy4e2m
wsDzmjai9bFqCsaHEGe+sfWD6ZieOyd0Byfg61+2arTylQg93+efQuknYorU5N2QIU80wERoYpOq
sMzxAlA/AVz8RNQpRNouPLnc2J2XpOIHi5B6mtE95o6y3A7kSnO+a7OXQf7M0JXNeqlTlFEUEH3D
cMmf0jUxGVKrAmC38zc23iElW6xaXWQyIylFLLr2eIgciQU4DuxHn0b9/mIWZxjvG4iDi1VIZq2x
ngdVhXAshXCyETAC7lzrTBCB0aT0rY9N3H/EpIRynYpzoHe5R401w0vn2csmx98nvjToNEQ40FqV
KI7Hvz+HHMZCULr3dvGKV6/qBgpVmv1GeflyZW9xlTpXZaRe6lpJE7Xcr203pEZ902TU5fiKnZ+E
ITcTMMsNqhtgXYHY+GJYq6nfvxIThLkaHB730YWz9hqHPBSg+l1KtmJbkx5z2dZjEoum+L66h63l
r1ImCTVew00eUQ/SQxfyb5hwuMDsv9pKkjaQwaAFUIoAszc0BTodBOPMggwGE9BxNQDwKZkv2Kzj
qW4qO9x83xfIvEPAuzwURqqHwErIpSTRnndzyaQfh2RZLaXzYQo8TzMqm6hMrJOpEDbLzIwPARn1
aYHW4UEUHu/+PTP/dBlzEYg9ezgOOteGeHX1nvAvduFhaCC5DZvkhegTGVxSERn5Sv9SnHKoMJ5N
nH9Rs1cdYJHTjZaiha9pqL5UcCKoLRIv4aa/1haU5BHZQQJ9lzEycCWuFt24wBC86t4nIExXsR9+
gohsEVOlUKHxQ0SPXxoBzerVAQqNHshJaLIQrhMyoRlM1S8Ak4qADjhSZR/5x78QfcwKj7y6NLQo
r2OV6X8wTxbnfQXgAkynaMcOtnwMZ0fk7t8oxXJzyzRh82i2QK9VZ/ripgWPI1WAEYwn4nNK2I/X
TmQSJ9kLDfm6PPMWazJOhM7EXy+FlJ5EJau411ANA0IfMPF1kTjCWRxvzf3vm18EadezPQWeE8Pu
8FOoddyBreMUy+6PTa1+xEQmZlWfB78E8uRLdX9VwL+9RcclALNRjrVXAzvhlKUqljn6nX/Tj2C7
dddiVBIMkGdr0OZZ/IFGss00QNxf8euJR+vHm3uyfEA0FGtUF0ljUAAaITegyF3SOdOVlmnSvB/0
0SZ2PzaSQliqcu8yFZlWQap1+/ttGbx1UPoq51qNhqX5bKoIg0W4+1CVLXzQJe5DTPH1DDe+3nfa
4VFO9ibK6YFgoZpedPkVR9ob7nnNTm1vO5AN7dJMmDbb+1oMPLqKyB9OPbVjTj1iyf/Np1RifVek
yopzCdvU52o0wmJp4Ij0zmhZpidtdQB3x+JiRvXboEMwzm1fao3Sw3XQpj+7vOJtEPyulY4T6Ots
a9uVPbOyC8C6VJQ17o1NOOUpL0FjhCMELpsvDB31cxsI4NUtdZrhB5WvIKDDVH5/3YQVYOLlbNQI
OOiKuksB/Y3FRij3OyulS57jwKb3+y/tq6j863C5EtpgIo1nHKcssH6Avze/FzxvLfIuYE5B1nWa
n5nPfghv19NJhUjedy78CrowbcA1dowVJ351+qDgf/zrlyARPMXZ4VA/rFekMUwKAi9ZjHnUjCth
0zhRsqTIzfhrBg7Hxujlud12TbqVC5n8kTu+SJQD3VG3R3r9qrTNflevQUCgBc2I1kCu+wPXic0D
WxKMQjf96JFC2+jbe7SRQEzWmWsK6uXhtH/WbZ4yxh7yf464C8+x+U/zSGSBMd69bMzwhceisYzP
VVwV1rCIWrcH57DjsBcFL5qwIafhzQ8hdozlqKtaXzZ+mCmOIwIS++lhsEVF6MBTlnuV/XUq3EX6
UW7JBB1+b028OcsY0nv3c2WssltilLfIBGqoie1yF/1P9ImoQm+Mrd8wxX7mcqTdpYup5TgSiNxp
G8ddTDKkowz3fKLmKHeCbR2thfnLunncMtUXUZEmkZdHsaiSry5sNVnRxz/FSuwNJRjK83IkyQeV
HBOp1dMmi/1nax7ISoFEO5lQofChjC7+IE/C9vRl7QAJTM2OKBDgGSF6JXT2CbapBxqiI74P7Ozg
ShH6fMzTVpWZXSomzZohjMOsKUyh1w8pM3rz1AzwMSyhALhirB77P6LPryrh7jaYKogrM5vZzspQ
dke/6MWWBzktIYVtDCmTQ0rnO8HQY97bvsQqsbkrRxqafZFTFZBJiT1N+kL+9C2KY14gw7Rl/2p/
uCcGDe1287HltRtSb1QzIW8Iu3m2ZIiMrEIXyf+Xg2ZBDqOY/JQYxWFoAawabHKlrM66Y8qNsSWc
Ct2Ok+undW0vwfKVBFuM8IpFbfAlAQd1ecyWS+YVCjMKFKLxqKBNWIxLNL1Ln53t2QB6Ey98YUor
UBsG5mZemyGKDveTPlb7EROxRFjkL24KeQY9cOIjfxDBkutpxv6KrKWDFW/8OCU42h0jtR1i1PJQ
qnPQhkm/dONa4UUaCfvsaLWJxicbDhqYM4/fbsgyeJ2zFtU5I/yI2x7DlIEnxFca5rrBLMqiCo/b
QyG36VrKWQeBzU0tDPgUNYLxNpXhNbOCBAprbhEu4561Na227YVaEgWTJ5XZU/4i8qAMD0ZqnEEB
ftvRQwRJlF/B9Uxn4EqnLtgSerZrft0ZcvSOjNmAoMYu9h7is6i52JlxRZBjiTkq4ek4v3aaatfq
OeBKJ6QyvloLwR/LB1Ni/MhrN4ui4S0wSM8HmContvWNE01IBKnpimQdNQvn5JFdtnw4UvPLxT8H
NJGkmey79lDo9oEyMrs81r0uDcJSypnngcSpbn5hFLi7RODAqXnPVMxUQwoNqLFN/4sGsxc6zD/B
sw+H9dQZgoI+mG7lI1JR4/uP9qm9LoaekpTyT7Nj4WVO5xbIVyMwM+WVrgo9bi3qTNMTKtdFihgp
BlDra0DQd3zBNhYUUz0qvCXFOCbOlof6ueUkct1nEunKqmaYF2vZS7/GiAVn9UWqV2SqxCClOalY
dy6Ak2SZpcsEqyoLTHhooJ0ZZcTyIvJIh2gVZovdDq2jWhtzLV3k+izjuAPbCY38a3FG/NRwe1sS
hU4XiY+UYIZ9g1Ht68fgOkGAGZnohfQiozyVKiNW3B7WsviWN8PautFBHqZkk+hrvVSJTv31Qs5l
TOao4NOFvnL0BBMNuRClQTC0E3b5unQyhCPqvEcBBwvZuva4sP3mPBHMJSze2Hd9HKCfDfFYA/cZ
Q8A3qNUVyL/pPck5EUyYEuqKc0czcx+h4JbHVBuWahOu2F4EGux0XDFJLF+Q/A7Ov+2ZjrPfL+dK
doPnXSdhA0YZ1tZNgXs7pzTD2xo3HKxw6LXDMnCPKedp3OIoGMepMiu+0D3szSZ8g66gzLESZqFb
1iAQ6YKMCwO+k9IEM7fyxLCXnnQiNsiuUwaByflobKCxyxaHocakwucY9N/wrjENAdeP64SRVcHB
QmS9dR/XFjvbF2hVZtjZVjWSt7g67Kqqfj75xURtkEML3eGFuDjvjVxDRjfga/b6lpFUcU/iJnTC
1uK+Fi0tKKuD3xTgxWbhza3OKzGEPN0PHL9z4Bt4ktntaZJHS1yUOVB4QccLfhvwg51vh/bIA/Tt
oDWZrpaDnkPHnMz9qj3a97MnllaY6L3CjUckvA3YBvKbhV7tMNS/i8v5FNOJ5vZ4JVdrM+Gr15up
O0Cb81n1UjAu14f/CORl0kChYZ7T9b5ArmRP5Tds/i1DtNrSsglI+ft4dKu43cQbqVgDsgORpMrL
0GjOvHIArsqzpIbcoCLWlPRkBgy8vXsIdsRW3/lHKpDIVNoYWwh2F/CnGvmZqplmyEv20h/k41iq
jk+OqI5GrjNH8CLoHCqsLoFUZCZYsiHGlKjJrI4xNZmdwT0Ny72QYDdx46HBwZzQ9lHqsJcbGqUK
4rfgGKIsmmZenKQ4K/C5ATTUNwdNSdiSfDVg/AzwL1cZQ8k1F8e0xqq2NcKB2V4P7HEfEMkdqdmn
fUAHNfynZM6z0iCe7TShSB6xnaqFn7rTxKZAQ+g0lBFGTxmY1kNL8aAxw9qz8xXaMNxEQuFlCiRg
65bwfzF9eta5SLtdEW2Xi3PY/iKfDhOQ7rx6CKLxvEE1mQhyHFKBn4qrhNY7yK7jsUruwO/L43zk
A4iL+hy2k7gstAwZ4LPvNVRDDPKZWulZytSHeVJEQ6Hg8i5AyeUD6DkRME3soNmP51xAD0dv7Ul9
/dyBm1WPe+udq5xeVfWA4US9pAQGtNg6bISZGGphw09pj8rZ/MShLztDvyy6uBjCZP8q63UJHqdZ
ZPTGXdJKoiTEr2HLugyTe6OCj2EnF6SCmuqoIy1ONEMO8A/1SHK292c/jSfyyA8WmXAlO+i7VxGC
xHApToHa83aV9qHeDRcDjoiJ/gu5077/tmD08SuXocGfnG8KSL+AT44DJJChHGJY8b4IWku9Qu17
AqEkqK973iqW7ZK095SpoCGHskbB1TsZMvL3JP3/7tAh/Ej704fKMzP4QpEJdivsXg9KeyLTEVhy
jVHDMevwoyw42M5rOmboYegg4Zhw2kOFKIqUhvXBotVmzm7wRYtR26kLT/SM2tCMhxuD76BBWUWD
ZPjDRLjvFYkvsh4SJmfAzPLSC62gh29ntN2jhzY1HXIgmpB4wrkI9snO0IVk7PzceFe7Y/loZ5ED
a8cwN4NbATsqWqqTjo0XIs4eRD7PdgKpByCAc9GsTmLCvKWQJkzJYfceYtU6yfY0XGZt1oyRpLmC
WVDF4nO5BgUe0/F2ccc7ATb3GYjmM+U3ArzUSSQr2Pesvi8pCrnV0hXWvEw6dTSRQhf/huFArg3a
bIKnt98GpEF8pGzvFU19nh9LyTqc4BrMlcPIXzz3o+nTPcVgG9lfLjDVeWRLNJfcSITktM11YQvq
TvQ6r7KFm9XxY5LU75HSW3UsfjcUp0zWXlfTAMSbKqRh+J7Fg/V6M6dF3iJtup/Y4gARki5H2kmx
Tb00amwRq9S53MCCudT3cqXEL9OiPk7oiRiqrhtOfm6gYLU+b0i1Q2GheRE2eNl3+9pvNs7Pfuz3
l99yzhRGxvNNRjiRfNZV5URYXJQpelOmZH3bLC79SE+PEzkfDZbPZn2IjI+1c5gHjytmypOkAE7g
2XZpswnzcBQGf8Nlu+x7mhiwhBHIjeJ75USTYMA7CJdgSzmnpF2yy3hGJ6lQjFRyGymuiMptML9w
LBM0n623hX7+DZvAl7EvUQYL3WAIkSCvBxa33s3/t6uQHn6DKO8O4gmrdJKPbrnJPszz4lg12Ib7
PPAVtla7Wdpde1Ztsj+k4kg90K9wPt8XiqVteSDR/OpOOPDp5C2/aEejN2JOeXIU7ZoPq9zsPdWX
6qyhcTBwvuLw+OKGxVV7xnxAbIPzi0N3CayCZN1ssHIp2ZBen7gWgU14lBpt/k8p344TAXb/1FJd
1XbY7NshGenh7McFHwVHsCHcK5xbiZsbSYr7jtokYcdfgKU6ukzIyvJlgOH4WimR0jPGlPlEYTO0
CSdho7C/t/QeXltHjLnnOPZc9B369kNrFJTGUmrSym15IFS6nuTAzVoBEYv5bDyD13Ba8+IP0cOA
qm/CukOM8b2y3Fzkfi/4Vr6oJp97aVMyVaatQJopmYacJLrw+2ErJjIocILMelRchMG+19G94yF5
N6IhXX0rP0Vfcm4Gh87jpeazdtIQKthYO6LhUwfYuM+7Nx3SlkQGwiTrnljqsRKQgcB2E1Cqyyeo
wMaoYI2rUNFEJpEg3BfOnnbU5IkApCAKxZYoW1Hhh0ziG8cK8ZyhjG8NEhG70qyVodIvRilW7Sv/
rioZ5miaLoy1kjTSbF33pYfCQdk8LyekNL9YUzl0tg9ZlgbYytD82bgP4/DER3rcJUfXcS13PgWQ
F4xtRxAxah8NlE0CABcFX5ptaHkGd5MCY3hHP52j1qxeQgJc8h8/NVuelOSWR8RMkXMXaHZLetBv
B+vMgH6h08+Jl5hNaqL4blEn5jBMDbBeMj4pL01Ko34rHJlOAchWE18IGmOBr4LvqF8MSwV2LXmu
2ZHq+xmNatjpqtBW5NBpg5TUW6iOFdhuiDNrYv14yX7eI9eMV+1hFpjAglr8Swuo9yegYQibVSBz
zVS1LmCJ+VvbOewUe2xEBBIw7B9Q1GSICTs7eL2cMzKSscS/Ve6vh1UIIvah53YKN3jz2wZDNExg
sPnv3IEZPvWzaRjT46KAnvLdjxbmLEFzUa7ETf0BN/2za+3oQbO2YlYIXuEd+58wpw34PaBIY30/
FEvWLY2Rwio+zDDBPHHN94tf1Ywx9gsuOOnoUYSaYVUMNkIbWzYQG4TO/+SXgNM9X3GZsi7HJot0
3zWNvv8Ini0f+3mRUbNvoMrehZ7TWI2NX5Itu9FTXNWIIz0I2Liu/2rfeKwYc+HWOAejdGet/Wsk
ibIWq7MumfRl0KUMDvjYKM0NPa1t0ejLC7Qi8zpnaaUJW00Z8ZnTtErcyw/B9+QwFIMcJ2G9wTOX
lA4AgtWo3XNHDfNz1uc0D0gTQyn3GtjZ+Fhl+ENHCtq4NC7+MpIoXlnKHrKUVW+zFLm0rtOQSPhc
zqHqKMH0AwnSvSThv5zU0jTOlZlRa3PC7xf9yZfWaEcSC1q2sQC9lxnX8RyMmKmdcQCd+C3v+d3H
SwSpMeTKaFIExLC00Y9fHUPKtbn0TfRRxv2eGBf01+oBCSDTNVNvN26Ug9g+EMWCEQt71HYHkDx1
6eTypDkxlIUxlJ7Ww4iuKsjH9zy5F2IKakBX8aIPrtBD7DxqaM2zgpG+YTAKhLxvD01Yztc1nvgM
3Yub12ud4bLtz+lL8dJVu78W0TBDXnjgtLQGwAzVk974iHlJ2rzS8E5GPI045e2Nat2+b4KBFj95
MxCnysRZ2MLrzsksKO5Nq5V4nui80e2u7u+QsVIIc+xyYfc7Wo8KpU5hW4wrghMPzOlB+uwordAi
WqKC72Qw09LcbMQBgFaS7MLAGd3b3lGu0vWCgIWHT95W70n4dETSlZHBacSPFyBInzB0Ap02j568
kqgjpVhPbL8vaJOvKFMWczMXDrvXwrLFYV3HLuhkQQlwq7XhWKrzLbBgGpMZ3N+IgjEWJKGheQIT
MZY/7JtcTZLyC5h2Tg6LLXm0rZTPRoESKi8Kwl+XGRjCbYcGDCxiwwgJdiCGThtCYfb0z8bSN5NL
hRXlXnmMeb8WRDc1UEvpJ+n0XpWrk7G9VI24vN6n1ztM+njNhACQt7Oh6/N4/TkwG4qTw/tK2wL6
KykGW9pAzd/KPtIhMNUL9efLttkYcy/CGX2K/CYoRiVlbVA+V/tR41JG74NUOi0cxiwQbgBfnP+J
vZYCWQWGLacG/Pgabr8xIyvcWEM4Hu7InUvKeFkdDzazwjXtrIxkMI+eq4hAb0hDBjILhLb9G3sK
g3hDZLcHUhfZ7BfmqBjGv078hDTwKpeNdhV2XQ9a0IzJpfwF1BLR2vRyYh4VF+KC169AaX8x+jz/
qCNxkPgqZ0OmGVtxyas+ECKf+SOmSDe+DqmZjdI0RcdFsq4tFt3PfJ1C01vF7rVPjTWqxHR4Y7ia
foHhi7ySDK6Pb8fgT9mpsoZjnpOAy4P+zTHugN26E0/vW1JOtQ0k7i7fc/EUF232aAdbJGzcGv7G
K4ObWc/pUuw1zrB8mVrMWqhvUBmNqBAc0alZ9Y5q4mUu1iFbfPzkHzBUWAuxDGDoVQumXhSrRaHy
1pjCEc/Bb06LF4YCXMiUYHRXqOTZK5wAnY39l+jCDllMwleOStAgRDwRCDk5ycHB5j/ZvAYL40wd
v4VKhPCfSyhrUzB5OZpaT8JM9Dg6EDvUaVeMXbLt6cdBhNY30ufB93CVmD+6VVv1myWgnyLosre0
Ji2B/H4q29lxb0gX3JCB3oLPyv8+0mELSI/TODnABgqlEx3jtD+RP6cGDF1EddIpLe6+rvzhyUXt
fnO49l4UN94KamXdNWrrLJ2DORgoS9xQtlMbNCFE8HsoJZPzve/z8kvZl27AJtq58sXgin2YQhdW
LiOrPGvkCePM/q07jCPREZKtdJ33wMmuyqvpmIikN3bteC6et+Hy0wj4ygMupilgDpiUNxjIkO4j
Y2x8Lmi93zm1HoyJ71pIyf47sYvMFrjdi90mUoUoygPpUDGkQWjHSGu1/qzVTDIis8UDZHNBPF6b
hoqjnogE6SBw30C89XDdi/Cz1A4CCad5XDvMf5uTlv5TswcSuuRNwu/ThKjycyhbfUF4DI2a6FGu
B/w5HjgJuk6qx2kxEh21Vukd149TVlnlwufoBWJGvtng9gHKsi6eKzt9syudT4zeBho4cMW/Q6hW
Vj2ib3h59qr2x6bXXD7nj3qnkRH767ohUqBmnu4dPp47fbo7yyxl6IpVvfXu4QXNrT/8bEovwfvO
8XZK6AQ9cKm7sr6FpbZNFix+0dG9J1tLliX6q2Nlr4k1ac5OOSd5sQ/drTERaxF8pStzkYMTte6N
6ygXqtgcLH/QQe1Oamuax5ZDXgPZxngoymfNlW5D/TuHNXrnsrvNcxH9a8PRlE25kyoM1vYETVau
szfYCq83/KQNPGKvSAp8zt0GKQxegF3DrwMP31cBKQkVjSyUK6jBbFjzB51Ls/GBU8ZOqQ0YLavh
6gSu6MiEV8HDIiZDuJ3Sdvf8UwMVTgMjNkQ0kTzPwLXwj0ZLPbobrOU4QiGRlitR/fvpCrcoV5sh
kaVjHAfE5irTbmGGTxudHKaSnXD9ntU/3vUH6Okabuwh+Btl6KnMX4wDVQhrxz/8IRToH7Go77zj
VPbgCXUMUt58UeqcFFtCxVFO2MnJZ1mUL3knLYp+3QG03Hr0zQwcgRmN2+ikoALm28c1fSAfRHe+
roHzJug9VOecndLyV6YooqzX+MTb8Xq+KyCJNyFnC1X9jjbFTHkM2haECb2MwmGVwkMV+o9G28Pl
FvXA8L4HNBwCfFsJ8Y8NkM/B1Q/TY/Mzvz+izMSUiz51akFy/t2RrS+dVkJcjQ7vmi1CEoROJk0+
KbgbOMVKuEppO10+09IQMvA9/etW5EHBxy6Hw59JsJebBJKGwD1PLpDsLkE8ige8xUlrnmeNdF/x
YWvt01VYMUXw/KBCtHcDGDTGBz6pykenupudCsU3yHksAxOhGLN6ngjfGsAKIykAemzSH2TW4ZVF
YV5o/ftnzISh2w+izyt65cGhlhA0TgiYQQdcmzCVo+57yS+gmlOTHDroy9Sz87BcrUFdSlv5RDJi
R6BswTq8nx5cn+1h0TVTSstCtGbYWgISnGumD9kS4o07QCvwnSbxq6fCRPSU8gw9W4QMII0WFJyi
dgjbR84dRsNiU7OyDIbhG0BOXMz3Pil4cj3iAyg3l8n/EOlpWRp48iX3xe0rxy2ULwOlm70TxUUA
gbAFFWz90b1148LkdH9OlHV3KFFka0vpLeuwh4NxtjrEjwNwOM6NpdM31c9M9EEfv2B1Smzo3iew
/DbHK3DBddwEDljQvZkToWBvpLjzIMtwZ1yTNtAjCWIwX0bF/xXyC9dAXT3rzR4zT5klD0XseL6F
/vmxxNByL5Lp+dWhHXe9Qwz77rx7CzolkLedhSfewm+TGX/TYQJjfZA7jWR/FxHBozDBM5TbEZeF
aqhtb6FAksssD6pV0eQWOmH/StQBzqJKjJnslAO/t4sv+pvZZNyyHrTmRhC2CPzlWk/uZW6UCGsn
WudCdN/mClFw6SA3ttBqzEhPYxFTyfK4zLKJ3FPUUan6bd0XZfPxekH2Xw/rrb8VgS47voJUSMWs
/ABWWL9Wec6us86Y25WlfT5fQxwJwaMlC9T4rAEr2xZ2pqEZomJcDS8fxJNWgnkPgUDLLFfmRJkp
pR/s+IM2Op2o4FiRY3aULlCcopeOi8Tz2OXJ6d17D2XE5wCUwubZHTyXbAjiZnxmQCu0qlgf29ue
QlX+DKW8ShrpSXMgRHL802kK/A1LpzVdezmbyC3t/ZN89aL0iaHZ85ljKBouO8i9aDwz4CHdfSio
96fNAtVqJN+Nd9dlZPpt/qv5zdYtPN7EB+MHZkunFCM2HvsGrGS/W1LVG6URhZdZ3AVmcwqs7X7Z
ZRDjeRwawdX/mkxngrr+4zqhG0v5IJCCGKMYZDt5F0vP7G6WYZIs6nxr5uZQ67/I78isJhP394My
GM1GOuUsea9D0BdDdAJgCay9tqUvflkuR/p+iRac7fDEx8kHrhiXHN9l46f0JdAkYkO/kqGnvBgj
eYc4fQ9vIEIUJzJ4TpJNU4D40RgmKHPRDVZFZTYHb2ZXr+0RB6MvyEQLl+6S3mCrKD9Ea6F7ZrMF
CEmeQfcKOW31vqjINHpMwNTBUAShMK6t4GGUVvqDsS7OBmDwQmljd5Ze7KBXnhevs4gtbfrTaXRI
0u4ItiatNEFXR+APFVWgLma82vKTrCxuVDBDuT0MpfJgiNg6lNOY9It1IXcvrcDJbu55K8siV+0X
t0PIqrqD91Btvf1wpDl5TVaUu3BxiItk8k0pclD1i/QzHVN3ozOeoOK5CWyCf23vAspr0Dkj/HoR
5BSaSpZ5fwc9sQx9nKRIlYXV0f/MCDz8hpjPs1Rm2sBLWcxWkib6fEZLYCNwy+UVWFxPMgyI9mEg
hNh/nBunyI+k/lsONxbwGguuojpLnmzrjL5GfCdUUK56P/WuiiSJlF+lMzidzwCh6ff1vQgvpcLl
ylc+Y+iE0w9AF0/+aYnJ7XjYodadgt0hHS57Yq6w6+zha6QWT5B4+nI/BgYsptwsYVZTVfCzStnO
q8VGpTUsjaV+iHnLn3BeORYf3JNokMkEMFaFuGhJxYSc93BpFKvHUGql20j6u4rN/UNwFV+PI4lG
TFtxonv4abdqPsemLr+7QwAA6dGbZTKLFG0AA9R8xTYOe8Ex0U2gcu4Zc4dXre//HPcmvBmc1e43
N8hnkyAPj2qJhBwlm7hmnKv1yl5BK35GdzxPuFPnetpDuvZ7vxLqzD8lHS0QILj5xeGWCSVfkx2E
0LpOvIqJDkU5gt4I5BKQgLd+FklHdl5bj1sE1fjXZX6IyNudyQzyFpUbyqwJ666oQXArG8MnoJxq
If7Aqm9U3JCONT08o1ABxINhklXUWyNbsfrtYtE9WwBWnXrqgnGFVx6FW3mfX4TSRSRniIOBU24/
9hQ1gJCxbfn52VRv17D9N09ggK9pWRaPoul0qFxu/EdIJJEcmjYIr2H0jhPFysjaAZyaFk+u3MUF
AF1USGiuGCX5j2mpAH6ZCZnGBvzMeTqDLg+XPQfJXi2DtJyf6YKeWg54eC43PxbRW3knPQcP2FDt
bGsbV+FNbu1PyeM4YCr/qEbzgj6GC/aykK94pC7Pr6X1UvH6liqeKT7+uGzHfmv+5/Tv61qfdaYa
8HkV+gZ271nFuzis0JIt6KccdNb2YEwc1DJKrUFxV/bvs3MrkqxeiVRIcvHAFd0oVfRHG6X8JJcg
c8k0db4EtmzOPR2gi97RiD4+5i1aWfRYqgow5+j6xJTYtscjcmVZHBCIYTP7wovPccxicfwFhgBB
4DaDQ/Yu1V1/BTTKlS+d0j7djCVO989zCIkMd+Tv01g8OxEgdiGIuo1ZGP48ikjvYC/Xb5QVeYzY
nOanOvqq4biAeGYWiE6qahhPFUj+BH9/Cm+z6CBKH+LgXTqHFVAz45AY7ROAo2AJXVnu3ET6ofez
qgBIdUdmVM5QVzemSc2tTyyWaum/KAqI1jJRjWSFJC/H5R9XuioXvdhAfniME5KYeUCiCjUx5z0Q
xdUUGloj/R/whd/VLCHcTK0JPTvrzzXc2BLGkwaQKQGajbzg14h7yzb8QJ9L5UFv8dMQ8yI4nZHn
qF+NyXfoit/hFSnEfk+8FjptuE6wtNNdJqsB10nXt4K5eLUiGWtAUllvcQ4TCMd4YbpKDP/+nE5+
EaPQH+g/m2uz/ebRmHemanqkIPKb9f0PgSNJxTIKXeoT5qtf1v7/Hb2Nnl/ofjBw+ftJbhywHYBq
W8DRHqCAnk1D6NZbqHlfcs9lPG7/Lpj86w+z+UnHdkDHkOyJdytiwPP/o5pJUzBg2VR9sDtDmC2z
71TrsRkBcEHLHz0YFLygTsDCGMLl1mR9l+baPbnxJzGq/S3sv19bOPxPwoDU035zAIzlZHgRYLz2
2I1UpJ65Q1aE6jh4LvnjL4OIAaQm2BFyOqJJDB2AfHI9TdMhYlj/ahRPTMjC9px8bG7eHCHh/3C7
AfrPcRbylxxIaxkBxuTVlRB+RulDNLQ9nUqqwF0uYHj1s4iiG5N7e4H/58y+LvSj0vyiu2aQnvle
EENtKVzXlpw+ynbxKaBbh5t+jYlq+zNYUZpYPZmLvCm2Nw0ZF7VzFY25vDCOsMhnuKsKcpye69q4
bwq230UeHuJ68uuGs/P+KtWH2CUYcBWrMacpG3GRVm2W6KU4YBTYXEN+TRnkXi9Gkzqey+DuutbM
tABXZ2tL0bnaazfQbkjiJD8m4GG6iGPA44HVZP98gFtdQNLemw3qcqqWj41QnphEQOX29sGKieF6
PCju3ARUuqRGIjqVjXHDbp8dBd5XCbPwhZVdUmh+EmYSJAxP6XQ+h6BxucI6GsoHJfbLG24T3tGD
ITI2k2Q3wgl6gwqs5pFvRS0Z5JMJ8akHj9tFT54WpmiGiPKnwhnyGOAukRlaOb5/lldT3S5Ce7kM
taOp5/8Jgff+WWX+Q8S6Wvu3UuTQ47r/uup/0yIZrXZmcsTmSoJg2UhaKN2WwGV/C9oW5fErbzm7
x96F/nIDIxDBdgresOr6+2xXGPucZY0wn0e8hirEwYz1Y1G4loFbXgBUw6n4fJnCorm0CX8JCaAT
8BYRJjo220gA24DKEXxmlyk3t+tfauFP+smAzhCWdrQaTS+FeS5Vz0EebClei5DTYQncLger/ZMa
brcKeOHisAwmfMKZrZqoOwiv5O5Jd5sOZ+X1bSTZ/bG9uZLv7/MGGEbsepbRJOEerAh9vWx61hQq
81xFJaQENWfT9yZal3ssVE1Is8mk6Y6YPeaMFwVjQ7cYZ95JTeI5vSiq6YHBV7eT4/Z6QDi16iqS
V0LMWWxwOW6GOA3ZrNG91vM4jjbTv8+2agoxyzvVb71m3N98gMa72ODZOFXOPGX+pmjwliOWR1IU
dyLCLoFqIvRDFP2SuHOGjNl/2jC68CjtMdShnBB0/V0HlfJaGgfW53QMEGnRd5axNbR3FOV6IPKf
zrwxo7DCudCSR7UxYlBGZ9mq0sZ3fuA7gQJ7Qc/eIhTgjEPcxkHietpywkxM5m5Zy7ousud3+j5P
Qy2hmg1db5EdCwyuR62SNGXrqWwEJhsiOxmvaXBaW9B0KJKK0K9mLmMHioPjossmpAAqvQ9inx/O
NN+C+96AG6dLWAzhXhMuM3LSY2Dwg9b2l6zSrNDN7ehYMVWLIplzvJABcd/8cz6RklTWyw98znEI
ZvNo+wpnYvrBrvJX60PlRpzgHg4CoLp3s2SbJr9ZR+rbJbNj1X3k/ImOMoHJRPDEioPX4/yz6sXm
4ZSBKkc++cvdS8hRsymv7MpJiYHxWQSJY2mG12JLQAE8E+0lw8CoMsFgpNoAfYPKA2CViF1zXbjf
3qHCuubDxaOArKN3f66MVHR5tBdu8TK5lfNq7hQzheimu8LCdivjjNHTlC9Oo+17mHi2WVEs+frL
A4vvtoI8q4DpoENDMpc31hcG9Zv3r9+Az08aVPTnpIwYkNswnQgGLlwna9x3OEruwLf5m8FFMP6Y
x+JQm9SrLNcKBvKLEdz/XoHDRpVMhDqbV8TqberXVk7Lo8lqWwtny4YoBuEaPS6dudm3NNdSkSQ5
N+QVMHkC/NiQEi2RX2Bfyi5d12Iz7ujqlaWt+VW8xYKuzs8WWpHk81bAGTaSCyO2Let2ACOrYgCg
bmVZPWZEiTL6z3BP4t2x9YygAZf/ZhJ6EU44snlM1rvH52/Ln1NbHBoAeqj+7xv69ZeWVTG/A/xu
kQXJz9fRVYjcpxlfu24qFVKOapA4U+CyWx3nIrsWkGmndiZdulXHhlPK/Pq2jnMssPy73dRNGd5N
nDBlm/T21EoUWHQ28SQgCHi4NYUXCL0G/ItyYg+iWe4dOzGmLZ+2ZG+1aNrKw/JX4CLMe4P67RDb
ZptF3HXF6PNW9GDmTkH/Iw10qvuYSxocbWu4YrvH/mR+N+ICOr2tLA+km1Zxo6d6lr9XRQLdsLf+
Z7hIb669e/8Ue8BbGZblGTvr4mU+b4YRhmaOl+q+sqKTAStGvLKiXS3evcbRgkHknPG31aWCjwS2
6zHd0y9BORhdwmZTy6fhQahr2XZm+NwOs34p4SPLQK5T3PPveB73O48wnOoqhllt6UiznfylEQiF
Cds64XkJSpRq5GJidMhP3Fzel7n4r8h5Eon12orioI2eBcENt512muSvt8+E6Delhk11Bk7vCEK/
Kljn3REQBNb6Ek83abEy4tOKQX3nlwQdETv8IpcwbEmnHKKWWjTsXMu9jnNRmvKZihrPmMHXkMol
PlgKw6a/elM7HaUWiHtXw02ZvrSbVHoR0g85KowGt3FITncuHMb0FBSVLAn7lsCT8SVZKDznNd6M
1qaDllsLclA/mrwxhGdmYyPtpbpF9vYzByoZyKilwdXqDNPIPBHW3vtKZU6LLFPMyuXbOcZ3z2vt
cilqfbbzgszg40v06dB9/KTQys5hvksWQdGJ8FGL6rVv8gBlKBkeN+eIcT+wvLaRqW6kqhmJZZ4q
RV+5ZZaO2mSz+/VDOU2/8UYk3LX1VFQUOL+MyyGILP98Gr5HBOMh4IYss5yn7g9sg1wMDLjySfPc
lyhA1VKVe6nNvl2S7lkwxYEIOz2Bmdlmza+S5cwyAqpj+YzSDSC4Q/XbzgIJtnUS/tm4gStJv7In
pE74fA/URfckoleHPio18KjFvs0MShbbfxPnWBzNVX5AX93UIq4jxSOZVvxR60GQ6G3lx41VSKgp
MBBybXzeluLaB8nrbRegFrjXRpQYtmwmyBfZaK8xqv/Mr8RDgOAEfD5ouO5b9w5qXPTMIecT3TKc
Ge00oRME0CwJW82J/K2LIzhkG+KCpdh6UBgh4qNg0vE9t22uTbJUVJ/WsENLn4z/0MMeQrQLalb+
aXW9g2jdvhkKDZ+8ZTqH1NpEbrWOc1+QbrXuVoWpmgn8t7y952HICUAJZ+9Oy8hTp71t0s5CW/bl
yjFZ5mG1alNuBeDXLpqtoP5Tl2lMfytzYrd5zUdcGhfNtbuk21uCLdXTCz5mZjME1R0GOGZZ2AiY
D3ryA0GQAy9O/T7NQYYNaSRWXJJS8xw1AZ/gE+bLzWWDBNKtE8C/DzuLFh5aYl8HyYKvYhniJyzv
wrK9LTBx4qeha9M9PE73xEx9ZWAxikPLrAtTgJj3zplS1y5nEXCdP0sbNcJdeeSr/81RnaM/t9lm
m01diA+gIYQAa1WTTzzeHZhqtC5zV+j0tFcEjmayIeCmS5bnGlTQ3wnvsnzyN+DfAoeH3Y3kDj6A
D/MbApSKnHAIzMm9IppmOaJomG16UCqs1PcEi7cP/GXvdjVVlcplNGK2o7+stV6kwOgoe2RLfpC9
IngUDhAopuTXqCa3QGJLvlVRphzXKx0uxmuSjdW0l1dGAy0soQ1EfjiF7nUvjZ+ua1F5VW7mtY+m
PCQNyAnWTgneAMg5qJb+bgzTNaLXzU0QurIFLXrqFkeokluHccp4Pudf+U8aqRyDnPdpQ2bUy4zM
RurER1VTOGB9q7yTOAQRB1UTiKipJkUSglq/QEDL3zivG7vyWVOidj29uiDW38vKAIo0S67Tqqas
chOxB/yS1i0q2WsLEKyDQF6ofEU1JZxfQMU9hMeUnSrmmw/LJUDRmCsFzTHdJXhR/fQaQiF6xi7D
IAOV0gEtwtsonfaKTFY1WKOn9hd4zufVf4idVJNGa+cM2ABMQ9w5o95uE8tldPjbni5CpAbY8Vzc
R+bSL6dHoHofZtiVJQ2ehwRuOSr3RdBD50/iWXOPr/XjPxGmYuPA4JyQBgxKnn6lbx8XEYZyyeUn
kqsihvcqbPmdr9BFDvKDLukZNW7nOxc5mrJcLpghoSmDPNkjNTC1At5UWbDwwGoG+bywzHLCZAAy
205ttrkpyeD9UaHNbWSL5FP+rhdLSz3gsrSGMPC5GZgBrg8BUMx8d97qOlDK0tuUBw8j+xRMXa0c
iW2SR2gmp+3GOdxXnt93J1YelW54ukhGdX/ATKB/fAykGrBRsexfCNofmdRGuHGHA5Fp6eMnrRXB
0bWfShFGqSVC7dsz0wuIc8h6Bw1p2AaEdCGxlF1qJZqwRrkHlBpPZv9HDfQZSZr40aqV7rwdNi2l
TULMuDo69phASfJ2JknD3ZxmBd2oW/NDXudQehZE0tdegrnakNFcK2M39aTfyAxgcNnrz/u18But
K97YEQGQtE2GnOdV4mXcQejcXhPAQHwpaUo2FghkUlQpHMvrBVUzQ94hUcEKoGIztQO3dt4GyF3R
F+wxbt56o906kOsubI3htucfoz76j5ujW7u9hGcXhE2s0z8VrJGf5xXdO3EpD+mxf97ExBs67Y2L
bIstagNT0bIbsFfQ1O+uQ7yFhsw6XWJFK5wfel3QzHzPecGv5YZMUL2hKQiPkWCGBHoXtHexVklY
4ydqKo4kQUbbCAJmJc/JdJ9R/GYKf+wWZHdTeYMqqrAsCCdbGZAVZRyWJn0TO5tIxremSF70kCWl
IXEqTu/7D1OzwWRgXLl+yuAgnio1TzPPznUcFOYF2iXACfqsOFYu9vBJsdqUpaZ+wUbYVhq59fhR
WnGp/co3DUNgb9KXppeHJhvIeeUsdCUHSRcZrmXPmBHQeYpncfii3BRw8WWHmz+0FAOZcWswJ5Rc
AIuK21lWLZK8eE+XwRMgW86GUTiz7jF6N9j7WH94jvRyDWXqqlgR0Do8e83iIXQvAaBrL7AKosU4
1yO8897GKvUJDPaqLYg1xPNE5TY4epml2boqbYFVqRXUKyFcmSuW3CDkhWlV033WquVWDvb2mzQt
S9ejRmt/VVt84/TxvrrsrkZCYstyttUl1mNo2PDTEn73CIgc4abfE/tFeKwLhSNUKzwnpE07dkvC
FvkrJMl9ouVGf9UdYNsu37NIFBZ+OjxNWQtG592VfRXcEqRvWc/E49eqIIdVigY0WBKO2jdkt8G8
vJn/5lxSI8puSLeqL7y2Q1Ifl3/wjS1vD9uoCNTG3YgfyvyCFA8peJnAOfYrwuYm9CVxEAmhJAmn
YIUz4yRwr2uLMMddrq4BEy00ZRKu39WEfLMEkTaEPm9pzDPiVr1o0hCMXagigelePfz6CP/M+o3/
OlR1orES+scP1Ss19NuxNjybGWAs1sxLu69EObTL9fdB+CW0vSb0+8BRi6ee6ogekDeY0NDuntkf
Z+SHWwaB9y5XC2CkOTkp1oOg1D69BNiIguWdjkZe57F3oy9feudnNIBQvTRaVCPUg4/rZMcut8j6
tlpgW6nvm+qKLEzoYyvOVLY7BWdMexz5V3ZgtGCmbnkXjgyYFYQhAjbsFQy2kycnJ3V9EIkh690t
tByNfJXH/qLay3Yq409YDdJ3VbszQzIslrnqr7UFOe/cLHbmmPHUY6TPrhwJD9xr+DCmsLRgra0w
EB+j++aD01MrsLFmG1+sftzsxocFT4us+2GI37W0SF2rAFQ6wJ3VaaMfA07+4OjuVJFqlDnxuVN1
jZWw8nv/9ekyUK2pD/hFIm6v2TtM/Ra9n7K8ns3sApSCWI1GyQ3h2h3NShO014gg+0I5REgDEV+E
v47Ti889H6ga4WSjmNpF2NK1DdMq3EsyLCCBE8fhx9QRHcIwKt0LnGbkJ9U7R2tJCB99dJ+1//Vf
cA3nK4Ch/fNN9KkxtxRQ7CZnKBbnQ9QVl7c5o+aL7BuGWRUyf7l+m1FwkqZTyh/aFrPfgFUJh1Ay
aJ6QujnVwQNpWdyOEbL676FgMLc6y2Qt89T9Bt4SFPAKcj+rxEjxCo6o4eYkLVRD0aX+6o/fBqJJ
MBUwerYqyfpHp5APZ7HSHbhZ/lGSQasLW5mBE7moAvFeHQ2r+2SFj1Ph5WviCCK3BRnv3wthzM1D
PwbXvsklAW43MAG5E3PXGdUbJIAGtkTkRHpfaUa9WdOCyhhQ17FcvigyjW1ab7u6qv3BAxBQT5Jp
FDDUxPad2XEmJOHsBswHKtQ13Mwa0wQvQNNZBpbi/Op6iNIKGPXUPyUpfyq5/mwT1L6VuS1d4FnC
t2vql98epBGLTKCBgs3qLVHS9J9zo5PjUQxB+P46wKwi0rgdcpog1aqa+Krk6nrtU8JO0FYBT+r8
D+7H+ooZckugxZSFLGU7dvM820l+FdfpO+TOHklkF64EL6o8nMVKjGSq6XuDmdKIiT7e5npRyA7p
KFO28uz8qIS0U8StvsQU76p3LGSWDuDNEZ3H501Z5VlS3Z+I10KpecE7JMHJbLYn89fGt4j1XnoN
dFtvA/1VxXGovDVAheX8/gIIbt7/6/OJqIhEevD+9a4XM8aZ3KVpErueTDBOfnOIdyJ1Ki4JLamB
nOPBWKretSxAQAMripubUISbchZ7edo73/7erkcUdB9wH8Zb7ud5WMksu5RLtiqC8PRhDBuORzIX
wtttd24IJ1RQqcPdINuawZkXXcyn8FCy3VKMEUIijaRzy+jqgOslZFDBMz3bPxPRnAHqXTURp2eJ
p+BN2pnAx4m0uZhrr1jyO2Ra1eY8FS2sxAxkN9G0S731SY6P+yEARZ8uGV8RQvCEkMajUPsAgbO3
rR2wUQVpvPKardlJnCu6J8UXcgZ8MqbmCWPh7t27+K17ELyXVySW5lPH7tUh8occRkvNkRHQ6Epz
z31CsjNWKQ90vUb6tUPgOimsT62q5fqroyrqi8ZpSX25oyDqBFOyQi9BLS4NTCEaggr2D+3J7Uyy
ciNmYVBrHYtl4s1sdXM9gvPSyhjfWkb3qg6NvdVZlX6eN/g62J07CnhtGKAgCYkzx4wIDKWsd+xn
Ws4n8yQN6fkAvYWQlQspoZanc4pt5eGAoODP4hsmNg1p4sA5og9fohYfJgbJaaHLwYb3LKSn2bbg
R60MtYw2/z+ooFm3si+VbDqfDwcbopv5AydGay0R2ebYI8oqfCs2Ak5cjbe9E6Lf8Zy5zwqJK9iS
kJ0tNrHRai2fX7TOTEe1urt+yNV5daWjVu89im2mbPYJ+tXnedR/Od2F4RTXI0I+EEzv00LaN9vz
WrVozxMPyKHxNSJT1V/HekQitpZXPYDBMM5bcyXrO0QIRR4CK1c7ztxYCH0tZcXI2H3n6fLtI0n3
SglF8EkukSH+UJJBZkc4l5b4Hx8nTWLpMhMfTm1QtzIv8FFud1DaM5XRMn5Xuzrm2WHhh85kA+9x
Vx8CC/ilhuiJAU3eX7j+biYa2PjuotbXr/FUdvsEqQApdYwG56x1K1bLgqVWjDG39uK+4zyVimzR
9q7m43CUcUKohHj73dSiEM5kP62DEgY1+kDlpuhok9On+ZYMFY0lHGDTD5sLhj/p2SuN0oZoFA95
cr8yAjjJk3dkwp5aRcoUzu066MIF7b6Qf4ZdQbSWH1IipiOXosdPLKIOg5FyVmnMCk4LYTd3BNUF
RW6lzGWRW0RBEjoHXRLsWWVYtgZhl/N+mKoRkqdhGGDuahZVPCu2Jqas4UD12hfAZQ0/YS1vX8LB
Kap3ZIcD6A9RgCA6JCATiSo2FNvM35+sK35Dk+g+vKG+9zKdWRZMb+fGZ3EGkmLoZK2eY2e8ge/7
4Am7FbMvyHpuGfVdQtHiC24y/o/Y0SQTjw5mVSxyviG/mrHOCcWB3gyLsVKtEBKv/OGjbDghXXvT
NBiCtTppyO6J3zR8ssCyQ6wMCIqN/wG2bD5lEoQ85fOWGRRG14yBk8Www0z7X+VVhkGLFAWuZcZo
PShtpUYRbgjCEPYN/JUn+IzvN6Q0L2ZrfAE33BXUaQKDVnCbSMCcAzokGOsQULgNhpH+MnL8h2nP
CirHfEvK6HktXNd5ONsNNOokqYo5XzEKcv5+7vhPQvpAOCMy3pQjssnHirYaYgp8MuPojuUdDdbI
hrHaRJv5aMqGwygDqFqpYPxZrQOqTgDlEJLc1cqa35IYtqAGLotUmKrEVtaWAbi9VMmHoQQ2jWTX
StDyP/z74ZL7omS9t98Rt27QU7ExcLhMl4zb5sm+DchXDzX6oKZHFSILDnL4CWiKsHzv6AO8O7dU
mGcjpSmtGTZ3YDTiKpS0lo/4HsPyklSkLL/JGP8N1t56RMvgzf7rjCho/U+yrPcHGEFwA6SnQbV1
Ol39DMyzMKu5O+x2uBEX0LtZb5ksrldThJL03gVQjuKvtuZ88PBEDjcx2VkBdH8qcJg7t2rhJCHv
iYRriIoR+6sI0lAe4S9dIAtvro3EmqDXhveI9fSa2Yz31Hl44BVH5fWjRblO2bLaNo5uS29hp++U
j4q05ZjCJQZ8YGgY2w0X7J7EtZ8cx+CWYeACMJtakNaxqMecggNBcDe1/X+OPAmRYXJuVDdVvK2n
YUyLKkJK/NcmLGsDajZp9Wr6wQ3bajXNo8Tog9wIyKqZE4KcNYgJm3ItyK4Kgm41ZcgKrs+AZjmh
Zta6fHe+D/kLUxcteSB8Ro7pl+kj6HnvX+1jvCb6duPE9GR67wuq/x7BeqYSFHm9rxvz/AGY8BRj
rFUHGFOiRUWmOkDzIVmZ7csKaDuPw+CFh/V3i8M8FwV9YCRAc3jnzY00g8yyeTImI3EreUb+azKP
veZT0tj3ON4rTJCMs3Byc7KtuJRdd8UEmXcYAJql+0SOwkRMsCUnNWoKgughPkRn95fwd9xWYypg
d9h2sf9qVKn2z0UVgbjhCL0tsOGjF89PaA7zY3yn9PFSD/iyHwGuciKa0z8iisIehokX321MrCTw
6sWZ1XYaNEEKf9EQE+3lcoa4m9N5TTxkBHKK2fnxH9Png0NhIIBN9ZxDqPTw55BL7q+ZC+e4r12q
7KWK4tGlgwVq3QfTodkXCpJIH3cmP/ZYCq+17tWKceezEv7jVibV7+BfvAIYWqRtrV7R/Kl12m9r
MLbgudwlLP9Z3otnduPsQidbx3P0cIj9k0AfTZZWvLifG5GeGq0LKfuxsfGje/6+Gq7JlOiVmfd/
6nfyGklF3m9qjgecGZEr7jZaHtDpz13arJxQTbi+prah/2OR8w6VHAdK/n5JNjsNF+q1FokqJfea
9jQ67iDgcCtsLwEZdDICIk+1A+x8JyLdrza0Y9XbDo7//XrMvEOVcoEyEkLN5b9d4klZ06zKYDSt
+TMitZt2UgjPNDPpBrAYRlBaNk3w7KoVbHdUwgTD46MUJT6Qe8xSTxWzbObBdkhavood3DyybIbD
+pQ04tLm9gU7hR4D16KBseG2rRXBNiG8cNsq1Iu1s20wFSWh/9j4CYh/icvNTBUylrceefoqObsP
L7ou8rfXbzqqoZIEW68BbjxDoVIjM4o95XoHBYHGyhXg98oMcQOs9SKiPamcEVFA5RcS0wTfRGIv
7zHMpTD/MATRm3WPcxa52/L3YMHjA5iFxaK77/0jhwZlRdUzWeUCLgWtG05+IbMAnS2wHaAzl5g5
0JaRfvZ6ylOzwocB9H1getuvvOeuIyu8OEkSzvAtKQEQcrni9jEkAYiut02cFgcNlQL0kBq5NnbO
SHnXUeAFsBJ3WNo4IlmITQGDRLUqlmDmuwvj2dPA9mm3f+QxaD77QKKtSRBFhbwrtFuGjKwwg8A8
7efi1IVfXC0KsHVQ0DHqJo96+zO+aV1mgNmnDSuJz4O7B3hfsghx3HbOz3OiaMcjT5pGbjJIrYb+
N20r/RrzjducfDCvlsc3kZWqOg+74vksw3mEU7zEY6mWXE0Jqa7500aNpDBYe6OVZlhBXnonwGJY
ZVayr2sSWU9zvRPi967XZbocREr3Oqefk+auQf1MCZn0/+54w7TZ0F+z5Two0aeElbZFoWUAv0rp
o4PhRoH298SlC/2GDjn4d26WIJ/xFxkj5QIA+4ZV+Y5Y4z3xrTnrUj7aii/MlX17YBzp8+R8QOaf
9olglDin9lMKw77+1z5sPe97j7Tr9/u+0tdtZXmHMMvru1YEU+vqMUnssgs9MNAvOK1w87fKQ+dx
yBj77RZv/p+LZqlLc8ORVlL8rcOrcEIdj8D7msaBrB4p8phVLySD1TSX72iBof+kn9x1b7MT1sVK
NLoeSyx7bqYD4KkdxOr/ummZ1bmZ6ba6nyf8fcgmVbXPaj8+sAK3hgr/gi74YmGtMPRqmnjQAfxk
jtoyuax9L584Fr0W4Y3qV6CLYp4jt7j6I0JGxoMd0Z4lKcEkmMwVxzBFO6ghPKw7jeMIMYdVPatS
rsnj2NccFDhzCq1NObe4qAtyBipw0RfYY4fh2B1Wvwd4CcHrh+nWebMhFQGETKyvLjn7SVJHaAXw
3ZO921Zujfa+CEV4u8gpaN9tYU2w2lK2blPQIhV6UcjO6aRuC4fYQovPULUL/yGmttLiWYeGTq17
pLmd8PaeZYngifO3UA3CsACem8a6yPtdHSOLJUovUbqwaHZxMH4rqWgahBrvTnLp1Y/OBYIePXZy
tDpzNi5a8XCQQEZFEVU4QXddlvRQE5WRof6DxQUbkLv6BD8/gAttYG2qffjTy9NMcIAEvKq1p0AS
6Xc0foB/8WHUkCcOJABMqkcTHfOnhtUkYRwgTz/NtryLF7bQcjMfXbERGQLI7B45TvXHxBeFPyHJ
9PK9yLlaQSgmesQnZFaOG3wfbwHuKe+D0B8WHZW5wrKdAd0GqIVMnyvYt+P771TbVIZ/W/LfJFaH
SS2L36Ok7axB33cflfE/bEZ1QeC+VwhFpc1v/zBdZwjpAhdp111tZ2rtSR7/u94Ab6e9QsOW6N4V
09ZGl8ERzfkwYh00u/qfpYbxkvO0Km1dxOS9us9SpBJn1HJDdPWoowyEUykLfJjKxR9WJYkCEfl4
zCyxysnBJRiPhUGqh+AOpNdwsoUToEWA2Mhyq0MWSrIOif0K/7nYvmDgGq+dMzISbUAAI5neT1jl
q96PB0O3hUnspYUpSFYOYGPCa22ECyVOOjIMTuYmGav9aXE8VoWgeWRmNkGkLy4nhK/CfSS9EjNI
0nPIHhzruYKMlyGpx8ZlHCUTwxeIYeudUi9ft476BpFkRcYyyraDvINa6l+ABUzd6dADInC79RDD
2o89BxT++tlkqy+IipvF+JCy3bdRCkbyQNDBp7xQZhnwPV7VM/OzZvK/EveBc/MGICjO0wZoYIiT
SXqnNGXcJ7CnXAxOecj99CsbxAesBHjqK6jY1wapOQBpPUY/khRvON0WXIOVJivhzSsP+hTr/xA1
2WeSj2UnwhbSq1hzlSWcOvB0UDLM7P5p6EzN3bXFUPvrpbFED9w7rKNRLO67X0T5DwL79woC+rX6
uH2ORj4v1TRAX2ZrhzWLv7u7GkJeCwYEhVoS+tQyNntPNgC+xKh41IDhJN3DmAlli5y67eE5FFiU
w3aW/qBc8viuQ7lIjGvzrV9Ktynb12xtvr9VzVx7G6MjLh5lABmN1ReLgnezQSrv1w/pzp41kqZK
4shsQD4eppFbAygXEkNI/Pqp2mE576UhoQIEmO6jgRzD31X2F/klAAONk77M4Zyx1jkKxd6pCiq8
++PpTN6D9nZZIy5F9laMx8bPSn4mRr70F4xrjRxkRGG3Aowt5J3QWOZcIdgtpa+r8jGF6Msganh3
Xvtw/Iib4d0F01TR7GZ8MhYTMn276dXeL60AovIlWuV/FCsYXOol/Gcq5kqTgOqbx0MPp/csQknf
CXCu9yWgEB1P3eT7uCFo+6WLLE2MSwGsnfomHLr4OYRw7L7qr1mM3HzHf0fUJr0jbnLeqlADvwku
C/wadgYmdRIaADv7wYKodvIpxm1wR3eda4eCbKKUBMIcGDnBOWrGpYwzb95/1t+02HOwPQTMFtBG
mN4Aw0YKFvWqh7JqhJJ/JFJHYobt7/PaBFSaHieAZTBEG091RrvxzVsiaov0wdipE2+FZVF4qgn2
eXUx8PKflZ/ZOk1Hj+CwsdbiGvtu4ARp2CJ7eHtGey5a9z6mbwqZZx/jcaN774LtNUdPU00LMGp5
pHvaHSUU7mVkJ1sk35QbH1sjDvUNnCSRKMy0cUiAj0Mls/PAwIiIs5GhV9EQ5vb+t0XwR9Z+opGI
0QcKwcqmbkHUXdSmp08PlbFfZ6MMNJlW9g42Ed5DaOHzZ1Dhz+9EIJtJoHCHyKo/1211rPwZh/0z
SS/NicMG+FIzkYDcusNqpOgxx+up+55nsWbOw9SyO1xG+MMSJCacVmaipNDS5vOp8VFWerYsmEmT
4zOLUpahX+OyJJw94GVjhzLgTDQsiU7VS/ipqMig5U0hWpE/D0z+2uJEo2d1pv/JeocE7ZfJyIgA
lZMSar3m17O4ERgUi2qVDGZkzpQex3e81DzxGAzu7zZ3yZzLwWgxYNgBhfVIdFEzZ1Zyj3b3oHeZ
EG19JHz/fnZ7sZ1qysQV9phMJh6kfaSArXHcasuEVk5CJgXAhHJ2WiZNtKcG6EYGMVqLaIeqmWMM
LQTSquCDJksYgLBvtqZ53VXQM9jWUOwTNCiPKkb0QgSVOxb+vgJ4tO7W1gKZ2URqBtQ5qXN+eXca
mKxCC6G6OjyD7tnKWIKuaAJC+JaVlJR5gbe4y91HLuN+xjnrwRLfQtZFv3ssr1CmQWxiwLdBaSS9
pthAuf/6y5MdvtFcc5a9x0gGg7QOojr6PsCWqMNgUnp9IZsER6YE669ms9xjErLgMin2AS4ops04
oMDlsJ+1I7d+8XFDA2ZL/Pw+Y+Fz1NNQamrOtCeHgdYZcRu0j8Z32MyQS0u40tmyAE25zaB365i2
bZv2HGQ2T9km0wOubE8ory132OfEjwyG637uRwrIHzPqM3wewXqgo3v+Wz0jtShKDOzldrYDM0p7
dc8j4vm4Wib0Q0v5lWE01uHvPJF9JG0nfsP7eB0UwunVhctPlt3UwIgCXt24R5FZsIZYv5zOAAd0
Dddt78Qbb4IwG9PNSncyxsoabka367aqTKXRAsHqGEJUr1HWfoJZFx4QqPxYM0ARG9B1aC8ph/7e
koSpiYDu20PntvQcfaji94RZS8fdu90yWdpTz4To6cIRrerBxOiT/l4O3YSOKSexsDitcNSNRh8q
CtlVqYqxcStQ8esNzvwAOHnvIF3t0fq8fnXhD57eYoZryy61eY/Q8plgCcR/BtVt5mQB1lnaLjMx
9KBvgiEv93ADGED+4B2axj72E8+YxvoLqLdC6HaPun6T777Q64KC9XrAvS+IaSKLpfJFbrLde14N
G5Kb3tbMksBq/5pGIfMRiDkxiQvq3KRaPk7FJVf1mc6zg9FJHb21ix+tMLQY1MtSnEOMOOJ5nu+F
sY/o3+rSyd5W+/zvrHheALoY+IJRKN1iecsOqGm76eO8REGPMSf/POATZWKtgaMyOfB4cnw3U8Mh
xvFVsNLBp/JLaDWRbArQjJeadzK8nArMO0s/4ifbV6S+cb2lrH7tDZWyo1IWIoA5IZdp9SaIq0zJ
H2lRfkObgbzDneMcTTdK2musTnyVT+7MMGncNuntOM5RqLEjX7enqybJk4SvivCKwtkV1sFVqMZ+
3WNJ4wSKLA87YJ2G9Uxk4IO+u09ghjT2pzdGxM+aYiFRZ5KLVchtNpU8NnioICY/w+GlRpEtmInv
0gGxgALaTjeTDsQsDQExOQP0L1aep371g70AnHkQR7hlTZPgnNS+XI0d4uCzunvpL0Kcyy74uQhi
npNr+aQDbOgareSOICFMoCErFf6i2DVCXUaRz0jd0F2jDVO+k+K9BICYY0+0KPv3uRh0XPr1qSFP
QW5zy7WkImdXMsw63J5TjfouAhoc1uMuURnbL6SVztAKFirIAm1onPNtH4wPiIQR2e565Q1vlbfg
npxk/RBt0jiuFDNcLnY0aBS4ntZnH95svWeaLhbKtRiQA5HWjcrkNh6NcNjhkv85LDsCnJIVzHyC
I62kZZ1K/TN+d/6FGDASGHEvQiWmRc5SjXnNhCoD8zzKq2QUXFDHbF/D8L5qsZiszifvwZcacnQz
IVqnPENqlQo75I5a6UJfKvkCtEdCpkKeqsnCWnC+Yi1Rxq2FcDmXS7ALkzhVWdShsGe05v+Q32b9
7H8Ikfjo5UnGf/Dt7xY5Eu6K2mVkOGASOAaqgPvKws7MMJZrT1k1IMZ1AGoBwzg3KDaKi5ZWwTFT
mpgeLasyDfsTDdQjXkQKYf0TghJWk2rQrsNCscXQMI4hojjW/fFxcKV0CrqiyXLPR51Uj86GLIFg
RmMuytXDjT1dHnsen8VuKVPs+29mqdd0o+hqNXKdBnm3FReKVMcFBqYlVoFFnQSqKS17reObJckp
AmgaGL8FbpfY8eDWg3F/J0ZMRPrVlhEPq7/SNvgV/Yke3+eozUha6lY8/LUbakOlKwpY0aRRO4ly
AaHbyZLO9MX7DLvmi31stT5G0VDFSIHhk8M+1GSDZF0m3Jl/DXeoQt6A1rr66yuM5aPM9Lboj1Za
1UzbCRrcvT/vyAeHs601r5ZSwQUkQSBouLLEkrbsKDH7xC4aQBL/FgpCqFA4e8FARuxqlohTarRx
qkspgRDQ5GMAgZM0Sr7+ZqCxxTzChC4ITD34mdm3YUf7IEppuSe1952THTKm+4SEVEG6NKoD2BdY
8PTOlB/eh5Sm1SYXa+/hPHMS7yC/L4FSD+heHICh/QVt2AdfoG/yscaeeGYOj9Y7Hq0XY/R3OMrc
5UD7v9hFzvglct2haYnFqBcfaFo+dBtDVmVfiq7SynsWwKDNEHuIH3AFrJUIpu2V6zFLq75D1EV6
/IBVpyOYXNEHvZ+k/SpErc7/zqmMPpfITayz2eoIy3nlv7FOWioknfMdm3/mjkZgwWce0QYSYXfK
RDwUTm8Nbmaynco6FjKcJ3n2GoHFjKORw2Rf6ez+gOlH7p0NsQ4OjasoO4uJW/TdG88L8oPAxplp
3VR70hOFKKQvETeStJlN5Y0vtZ5wGRsP9JNlS8HZZuWQ+pwZmxs73RuG3rfZ4E1jkqaTLvI8+YOu
BuCWkhWXX2ZlTvWHunD/kyCiuBiGHXMy+azBU+VeXTmOU7GnRpS+VlSRfdzbOdeq/ja/x6/s4fJf
MCFI23XU3RnGRn0bk3xriScdCVsOdkRVsMRpORfmcfUDjlNrpCFpAuT+DXTA/ZHiCLQhV2/52pj/
LAdNSCP/NVqz9JfJ+OzNqoXr7qbw6LzWJkplObuldiqwggiyLrpujF8D7P/gKUQniu9I+ZJrYvqI
K29ssPMD5gZFxRL1TDyMC5omtgudolvRMx1mS8rx81/p88RyEQHqjzrVaG6WEtT/I7Es2e2CCzZ1
UoiCzZNfhQwRavh4M/xdQwUhMoWtGPVMJEATuIqrDla+pjQ4keuRemKjFRRI6CKz2pgj31wFI1MR
0tQzMxoG6J5fAD4IKhcCB6HzF3g+ZaNXBmIwfHpbo+Bpn4tau5ZIE3QGr6c0+EKQW4vAP9ICA1aQ
h+zdHyODP5PPlRyp3bRSfiBXMGWg0tlBTTqcAWMo1lV8cTaaOaMKLK5WQHd112uQsRCa1bqDqCY0
pDJiDi6h/V2mqSpRs2NEVTukl+cGYMFPnBogfwBQm+OjQrTGVLCUdMkYi9nakjNW4k9flgUSOdO3
Y0yOGDZ1cqQd49lv4rtw8x/+UAgERnlCTXkUh5G0fzHS/Le65jjvDHUv4qM3/Zp4aHGpl1zb7Xsd
UnSx9iehQ7gonuwvI79AV4yiJaO0EClMbjBX0NYQadGp9pxgnSV9Ks4Li3IlWvxWM3THSWZZur7K
vBtTekLNuiKX+2ixYj7t3OPgINQ0YjaTXoBFyv8pnglRdkTuMP/0qbzTbzYFfaqfpFtU/RyZTSxb
vQcm7LK+NAjkAUJ2+x6yjv+cx7QOMsP7ie7PH2Qqq+uDBgrUod3ADzCsnzrdtZ4n/70t/sNVtK9L
V4KHuXyCcGAJ7PAWMACNkb0Cr0obVZ/1FXvqRRQpgWMZ+6iIC2jojXiL7upZfyoVXOhJUl56MCBy
0QT+9eol4Y6boxBWS4/E46BtO6qFLXFUNtQldnHSx/+V8WUV2l2iPM+PmHCknsx4mWeykhlscMqQ
qyizmqn3ghjjo9rjSI0fn522QXYiEKhuIDPZI41fyTs8Pb2eftn6Uz6keR4HVQkFHDPFI5t1Uc2O
xCPkAinoXNgi6QiXDnoSGIKpZpI43tkMdkgVF/laeMmwBmKnZ6XS238pW3zyvV/o/JQItqkRtaTT
Woj06yOO/f1ciazaqrak7uFQ7AQjGxLu20zPNpV0RKg7AICEp585dReIhLdK7oDxbCLuyoBw5U5U
sFBAHkWrHgCOUGlEh0n2yHqbKOl6TCrkXPfumywm/VyMERdcZcINZqBnlS0FuUNjILKZlhVKI/Wl
tDSAr9ilf+EaEhwBP5HMPLWJkNp+xSuEpwtMuj+VUXMV6eLMleEhiIKIhl81iUe/fhrAiCHXQXBB
7SXCa8dSfHR31AaJXEEukJFFwtoNpGrFX1XsVomVxz2EONYWaCclwTEY2PWdQp6CO4iHyi6B79BC
7AYrf9LPs8I20OZKQ/kHIcNO4QIHmeBzw+7pLTQkIcJIKPbNU3BRDM7a56QhiEXa9rx6oNEWgctd
15vorGJ9oeNmA2SfDAzc1BWwB/TUW6PrrP8/xFTebMJrR7jzCI6u/4UnJwt35w+WPlNgPjPvh1fF
MXBvaHuA5Xi/Pa42a//WWvaYkbbPR8GhvOEAP7mU4EzQTr++aidzTanM2dMX4IxAGtr0jNH9+tPu
HghTn0fNtbgucOnEonch+E2c1hFSjalJKPx+X+xlnsHRWG+zQVJS1yA+KzPoTxdiNlOolvGCpE5i
ci9id9MvwqpFADta25K3tR3fGcRtHVf6K8gYUGZF2io5RSwDRk+Tw8oajpaE2PSRcjSfsYiwkfDD
+sJLSDDEvzJ8sA/1u6SbjBhibnqyx3vcGsFO9lrxxabDn0Z2aKfutvf/L0ppcoNKtaoPh4YjC+fl
UZZeRrJxdwAG4L43/LU2qOb+QqW+0+kQLNmmcE1Noi3z9MPztMi349bSn4VyQXCeRrSC7/ceFDET
FtFf1qEb3vQh8sVuGY2TWMjhNGt7tQyh+E9eEHZejBtf3YaA7EPMjs0g6fdUv4iOd8d+CLYWTuP/
gnrwe/82qvNE7X5LQKtlcfwsq9qbmXK+f1QN+zwDRjCvafYYnh9WYF9qDmpqlriUjvsHhQi08yfK
+0Uno7kxozwJud9x7usMuxyWXYMoP9YMuM5786tOAQBc2iNaudlYjbtPr3AeRhOIrRm1qgbsLsg+
2tdoMU5Ot8CLzaQeqdMP2SHEvONUiMvXU3I9qjd6DpoHoj5Js662XWjJh2yKH4MnbpqApZBB7awO
X9iMqjSZInx56xnIhyTpEi4CoD73Tm7s8J8IQ4H5wCwMhub4SWETAlUot0u9qMc037xKC7KeUsDD
erDIEqVlpUAhT1iCKrwzsLeHl2QRQQlqV0d8DVEzTov0fSgIq0jqHGSYf21wctcGPNkm/qXUOprt
0NBnogzdGscT1GRcR2lrRSee1r0j9/hDQBfCmjiNLuV96mkjbOkT9HiGgpl2a4YqpB4R5DQoilwv
AskCZKd2uo0phEpHDdcuKkHikt7aZCjHkZwBEszPOCsuBqp5QkM55Rz9QZllkhEaOoPCpysg10So
twhrLTdC4Pto3YNSvBc/PqTCkMyZqKAc8LFSKn2vJlPt54ZlV4X0fe4qcv1JBUUHEYLX8Oueyrtk
l3ONTtCXMQ1LDk2uJFeWvoT/SlC6nORaGBYcg0tu2nYJU1Rg0Pq9lInFl6x1LdBsvZ/G6cIxQguW
J5xkCSoUhpLNyIqmUKRqP9ytUQ52mmDnERUxrVAzodpMC7UgGrOeVjq1lPbkGz3ZJ/aRtxI55nuz
tC0kLthXSBPJDnl5Ink1pE2TRuvimw6R4n3OMk5XAPsgFDwZpZUnqHVSp0iwfAsBnTUL4SSa96rC
axKum3rF5sMroRlavBAQeeblo0ow56W8hHrQudUl+rwW+AvjN/thO9GM3fPSYGBNEVobcMGTJ2Cn
93XUyRxJMy/7lFuSOmeYqwDdD88UAxa8F3vP3YOCBL/1xiebVAyRj7ld0ZUreXTO9i7XqpgFVxnM
vuFAmCBisgGkEpQkVMLkJDp5XCos/8Jmn0YU80ZTGT0YDvtolc8JhQRd9mskR+mvxv+44cHq8bxf
787SJZ5BAKnJU4tENbm8Q8NLmssgbE6LFyntHQYNQTkJc8zzFFSVO3q43Mv2/nB+d7JxVa9NgLgk
7vdnMDgQ5tdaed+eqdL8Yb8RWkwpHhPC/qpkWRpZ+0cKmUfVrMpUU4EP3kw591stZAX+wlQdfDup
1Qpdsf7iAXYkd11nv4xDtk1QqgGR5KNs2bKFQWeowmHEMVEer53K6C0aV3tIXNN3EcaHT5P06o0y
dXAXOBa/kLxlEcE6bvjkKrarbSyrrs9NURS0WwoyXhjx8XxuHd7d9e99nnrPrlCUvIk5B+d0zcc/
Criu9lgCWTyB0XIlV/w3+FlBsSzkDGZSdEXfW9fxHf15LEdWSP2TBGTSNaQLYo9p0TD6vB1HWp4F
X9pM8CyYmu2xwzKBkSxK7bCxSWS19oXjxXbo+TVrmxU0vMDM9SrvDrl0JX8uHAIPYbOEJumDERxn
h5SkCM42h5oOa18qJlfAc/QQikwEqr19btf/J9GfEcje62gs1tr0o76UWY80mq5CN541HVGcFvjG
mOQG7Dwq6Xp1nnqGrxOGHv/xFgUPCJ9NCKwFSk1s7UpW4MTY7QtY41oUTzmt8G6WxcauhZLq5/go
WZVLNH1buN0/zWNrdhA+f+MsDjzc5hwG03ioUYqVPgb2/M5+nviV7tV4utGAmfldeKHr6EL4HYaD
R6W2h/WtV3aAGez4Qv/3/xIdx8WpEIUZN/Ti23Rc+IduLYoQv5DYhgPMY5qPr9G9MPeKzcpf4uv8
9GE5GfCpaspMykdAZClaYiOgom01X1Ktq80zuNuDJKbAwI865lwNc3EAkdVac2AKueEFrKMYMILi
F7zhIfbv0AZfe7tkSGQGvPj7/Q4hGnQI5OkuIUKumOr+THtlTySZ8JfXa5RvfULtlpCHyR8y68ox
S1AgyBYSpxMaZJSVW79pOMOvJ7hQWn8q25OVPzvpYpCNhev8gQD1huqODGFG4IFyoWch96iYZgEn
9npl9+QiVWflrvovxD2gMxK/DH5b+dMzJfxIh9SEAtCCbZqt+L5f8DMrcs9GP+/yy7IxsUmBa2t8
ARyDpqb9bdcW4LfEMDrxvGWTtqnyvoqHOl9uU4P3plo8PZU/M2bthPAXtxqa7IRsjz6SH0RDQxLR
mDol0l0hpzh1Yfh2uWxaPArDaRvUj+iySG7I0oTPITpXrp7dU5wiQlX6vfJzIPk2Kx7garkWB/Sa
JDzrfXav8L2TcztnrH0ak5oX5DI/FQREeozQOBGo/eislWsB4hbtMeqRjn8L3KWOY93hX0KJQaGR
g+uMo92fXaO5zcskWLmES+YPCM29jEvW8BIqPnyyyoM5cL/QG+31KiMPxkaeOOVQEd+g7WLvEIYy
kedDco1dh3v+BDNsLkpJnX48HlqjIZOU5m6lmtpNZRrmYV6+ypf+pOe4wGyJExnoN8ojIlf+B0Qb
PVAmyafbhXOsMQxsDsF0B2AuiBtXTz9rnv3MfJEgVJ4dvgd3l4hsWd8UDgySKwZ1kr/9cpSGt/N6
1THWddwT97POlRwcQRCrXt8e35dBO3t/yUH69S9Gz4aTuP/PvmdWhg79JSAYf18Ax3z9uHsguZoH
jYBZsm3np5pP74/BpRPJcQMNEr/Wy63h12U8iE9RZ9Kt/UmJJ0cAfOGRUI2jJyQMIPgcASrv64Bl
FEhQbjgSjGYQQWsliRdkN1c6Lr0e/XSdCD4yfLXYFn3whjjJiUUEjwznebAMo4kNUC5XFyK8J8H4
k1tFKtsmmLPvhSMkZBkSzbWlakCzkuQb1UUztsrCwfPIBOI/6GHRG6DV3hkHvK+nP8wTNsJwqYpw
lqWH/QEAd7GWJjco24ms7BmwAQtn/Zx7FGnzM+RkyRR5f4UhqQNvEf4noqI22Vn9Hq8k9I1SyQPC
/gBPndcOHjMuq/chxfGeQi4NIWbrlKtZMmpNEd57mJ6FenKaF0FY1By2iuAiJhqAiU/iFvbGKjPH
IbofTcdUBce6FmS9NN+6Kv7Vm1UyqWw3tf8Q7f9ofKmPhujd1yjmve4LtpOh7ZE7gBN91m4ySYbI
Xo3bIZzc/aJZPqHZTeS9gwnUR2T52ui4BpsXuRdDnYWmYSehSA9qWXoRzIVhKt9+TOFihITGcbCi
5JMY8UYfHEFJEAG76hmulk2Xe1YOuBjimZyUhVWM+lX2JJ81gTbfxrPgkHDucqzOqDGkvuJDfEvQ
7kN3gdGa8BgWs0V+ZIA1NPx5700R5QFQi+5ZUbHL5iGYeXFVybL2h1qL1w1E5xQlsNv3+YPzWp1u
KWQSqAHyBzZNTXIu+oIy+LjQJZ2CfBU82JyzVXzATEbjXvhAmVAopw1hbks0L7mHtZp8Hwag3eOe
JX3ak/FeQgOPkomatdZqYuIIzOjUDgQRw079bEewvsoaJzqJjbhP1fnWcGtuz542Km+Pj8MlOnLA
kgfyOPCOBRulFM5JFi8RFntRLCpQBs13nBBhNAkF+M+wuR1++6Vq8NsC4NAeGq+PMm/VM0md1s8G
tMmx5oLf2gsu89oRZcfGvubSxZ7cxKoC/Rvu+qxxvi8eavuHEECTHwmfo/tBDCG+6k83MpE6gAPK
18FB3+4VMDKlXm+F134JeygkHQdyNNRtHRC524riGPm42YIb9wKqcaj43Hys9PMGfkCIaGZVLlMQ
YUlcou7nYX/myBJyf5/yQ2fW6kOvaxZGXOkRycJhWn0EVklvlvdbCjXFBf6r2EBad+W4rRmfg4qi
OK9Le52SgJlMPPcXOnCDHeecdiX5/18oQnyZlClrI7GD1rRO3OA52RBxV3nyEMaKtoGzxGFETYhs
jn1wvmnAPQaYtdXn1WgJWn6eKJYAvpfO/6O3wJTORB/SvB1VPGSR9Q3HRXOOAN54GO314ttF0sHH
PISpp9R12Rx5wBNWFLFtqMsW/hBjFjNfjxK0DMmwqbT6wdN/GdGeisO4FY4ZZvVH6I4CHrb+AS3T
qv9Gk7jvJBZe2w8KgitbuYh59aEq77f8i/ucMXkqkHeL4AxknLxWU7jtpje3k985BrxwY1jQo+G8
/lyQI3XhNet9Fiww+hH/81V2Ipcbiz1GQh/byCgeCdaAQNLUFnLKqi4uh1dYWhSDUMxu5drU7OnA
OkGoJNZoWpN58AplpmJTnGYrOORK/9ILWCmv4LJOYB9jCQLIMExWAfRVJevibcnWMrPli4udHiz5
+ZLvpMNIuenPYCwOsTpnBkSVOEmChxO2rKdi+ZIagty7Vrhfrvgrf1x3kJs6YuwRQjjtwa0qEZE5
e2E0bRywyW7BA1yPMemaaFCOZFN1N6RK2xonMOEeFRyeQgGafv7BTefpjRmeJQ0SwJYSf1t5AxgJ
2P0RC4d+pXQ0sXiuV4Q0yOIyEmv44UILYj1MqItw5SwilFB5rj6jHpyyujbrTLAAu4RSvtlbeeUd
1gqPOf1CXGUFNfMjjggpf4apjebUze3t3iO9dm2rtJSDA/ByM5VsCPk/g8Fa19XvaN0S5TJ3dLnf
7mVJew+GJl4HJMNrzUh3WITh9D3TH+nUTp8dh0l8m37GURhoIq689s8MX3iRuE6jrLAArUKs24ot
D8ffMbS7hoIy1XQcHSKk7UrdPxzSneo3B2LbJmmam8WRo9FlxmXCh10BmfSGqnlHzYJCkqH3VV8D
WjrwbGA5BVzOKXu4OXNX+/gYebW3F608nKOwPTPIm/7OiC3O5xQjTg8VWiUEOgFSRp5mv29SacOL
UlYqFit8RgRLpyhUvy7iXLSqrCgATd8cmqMaXowHnG3nMvdQeVZ7Duuuq2mCdblUUja6EJ2a/hKK
3QuNfGVFl9q71kJykMUlV53S+Es27zGuA+wDzdzNobKREhIlaV/rZBzP+mZb67isscjCoTxYZ5EX
fvOJs9dnvL1yOtoWBWQFgBT+ycuSfuvSsUTBUacPtTK/wILxOTSbRh/iZN544hBtyH9HG4LpqZJG
1ULwmpiz8vkooDZxrNcNErOozTCjIeGFIa/qthBWcAVlOXrwuSSd5qhI2QEgzoiAc9+H1AnJjuyM
ZUsUc6VyHwrCPKsq6GQYV61ufar56l8sXhMfVx0l5PgZT8WNPdNCPxybMm6jxqwxzfZPWyeD2zoY
own4AKIIZwpLeZJZIm0lti/OYBqUItqdiNDIDTg7jCpXJrXKBirRE5WjBUftJpx8B23+xOnHKWPZ
nr2SOtD0aRyfxFsh78YnA8p//zfJzevaRokD+SLZ4uvFkQJ0SIGw/DIa3hoD+taZYbilKlWr2HHY
O+0hqSZCtgiQAFEaDUUHEWLStpVBxed17oY6XBBZyvM26wdnb19fggZWHQneSRBgw0NwemRgWfaL
xNT+L2fgho0otPGorS4W03T+dbRM/u2wQ4RnAwUEgwsEjnSrNW4ZJ+3u9B77lJJt/ciJSOAz/R2s
wffICsDlKOIfdPk3TNdOm6fTHzJgSTCFCvTE9yMujI9+f/IHkuH9zkF8QisxrJEU9By27wq0t5K4
iPFV5fFqs34LG6xlMbVKILCALGL6ZOEBwO7occOxgBfHtetspaicXeZqcOG4P7o7tSgVvRCFlEdK
ZpPJcRyM3Xh1/6GrHNSEDb+wBrnqn50rtdpSzyL9Gfzb1GjL/c+/TSJZ8keZeCCJeXPR1KUc++/T
8v59QzWrJU+AtMaD4p2LXBPHrI5QEAF3GbSXNyQA284ER3rGfPfNnLlkzfTBJ+E/hLOELlykgOEc
d1vARJt8AililzUOeR+pYPFZxmBZWjLH8Z/WGWRGQoPEvHZKj0ugpxxvtWdXXTkiRbTWXPcXHkmL
QqmddjKg9meylj+AkTnYMECQOIL+to6jU6yNdBnfx7FxMpGHv6LN/1RyuhrwjhnjSahbPS4cOras
rRfArxukxTqh7XIJPAWyTw+U2CJm+zJXV5JcIcg5uQD20YU/I9fzjMmjYHlHU59aCr2bEENy5lGm
WQELA1+a8BtKVMFiHS1CI3iimg1iGhINU5L97toAGtuYuvrlxZ4bB8kDhamfokOoHGUmV9+vCmnQ
PRQgLU1LBqdaP4GkgGzgKGnh/9Qa8WTXHV6YuE7eUQSPLxZ8akWhV5UcmzK73MrkQZ4Sj7prmvhl
SNy4cF6FwmZWlQIMgpaZli1rBoRAlNtBF1F0ujyFeNAmkVWjjFdJ94uXGcPp40TegJfgqxiN7RPU
HP1IN6mqblyMI/x9G+JLmAXIr7x59O49HIrJSHu2CxRdgEmYgegvT8N9JLn8S2/mJl/d9vruD/3V
7nYhcnFTr/0m4Cj4ep/WMGJnskeYmSRIk2W09O7ljY2kYuWVj07T2HBELR041zeJ5N/7JcurHfXf
dRieGEheP6zzhzvUsIvfVBmyWzLWqF9SETlNoJ9+Dz9dBtBDCf+bAflUZK5ROnfCfYWThRPg4ry3
GXlHPl+x8aQu44EfEyX0+uXsrj/J3Byt3bR1DOlOMyq35NWACHN7jSXtXkFfd9e94P+2DpWoZRD6
YwoElOYHJBlE4EUbo6OjlsTvvpGlX7FwnsUzc4/orLIt2ZIbLWi69bQGh4M1bfelK+jXibOOQpak
J3hndVcEJ6o1CLjSpT/HeDVWwjKosAHhzL86KVKEQtAQkuRPIqz/kxsd6N7mtQ3ZKtTwLU2MTsQo
Q+c/pTc4pawdEqPmV0eozWZfmQ6je+xx1YigJvvOBJIWDSNzlW9RD1t1jOSkv4/5O5Xbm+zaQ/fC
yoEpAZGLME8AWCiUPcjUCF7QvhHofL351VlPEh9Sb+o1vby3FNt0tdGwb5A7Ha4GFoePUJfiysDA
x0WtPtwAV7sOPYQ4QpBvMSyUFIUwbQW1flJW2QFKI+nHnxGhB798Ba+yL8qn7WIrPwrNiqzAAtwb
cKjG5lRsKllBHH+5ndSEPb+eAqKL7+iQwE0SAcP7KNZBxqNDh5WMA4Dtp0MMsEZBUFRh/yOnqYfg
XK4kuIf0cUqUpQkqv93vL0H5b0kaIw/NdP5In6F4cr/6ybaSLsJqQvYAHm0TGtYMjX2qbL790Ixk
kEuUlOIsDgInNLUmYl9waJaQRCMDKZ7m2MTNR7GCgcFZD+Y4OYOQ5v9KNX/aSTDY9m+jNq64HkvV
lqtQ0G4rRkiCajZ3MWJYtumJGrgzGvBRIlfYyK6UqYIyjV+JDuMMEzEqy77zoXNBO2t/aCQ3YOHi
HGyNJsV5PND104y4GIVcJXNdqqdDQQ98p1Uzaf5OJtSQVy+Trd9jGWXrhS+Z5Q3hDsuy0HAIOldh
UMZmftnlnoL4uwTZqZ0yZw4Pti60h/JqULdzGZH4WwNqrDL8SQtLirwKlfWaEdpceuxX2bacVmX+
45ltakPkVHePhgG7K+FN7bLX5h9AtldtCuPHt/jWxHc7dp98hvZ+eehv+BUUSZmALUep+LMy+zQX
SmCrqQaiDR39XfyyJxZG0vh8SFf0chzPtGx/k/rLl480E4/RQmiLpiJrrxIhC2MVAzUSud2iMjDR
2+9H8ofXgCdY2Og1pn2OuAQVZ/VyLjKz8XXbBFcqrreQdgnzXWVubLihaWz46FzMceIlf7ixf/Ku
vj+O2Zo7brmTfptq7W7MLfxp2gLKKkylVuJLpLnAtOgKCl+EmqVgRpkhT3hwCqZQWwASukr/B0jU
jV2fLQwjHZrRf1vWQWYXYUwnJN6EPKmPhybg/93KyNiNZZJ2vZsWEd0g0wECBTfbtv8k/BcBp1IY
ofPEuaUVWdwjy7RkeBUAjPq6sDA5YKX123lHX7LytB6lPxkRqs8wxr5qX9YIMvsFkxI4Cp+ywuFX
nhDJ3c1VYnHwZMG7wJjB0tOTdeUznAvPH4SxuPo7qmvBr+MUCTjYAC15e1WjpRDqJG++YC5+whAT
r4hMQXJnOAGUobSu7SLLk9bSOjvNCTfE1eD4HEk80B0BXeJZYDuLgNuSPGqHQLMahA0Yl4AXjzR5
xNUiQZCQ2KZRtUrNzAz572exzCT7Ks/BbfGYTFVXGJGeYJcJ8z8Y37naHZKFu9cLfECAqHodbVG8
80a8DEoAGx32gnrNI50erqURuBVBVb0rBjjSGc23FnmvJ3IYyYKZfP5lQiAxlMRBqTUP+zJSbzAX
VfvquyenHdM/UCmHPmc7Qma1pEGvtNueU2GZZSVSpIdMfYaHpFfTxIm375AsljD/qZZxxKjgOr1O
DuIdNCf/5WwbWiuxR5T+57DLbJg4tCHJ6WbWqRh/utOdXqBPETVJlx4o+xdqYxDb+0bc+v1DOVbn
c1kJTV3xj18C9UlZiBICtPxLE0kGSPe2sUyHgkB7pfEHEsgiShHQ4B+25Q6lGk6zABVaH6eLoWZA
nofJW1TcyQVw31bfZW/1OAqAYP/yup+q9OsjR8Jbeo6Oil5MYIXWD6lVJWULFPuHYIkw2vABXJZG
LlvtWg3yw0qWA+4sBTWAcnXvP6D5o+bI7Ya95T/T4UUSAAbDiJcD8yIcQVjf5fOeqD8F6tidbGOd
br8fWFV3w4Zx5DS6g2arET69gjtth3xxIVX+rdBefz8MAUQ+7Rj3e6E8hqRvXcRlIz9nM9hmNyeD
MLVlq41ztjczNdf+Q1W+0JyMKuY7OGfrKhckdYTk2PTqeiecftYQyP8draDd6xxI0x5mLIBvvVVt
GUnnxsRW9jTng6NxjXpNSRYPmTaCm4yHWKvgLJyJ+te+PIdSIbP9QWxFzxopgx/szRCauJILzVD0
nZhoWdcIUnhlkeG+WVlF3O/qMC4A/ep8pyIes9kjZmX5kk5FfYwALh7w2cDW+aQvVBtapaGUlJ1D
ZwWYSDVu9AfkRsiIlxR/69ADfmd+NYp7/j+GCY5wcOhH3u/6l0VHHv577OkTPLxf+NwX1wbhIh4c
KnoyKqVwsRjSzNZa87BnucZ9pNMEZ4Nrl21NNqvTh/QDkhpVKe5XYh7aLP16mvGuQpvxthOXUtoG
eyBQU4p5bPP+NrQQLPUW7gV1xYiZd/ZjMgrouFDA3Vc80SX2Hg0fbm53meGqdM5i/rJdjKQOVnCO
AXLWEsaGkBEQSkOktbaaTL9yH0ywHIS5xSeHUfS8YePp47gjNNKR+sL6gxUBlAmiTVoo5CO0I8RX
nykiv51btULBh7UlR9/ycdrP1NepW8/GXVBCr8Z3ry0HRAToZrGNFmLSAVQbl2+dDfJtoUpoUUpV
PhR1opHXA+czBveH+I8/ZcxaouViZOYSivfYgC+d3tpUeRG+eMQ35k0lPiyS0ACwleF56Y/R7UEl
fohiq4WJ2IG0A29YksT4FKGiPIg8H8++tELHkqFu3fm52i747Uv3TGz3kz92Tfn4AyRmhjTRQxQ2
b6N+f5/aMSpu2AFSk4xGvknRGJv8bNO0b8VlYcUat2qlZ1dy+iGbw/PMoM+gPnDEiXBFwYpwpesl
RVjeM4ws+5ZZXIf/Z6u+lfB98k7TvnWNF5Q6D43Ua29eQAwL2l0jKHiu/hAoel5qZpuxd/g8AWGh
eX36F2yUN3Y/NCL58/tlrX1Ja5jdonVKLbKSpMKxifRejTGpGw6BdRM4WAJuUdlruR4L87kvAh4J
gzj6FgDQKwzzUnHeuiTZexRXl5TUkcW2ttuWA95xVm/rn/BEda199ZUlkDdRtiOUXBZBsb4jUS1g
yGCJEcdOChclOZqS0D6Hrc4lfmzz0Vag1+/7cVtlVGHCX1vVTL3uvt21jcRpL+jL817fkx1K7M3v
zQ6ZJQbAndiAxNQYC7d3w/vJvyX6kHqHGqtKejJIOpqGU6Y/9WX1WUhFkskaoemUghLvk6E1L7FV
ZvU5Gnty/WAOKAiyRga0nAXhYJw+mU1UBzzbXB555mFSs9F897aMM6SCwh0apXzkTK2MwCH26Qv+
y6zLIFnWfPzzz8eRlD1WZ+7hNPHyrnyZSnaR4xyEbDZjD4BVukCfFMomq9gn+UGBJOmZK/sj0V78
ll4WRSoq4NaACGinwF9CvbfGLg8zZSCQBpxkPRH1AknpAaEviIgdC4nbbK+iL4C0rinmcwjw2viR
edTHEQjiD7XzE/GJ+md7sAOOpDzv56Hznk564wCkVWlYP8WvvOtUSbLFIDE+BaBGpO2MrWQuMqNC
RuSCogt9DXdAMyhTVt7EsKAPxol/NgzBgNa+GCCQ/M44fv+3ix6FyXrcYvFbzi+9QuQK3Ev8/RsL
DJ/9PHvJPn+7mum47Md2hHz2PaXWCa3gocd2sakU7VTwQ6hix/KokGdHG8lDg8XL+CZ5LlqBAfsK
mwZ+01Z8dl0KHkJjmiGF9OcMGnlHLbZyl843DI6My4gkZQiL6NSeuw9nsS0uRtA9lFKgOTw5wODu
yzvTRdHHFLJaEaCaYssxXNhXaL8J3zc4oLemR0nWP77NFSnYq9fYzsytC/u949m7MSUO37uoQ17i
7NkGN+55Iaa608jknOPreSfFafWVneyaD0uSye/V1UonaomV3R+b/7sPc9gWkJ+7tu4ee97XkrCf
vwLRl6MPJ1dt6ds8vFo+l9S4xk/FoBJtPUH5bNzy3Wdo+2QCYAYII/5vEvZcyZVjqqztH2C3mvTG
yxHVuC1RI/0PZLaQ6Z1e9psOC0KE/xXH+fWr5AWNSi2llxr8ts0MasWRXgmFguDP6GuhLFAEzhQk
0TffSLrlK9dj8ck+FjhkGvIbS4ejR/Cm8/ju2wPYhaYFJVjJvpccqHw1jvGv5667uQmFe/AKTKJT
inuewsXK6nUPmtC9HCvwjPG8DN2ngGyhe4HpEUIlzZGhw+L4ag8RgL1WadpysyeRUK4+bgFRp6uH
jrTpr/JzHLgPwj+WHBDgaMpQpkD/SLHX9m7/5PdF1eRerjvzSB6S+RQpO7wMwtC1Ah/bx9JWN83v
C4xZB7xs+LBmFh2K7IWXfZdVU68uVjVMcafyn3qjxhEwBlRARDvdvJoxO+xD3PJrfyF3dr9uQDeq
Ubyfms8X8Pf4TOuVwM406gKBGGSxFzKBq7J2ht0NW5Si7kovWwn5xQfM0q5Zfaos2cGV+ttThRDs
+0pjJrGE5+rRCr0TUl0Cpg/9y6JFVmt9rqMfMfr/61edTYXVQO2UvUibBAJuQY5UsJHu/wn2IaBV
C6JZ0DvxFohbAK+hkP7lHcEsfK9jbadJXUMc7Xnas3zxetU02aSnZffE4hQw+WrBi52VVfuAD29x
kWzFcVW095TW01h7crJJnUunpfeB2C3rpNVYgAP9TOi7U4hgknezSzDNGRpwkTM2SFe60a/5DIMv
uuy2A2U8d67MY/tZjnC/NhM+2/wMz43nac3FI7gdTNtPLPqmvwrd9erIKeozHtoUyGlTLO5REeKd
v2V67UH4r1tU6VsZXxvNVnt4fCKW8M2KH3MtB+s/U1kTGuTIJWHjfUNHVMVDW4RBO8N92b/36HWe
xAZecu1j9dtJxnXgHpr+rnWdEjwHaBrB+h3HMU6uw3cgwtXV2DnLyfjDfDA8ZyfV9SM5buyg4M4G
e8tbDQr6CNxWfnvnaJVGx07vxwZuIvtZvpu3Kynl3I/PTCgmGy5cAU4HiPmExT3wepc8ul5NwwB8
Tmp1AtSN0vRL6iisNm9FQQ05h9nIvpsB1I67qMHXZ4EvZnaisdjlcThabFVBn0SR0y2LmMIBn/bY
Txmr9uz+DEoX3yDs0NSgmMaulqJPdpJx11Lz++2vAI5SpufT0g7tmOqryDUarA0bND8D2XRZ444y
+jecHt6n0sFtdG27WCVJh/uwYYrMZwcxIQ2CdSefEO3ZMh0huf60zEiTArLoZJ0mlgO88LQUaa8y
DSKpaywrDcVFyzTThR0HOK0ye6xFgLfIZ8RsC7BeNAaWcxdxWtqGfUkXX/UFp5EP/eXr8YdoUi5w
B65nmUDXGY/4S+d1J/kPBXdivQ792DKlyMed0+6kdYNct21Zs++ZlMKiHsoDnQAcCG6gdzRsz6g7
5eSyui+N0ZyakU9lU0D7S363R0/Z0rqGeIzclMoh9dbkXTJwcfuq/qj8j2aAIvit3veSKQYwhSOZ
6ItUZvXd3o0UNIPRRCtXsOtxoQ29tWQMggnAtpCgSpdW8xQXpBfC2qtjTBAGgA97H39vh5HpopgK
UDaqhUgcSenhpnVriyyUOAYgd1YRCYMFlZOlP/lzxcOcQ/nD10Pa9VKefnuI8l2LaB5NnktTmHho
fzp530Yp6rQyEYbwV6h8D+E6LwL5TgYM5ZkcfKqdrfcLj7GcPyuUrm5yu86bTosne8eG+z+fiwwG
zu4n5cJaLnIDcQaH1r9ZGyLnSOjqOrPH3+AfbJeZv37zEcYUnBV2lyCsRsK9KIheujGHkOxeUxGg
nfDvsjzCpX/rZU6D6J9KXM1AJMEdaSEe02/OxoHODHgCDiAZ0cNJYnECDYFVrN6rp0d2vldP2Qgx
3rEyWvQ1cdJKTFhX6odpTvbcL87931sN3GMGceI79nyyJJAPEHjK8A8fzOZlp1XHZzEuQm6HNAGy
ym6fd9120O84K4olVWt7bWa+WHjiLx8gkNv5hzCyyRbE1ShVdC8VWwRBDYTcibG9jUsiSB30u2WO
yr3YhAC/99oVqxcq4wpehz2Of1KIlHUv9C9Kv/dpmTgQv27lhBNqTvFB/gVRSK2F+Aji684zvf55
7QoPcA4e0sNz2xm/tNRO7XaYYVwiacBTT3tLhcCMJk8i746wuk8CDyInlzUKsS3fmNHlikBjz2W/
Lhspa0M0ZDyz6xzGklA5ruR/3WFvtvbpg/WiDDVkkj/mJ1hanu+UMipe70ehqwYUI79cGsAU13T/
j3k2LoprPnvII/AozJM/7EsQuRdnq5mV9qVX2R1VrEnl07pqnBR+EtrYVGBEVXa2mdGRJUKEF63I
XoAGLBbu1IKZhhA4sV71HHsTvfn0Xlwu2SAr8jynXCXcyou5ibtLPvb/S356z/yaUXr8WPfc9pF6
Cudt1gzafX6n0m51Sv3DcWkSJdojr7nLAWV/Z9ltbuM9YBAOz7O5TFWNK8LTOh4suaiUMBHGt2r3
VPp0T87X3AeT5/vV0rFHvvhhm+ZZq9npMd5s8Q10pf9e7H7T4kIF6uSpd1R0HheC7os6HXZmDg+G
NN3jn0hNTyn+3qJetgRAaQQ0XaoXEXaWXavsRQhHey0I2hQ9ykPinYSk7Tiyrphd6tJr/wW00beg
ZswCdqavOFogaF7ylxQ+aC9ARGw8snmUkOiiXIqlzNwupwHW3iuKXAdrYMrnF8flwbZ2+hmCWMaf
9uX6+XioenlXve8IuL2+eDagrlfiQI/5mSkMtNEw+/QCX5ATXZ3GovozXNWGlJjnuMyEjT+f8yxP
d+aaAIf8D1F5YLXaZly3g37fY248NUUpLAoT4K69bYfPNWDuNFLQRYMg7Wm7AIEnFAa5E3Zivzhm
wI/qWjTVrIAA7eNcfpm4LecBhtzKv3D5hHOt2HVsUpYIcHyEIB9bxDK4rG5oCc60jHDuFOS1nqaw
DXdag6/uuAN2yDLuH3LAjgp1wPMSJzrwW0d3tNgjhu4OvcQLlXRBHVKdhc04xHsPJqLBCNviIcqo
C19nyjS12vIfwdyd20O/ztn0f5+FW8yHoLWRe2bV6xF3qyXBsdTenQAFz3nchgQzsBv1wJwH31lP
kdisLWKPfXdMu80M8XJWm2WZ3VaJhnYDI9d70tKHECKys70UjAIZi8qaR91BQd1sbKCiNjPGwJox
1LCmmeJswaCYvu3f4buZBx39tZDYqY/4H2HcYR152wpYpBD5u+j1OMZNc9m+iuPUCyoklbycq3BY
xeGMJ7qDB8LXRXIGuhznsY/7ZjmUMZO6d4uPQBmegZTit7ZqrCvmecF0JJnG5d2rUgz3wgb6cmtQ
PNn+3YQo8svLyWR+UTz9AfTxwP7A0yK21KKSqJivrTKAIofIHQ3kM4OROLYkZ+oDq7XGIGjko7Ry
SpSGLSsjPjOBst/Zf16/VQtk58DW71bfP0M+cTvHV5jzVIqvP2+21D3HRDuPn5Qa4tlYqWaszGd6
/Iq457BC8SGlvubO0pGj5jk6FHTBfuIBkfd1d5Vi+qSQOPaG8DROwudjifL5QnyU5R/Egk+qg8bc
NgrCgv6ZQaby9jMUoQ9VUI0M8rCkjcdPC5qKELKQxNZRGC6mXse1FeywLa8gTpmQqM8OhBi5lFSb
QL6NrllQotbxxNQ88b+awLHdNkRIPzVhMIGG9BXy3iJVOc5H9UhN+jnRiBEWBCuuexXuSMdhpKEE
iCYp5RiYzdYmqhACXP3hgE2MyR8KTwDwGbZM6zn1yLQsi2TJrJSGeMHDoGgU59hM4J/UWZ/H6c34
l/5ZPOHABzm18uaoxzBqgxlsi2V9IX2rKEMrBA3MBgTd0V5Upmjn0pbf8f+xxAZoxwinEgO5Sx06
6O6iP7HvBXOl5+HdCL8S8wJNIc9CV9KIiOtYeY+gTPjDcmFkwHNStLXbXcLxWEY4zL2sZt1B5al1
UQ04sXDdVNBeEsy5TO/fKTBada7v1c/+cUbifv1EXoFPA45F1H8WmxLXSqDUO7Ccn37Kna4i1vA5
C+tPhk3b1jo3hL02GgFyoE53fy+T6YAsJEvSgucWc1aoY7X33A8ug4co+ShilEA4OTSAWmoMqxHE
anN2oDiy0O0KoPRfyx8ndTVtfCpWkEKlqVk4bKUsHCDW3TnPanRD6WNk/bZJRYjjI1730V0aUbbz
NvlgHeDXjZZWKuGlRjC2St7f0ZOR9j8uvTKC/3jHbmPBqdmTORLVpraKj+cZOVTxv6RHbGqar9jg
ZK/JNMCbtUPXhw0MU8nClW/hBnvjcxXnt1OcdOVsRDzfhD9aRp/EM9UUHqyAGzPBlsaPV2obC6DZ
9Z6JoxnElaMh2iOLAHF8qJzt5z6Q+bzJiAigpSiggYPnpheORKeRHMtsJO+p69CBS5c+neh8pIkD
jvJZ75FV7x8qcSFJ9R+VtfXGj/QQ3CrbHZKJfjKnEtYBBWU3WH+CabbCKeXBN2ZbsWI9w7ZEkdFg
5EYzSHiTo9Csl8/j2Qy0rqmCNANzbWf68PSkkuOvGBxm4ok8y4MVneILWS3OktJkCUHmfbhsWQuC
xudF+rz3QUzUq+U5HupV/GlPeddFlKnZAqWdYMpIkMXEvpofJE/mn10pFrzzgsAu6Q7Zb5enQ3S2
dYa/xVw8Xarq5KMIeeVntKkjqk3rlF2kbjwlXwvLRcpPMtIz2h4FKHKgBzRedSyLuqigDElqG5SK
ull0wqHzi1rCWVVmCkQlDLOvMf8UGZ/ZPHpup4tiltyvKmV54ouAjIx5s+iYDTWSz4fJjE0zpxlm
0p+4CILN1awn29BRnWRwTjcXlGU4/jpON4xwG541E0Q6haprys9E1u7yXIwTgiZffqlwVkCaJzpG
IzpytNOWsi+8tyACFpQ+y3Z3Hporco+NghrqwC9nRPzvyl7qoDtiYkeVnzaTw++ZX/oRTdmpqNNM
lWLDr50iPcIMp+LPWup2Hua11N7fC7VnGrO7EOl787dpk5yyomdN7HkhvWwai+DX0MYNS8nybtiM
kJZDj8fw8EjuCtL63vRLKHateMc7S6y2t4ff+HmanI2wQhYJgONyZU2v0FinE4ZHfsNLIKDP0atK
NX/PhrlOoxyiOcAciHzvcMaHp9wgVDfoBxsvjjVnFIzfsuDNYT1ppJH7hIRcCveWWFOXU/I/rWxD
/uEttoIBsgqZTt/79TSx0JaEfY7EBYK4NP7G6z6E4BDLTekb/1bQIKg6R1yKhI3IvGKFasCPvN+O
bbb8OUrjL2i77mY+8zpicQhT7EGH1l3PH2q3gul9ejwOSsgll1ziOfSrHCcFM5ah7naOolFHmgjN
VYGlWDJtZtWTpv0sBaCFDCdkpEUK1Ly5Sa9Fof2pAzttg9ZdXUTNBA4YU+W9pVYZBgDv4OQ5t9Tt
uZ7hKE6oOaqlgurHxrdhUVSOaHTwWb2lJPzf0Uo7maYE9ytnn3W712vS+Fb+znay/mFAMmsUPOOz
L7FUAzOf67gU51hx5MqrPoDTlux38kBR4BXT1/iOONTjah7G3YRpejEJysO7ch9GEOz4rjddNI9Y
1X3kWWKJEoaqYnWjlIRMyB6NsRhOoZsJqiY89G2W8eT+a+uiq4WrodT0M906Ixcu6seMu5pE+SM6
ZdliHfEUOcWqkzqbNojt4b8pTjPBd0a/d8lOozfjKolbwrp9v9UUY0i+PyZEGUXB73kYObXYDvDd
5XuSvGZFTKXvfS67qnu7B8BLaZ4NuN4+niBSN2EHlz/JgyyDYtflnFASfvbzl7LcxLB4+/Rfqtg2
qWKsCRqTxNJHYGD4mvQpuT4VmWALul7/CDX3M50MSqQUQ6W3lLYkaTerJCsK3E48KciFgxJx1P9w
5vfxIXiZlSQw9o45O9zL9FsqyoI9NjLY60VJ3gzxFLFQT8qPJ26wFMfTMg6kpE4XdbU8I/y6n3lU
MPp4QMDzRlzsZCkqZtc9LaqfSA/VYHZIzeLSPeKp56PA9P+0PRcQ45mtNwtiw7jYXOzKRt8pIxNH
XdvhBKKtGys3s/QkqKjNdJ5uap+zzkzvJJsGjCXXc1ytZIk10BJ/dLDRQPf2sr7C22N7bGtbAXgv
HxPFqGkhcc+4M0S/+Sf3zxkqGXrpGmpDaOEjxtACEl9hYkQIJiTBLZmMOK3sQkXV2YKa0DqtCUR/
of2GtI/X8HCjb2XZzOycDdWZ0EmmLSjKhioIEkTqH4duZOYiCXg3lNqAlzwgnJ+eZG309kw1/qRC
CJlDVVMVyTXuSZJQPYPCVbNMqwrGFjpgvDPmlUAmGy2br0OsEbIt4KhoB/ve7gRAB1X+QJBz44LO
dxIC+Lu0S/ZEzSNU/uz/YvsrtBK1oiAqyRD46gqHm6nk5ftM4u3KdxkMkjwaUg2RiEP1tIhwwhqp
G7xY0X6DjZxCFmVbGtXVBkrYVaPNRnDsnC/1lFSbx+AO9BGxx5RVKQOYaRpsCXU3IzAv8EyPmoh3
XoXZiuSqLQfFGhN3GAURItii9nRR9ltNBrcNpbEOWCCXxN8rTvhYFZfG50J8Oex2+mFY3AiUSonU
zZjIABCwDZ9sB4Lk0CobgEZ+uz4dwqAa4j+JzetH7A1OGhaUnKBmtyoeBsDrN3zKgCC/B9IF7Iqm
a1Voju9PKlM0ua0Avjx0fbTeCLiXoJiZQgGlVH9U9iWb9HjrgYl6UqSvkOkNtbxv5LXBKWvuHXIn
gnZwds6GSI56V/6jyEliOnHCJsU96WeytNjoC7INLNf/gXDjL5ovoiqu4O2HU6rl/7Ek4d467C1f
hXnq0loXLAX7O0RqH8/vlMsMuaI4/sAvqcCxz5qcl6dhxJ7exQ4sTB0jFAlbJSFqcH4cMTvwC0d7
DMN02HnBp6u0BNDGfXfGLMqT+UT1U61n18yxYdND8+dndfk40ANZc5/fHph2i3jS/djK42elS06Y
nmzm9bhjX8kWQQ0Hh4j4WtqxNKaynh8OsgnkDimwb/LMbvjkUWW/+eJy7fq8DFIgird2J5yEiNXD
7jzzenGxKFff1TYTDPEgQWabrXOJrIAI0fc42TCZfyEbAsup9U2IH+IVft6DoLaO28U5BwA8F/Ah
jVdjGfb8xr4m+TG9lvHAPirHC3ukhgp3grOxaVfMDr2MidFxFxZiXSRvqA7iXPcbrNKoTacVPR5W
ryN1nTRFB/OTxi6JRmvk4y7Yy8AQe4ONziZRalsLhc7To0rn9JmP2DHWNghSGnb9LQ7I4/6Cs9lF
DnkVY4jS+9wTDDQzQc4SRMhq52PFM2tdssOMZS+YBPt34qovWzhu2MUNv/loj2My7O50JeIEJ4nc
+3qPwSxPJLHdqhi4d2h4J2W4t9TvUij6K13vwoe62n2+mjVJIJGIZ4IIT7yuVpk2y4MAkOQLMAox
7UXZclp0qtEWlAJ4OlXVPI6ZYGyWbamckTPPa6DlpTXS4bElCFqlJ5QqwmD6zS2Di5DHoT6CZ1IU
lGb4+TUD2iHP5x5tAZOiMAH+RzfobUYZAigfH/LGTx/wEE05GQmHI9cKn3ufcrzED0yPWy3phPuS
XXDuA4rP7iwZLIXSAMWVLKYP7KhN+jVkdyZC+ySp+KvuIcxvmOuFHMzajGOEKCv+VM8lHFR12zfS
3ibhT0s1ZoqMdk/jZyDPxWm3qKUYwXFrgLClF93ZQ4qcs8i5QFEhMbTe8hmJakucedFbS1sYst7b
UUH3FcynRnM9cr3044Aqov4ltQ3pDVvJ6l+PiPXXnj33ev5lDjMRL4guiX3wemc+HRzzbBcH8+23
aFm1/ipPiLyIaFysDF/ZU6nuqgAoxBXEHmq1+AG3Xvj99S2Zf2757iwPD8UUx2UXHK+FMZvFTxr1
An2NesYtQBPesywBbh1pDvabImYOsA2Gxv+V9CS3dQFtVPZQT+pN004Gahh2RvcrT63+389SkLp0
97VjV2M8WO7AjbwAC+yyGMIK3NZQGd5fVVTyQqnINFHuet2hLi2lPig9ziowL2euyPArkZc1LyZ8
SOz9vfk1Epis36/Cyb+lGZO2qVN3Oe++uVznVOTvk1/j3f8NZ8uylBPQ19zFeNHa0giUjH2X/T7B
95sw+eI0wFFvipizU3m5BBsbjEc7ouZKuQzgAMhxyCNyRFUO3KKpxdglK1RjLa103/8NGcuKn495
7o38ZrIvP+/gfTHMfmDvTjpp96YQ+EJ2fg3RNzGahmdFjZ57Tizoj2iNLjvrxg1GOL6wzIwczIk4
Wa2kCwW2UFO3z6MitLNQ1atUxi8PCJHBpTq4qhl/QV5DsYdiYX2Qi7ejWZoGgbHGHc20gQT0LDwE
6mir+XH1o9ekPzUBkvt8ewxWLBBXOP4EgOdrWdVQxAmvBZ4Did8KlDtUWAK11767kv7PKXswWns5
4PkJUdUnNfj2/TZe97lKq61C//B/Q7e8nPZg2dEh5e7S1RVmj8rnpu0V+agt0d3nsc9KYN8DXJM/
BrWzQTj4De/r8DcfnOINW4CGCnwqMALv4fQoKGfCcnLMKNLg80Oil6UEfRv65uUT1a/py46GrNjr
KV5fg6Be6d2w5GjZj6v+K4gs+djzrViFWkOuhOb6ZFL+GV2pKqU6OGJMKcV2wunNItv6Q2ivNWJI
pcqTZW+KE0fxmPWs79EOQZPrfVwqDhsLFvhjocWiv07qODwJPJq/1sSHDtZ88qox5ge5eWIftIDg
Pc2l15uDdmVehXLuV4hLhVYg03LiHn9G8vj7eM9foSXVrDG3b4oMvMH/pNjScNFJYSL3D3T1dfy2
yXROnvpidxVzmM55sj327ViFsMdCNf5TsE/m7qpxgMj/0lzaqZk+ROMItJV+y54FOrAVpoKJ3ogf
udS5XP0IYZEqjau3Z5HldcX0heg8axdPp00yd0ljRlfPI8F+W57juTsOpOK0ujc3caVwLB3FW4BG
qmeiXnQBV44R64ZYcKqATQHUNoip3pRq3nU1ruvruD3+p6dBrLdln3Mjbe2iZZc66BA6O0CKfvAh
UGxS7ro4L4fddNMyZcPpo1wGMForS46wQnUrEkwAM96ugM5kDXqPrXKVyRdlKuy6K77sbbMlOoIc
RLSFZ+/xx68wCwnCBqt6ute5xh31rK3E+DHiIPdPlwIGg7zht//BkUbeKosonX8cm/HGy7OKY8K3
AUquD2ifSm8mjsO0y8L2ulr6MaWNkKeY4g/itprOmCNg5MJeoDdM7ZJ5y8PuuHUp4vGgvll6j+qR
QcRD/AMnaieZV143dHzFlq+YcGg1oFfMowYpZ77bvNI+LfmYya7Qo3RdGOMQOopr6+qKwvxtE+N0
4oWzjPSWpPXb97oXKGNzAn5Qmvi/RtG4u4R1XK/FmMaDevepc4MPrChG802ISdWrcSYqPIIDgLpi
6g2fyYfezHqJWnBlc4bJ4ma8gMv0ha30sVRa84LUVtDdDQViOtEDgMlSkGdAAzx2tZd5uyAN40MX
yjh2AEEOiJIvyWKlRW51UV+zOGozwSqqxRApoDnKS5DHtOBilMgD6rNMKYrocLjZ5Gg6kWILyqUr
HbgOpQ6Btnz538E+20XAb8MZniDvPbMAJEwJJw1RnKZfv6hhYcq9kjMsU48VUrBCdZIVlnfyepmQ
vL1xMPW+cMHh/eZHnYpxohfp//Lg/6N8tjIrxo6Lq/lxF6YSlR9EUrOHxD76vmLTx5ZGXXBT3zV4
/3uenlSQjhlPDTKKUPSuue1c8PumdRAcOJvcg0jCbcISRLLS5G6/nhPz3dYaypMChye/AKruwy/V
xLcbhAWjqDtnZ267rwr0Pb9WSBAiD/gPwXKAYaxOOWr6VCgYegOl0fyorDq6njb+TItFAQTGELEq
iCZPtSRemmvzcEnH2S1yjHetXJHScrvOmknsO7oEb+2jdKveM8OticmSL6QhY1uhtCWzAvUgPPAt
zzxCqfr2BM2GNe2uMFhQmtVpUht+DNzJFCq4JQbH8AUkKaUXEW07DkHt5XQPPw2L0HqzHINPcWcn
QS5Tjs7PQC1AcoRwnAZqplhIVPmKsVTF5+WpzLuRhYjIXW5BP5xKdS6294sl7bduJQZbWJHoCnkd
kr8FH3jaYppc1UujdB8JaiMildBgi3nEDRh4V8KN/qHpdjKA8w89+9cfLz2Ss+h+u1OrtRqPnfkY
1hCBfSsKZ1mw8w+KGy7Y5X7IMupOcjd68nixRz2at2yIulc5t76/4kX7EgaLdE7dliFTKBOEbvZ2
j0K3O2ZpMq7eKEJ8LogrPLHZKDL1jF0Z8pFsVS6IneTMgnsXdf8VnFDlbFxi/MC9vxWYYWaAU9Si
HELNgkjBv2jIo8kPSa5Qht1z46pBPUfkgm6sbntqix3SK7Bmv1Yja1KuE4vJLKLwp2rofbmompqi
gJC24a9Mu1Jd6+pn2PFbTlhpv8kI/fQDEnfEpF0rXoM2RdkU5DEKk3+4xCsyi3XNLDdyiCfY/FtV
4BFUA0Hi3qF5z3bf9o9TNDiaL/bwtE0Uk+T9Dev5+L+/wrwPTCSSMtXvnrCaodIExg2ezy17yGMH
538kjIuNdI2LRsmkTbini0Ty+McBytc4PxZisrSnlIp5CE1b3KXecL8gWiCdgP0nf63vsKft7pp8
TnZBunhkPPk7+AlgdtEwYciXwM96KQVsFJLMyX84wl3jV1uUrTDUV4xjKwVSclIVotyZ612KXQ7o
lSS2Igxfq81f+yAge7xdu/GcPa7tcDu2ZC5UpVPf+6tAAT/njRyxpanz7zHVjRJ5ULOyVAxb+u+M
dGWVcN+4gltVHWbC0hX2nHnEgbzF3cNCTwCeYTf78gl8G9VRCa3i3Xi9xOvasZEJfWeDSPN+YsHu
x5rJHelaeN3NPaZTynRikdDjNR1qjbJ4jbzeptJh+p+JA8hBl4LQ1JH8aQOF/kXs9ob8btb2g7SY
YJQ+sF8jW6vkSEP5uZ1vtdeLrbIoMMS0ZMQzPiLIes9dL81ATyIc1qXuD09vz3y+CQOx9/22qLyo
nNN1F1bth0WTUtXh+NEemfeP4TpwWL4tR9cLiIAyTZ28+iTa8hh9bsfHOeAG9V8poexk2SwUNtji
BpMPePBl0U+bbTu4o3d0ETeRoXOyYVlPMSNVtzMIFp0R8CwM2BMi4PDBatBcaBIMK12dUhdBzEDT
FYh5OqcKUARoppU/XhJjGyFvdVdtfxzoR16D+wPvikuwOF/JkIv7U+CgngqRzkE390YUooitpgbM
jJJvkl6TbCCbCIBpZMydgGZnohiviKvX1ypJXEeAsEGDpnllSzQo3NZvN/cQMcx+/VHPtfKvk/Sx
kQp061kbsi5zGdGoZCN0O0g+dsl3k2H6o0ihnfakN3EcMKXQj2XKDvDEgbbReRlbnPeiHS/qy6G1
q3HDL0xPNhvhTk4HLLeAC/+ow2fggkEDWDdwUO/tRH8uHJgearpdGLGnX9akao4d27Z0VwMBTmil
FZ8PY2g/0mzcMs0U8iL9QV6ELrQAy/yl9xvOSOEyMNdbG4W2u+8Mgrpas1u2OVGKB8tUsl2AGEAE
PzPekuAYkCfpem8qJDhCodnh0iJYfBn516cXzMEik1HhpREAQfYfDA9fbrM8FfeWvkafUi3Flq09
YW9V6lIc7+4rNL2YULFdnOXOKtJsxYnFlafrcfWYd9vOff2SBiS06EZb1W/bDJjZANi1vIEetKeR
AzKKw5dScHirnnO28wCzE/4VZL6t4KyMwtIN/k3WEejrsYnvKdl7d5/a2qMePcA21odTKFYzc4FH
httv6xSQLl9+3f8H7EFFdEWwtnVpnDc+7WMe8ibke5odu6bfyBYkxWe/kCL+Lbe4rmgWNQhuZV7s
mteDCuhLAFsQjhTpNvImfiSoOPWkBqjhQYXH2EjyKsvRyWA4Tb50c8EBcSbKOW3NSfaJBsZdaG7n
D+u3Eh6fW4IKeRV8oM/bGppCkBC9Hfu6YYnoPgBPJSYxg5Q+sTZFioEGybzRtNxuHKF3aD3ye3KE
8uxetWYWb7C6lfkNVKkfENXGoUjaypq19srd8VNKouPIf4ITz0F8ycMny2smWUDWtBT00k6xwRz6
cHr05zBPXYgt/hQ1ViHXW3c6lmRDHiqK3PEnj7oHf0eckpbvcLr0ggg+JqWPi+A3fXiNsMBqkb4d
BdTVVRBXw3leY7AT9ii4lepwnw5anKqA6ZKgb7s4gpq8e+bfKAH11Kc3T2CNM++OzTGi9AuLeARh
abuBbJVesELSYxCHWW7zwwLyaK56pfa4b/o2bl2XNMW6DyBnXaEgRDbdK1epYd1nTeCKUtPvXV/q
cOKs4nKETlyKPbvTaZZh7ikBO+zIyEkVnAJMvDJc+lZmJmR7mV80tvXjO9ObAiMYFele/gnTuBZb
mupMxA5qTfymoE/rZcJHQK4a4R9e+2MvdMhpHGCQurWIilbzraiBp69xaPIRjEVRhbLDLqyaW12b
aXjhOZCba/IRz69HQaDy0sxpWbAydhwZS7aVIQX6vq9I/t36YffRIuN4liZW6glLvsm/0zQsGUku
qVzPfrJwtVveaH2QM9oCso2yy4L9DSg2XP8UJExW8l0S539hbq2kqH7fUHhQ8XvaoCDGZ+4tLaRq
QJl2rgcRcrd48X/cBm+QeY9b/wSObjo2BxBY2mXz315k9uWIg9areUNNlx+n18gDtyMEV48fPyo8
QjRd9Sor8wupz61Jr+uadM/JlEopC6JRrsJ0QSSKnjvpmzdvVdXKyc8p+dIdOT220AqqRvkDUKVG
aUXx9qwxsbD/8P5sUbX4yMVTyMo8Yeb7wtG5rJSKH4nBxmM2OVI4G5H7Tkg0feLtpVfwTfoKeFga
L95lPd8bwk9iMmB6JSQS2rFEL2vviJA0nWOGgKKTF9B8Z1mm5ngeFDs33WvabVcQb8RXP72VnRhw
W0Uq90fPiEpD1uM7TQ8XxJiEyJfrR2nBYPLBITO7Bda1o7sRFE/FVcnMLTPuuKQ7IB5EpHFgzkFD
TGpR4WjZ6s+7XRAUrpQT0TfEmrBovWS1fCt9shvMW5SIuQt0WR1Kp/vAWgMFl38VmDnyiC3i4F+1
x/heFVqzD861XJX5GwKyX896HnDeucHh+OKSuRR4O/NANmgp4hBgdoYIahVl619DU8o6bcgNRp14
a1qvtbitoNMq8gREDcwVUyphwORppK06PUVVrHsw6kuUzYKdAtLFt9PgQOBR/JpZjRen80P9bn1G
JOIm8trFjv5CjMaBsdrtKChaCZiedTKaue5COxzRmxS5PhPAEVlifY4tvIR1fHeNHWhwexXn5tVR
LRtAfDLOUvoNJbZrPb+y8pOD1aXvDx6kMp0fz5AaOhFAr1n9YmnfNKjjknYEHvNMWj3MnKE4uzQq
CcpPe4Y+uAYjvZTbJn4KGHBC11kSzvmPvHg2Bfqdlq4QIFb/BsLCKc1fAY1cHRLXrbspSlkD1gjl
uaGdk5nA8knSy2LP6HtqAuph95E4wcjlqkaAzuurOp2hLf55wM/mfVoFDNxC40oWusPW+uc05n4w
3NUhWmiYglJ7shh+8bVb9b5CPwpfyRNDS8XSVpKipNkD4fdCtpNiVi6XBn3mbO9O3d05iuNRPgTv
Iok1BdRkkf+0NvhC4X9qAC1tE68imSnCLc6Wi0V7W23rHJwD2T9B4fg1WRkCDq0sHePQLZTHFKxX
H5lH38PATlDh/qUimKWhVYfhCGeXE7OEqDP6rJ0fqmUFFXV4oBh4+8rYlleiIs3cWQsKUhGfiISi
BYJgLcHIwLbMks8/wNFf+ViNjmcpb0uR5pBK1i4uUclZR4GKnZN1+mslr0n/p5ed/sbs4l1ZA8kQ
VaOWyZzYS62M0E72BoM/xhRJQH74T1oHevhbxmE0bz0YoEiIoYCfZMPrG3XpGcpfkjUVyc6mbuy1
+NvX9sKsrMC2AlJ0dIYvY0uNqSVmtspPutpz+8XFq2Uc6AAfi4ViawERmCkjxQzXQfuVyhYqEWap
Xh24pr72qlVUp91f8SmP+rCY9TyKYG+SLM9LWRvft7fxi4LZ9NDzu1Gw7BLXnjYZPImjO0dffQM1
cs8JeGVIZF/21uYBCLjsPbeGlCEeZ3jTacHqK7k+8R5H9j8aISU6dSo33X/YY8PpaXvBFkqQX/Tm
4BLIMfkl7evDfhopBUZHsTtSeM0AOilPnDuu0s51tMmVoQ+4oj3qt/Z37gJmdwNK+qa9amEHyA30
ZW9JSu6H55qlPDPHO9q0S1w10fu4lbBEiYy484AmGT5fGlDlOOXROMyLUgijZjiQ8/grawf7XzU6
bjlguvD4OIr2f5ARLVOl9KV6r9Gr2fy18TRkExw8RSdRqbhUXb+Jgiiz0YpLaAmPDODxFOusn6wI
ZIirOALC/Q7u/ja+mvMreXyez/HBzYJWsuM1ZaKZ9uIuo08UPzi1CSE1d9Ta4AlQzvdnb5ufjQ4k
cOfl65TBbqKPoUxPmmRb/E+Vhzg3BQ6tvD2qNLKVBDsornhrpaG7PIFoZ3/sNeFA3mKZBFjxBTns
V2QaWIt+geR7+nIEL3Nx5BMQqJGj8w/h96IqMULxOJ2pR56p4C7exHLgGe0GG7BHxmMkECpRrble
BbjpFl0cq9gkA7CkfFlLfI+dbiHCZvL7XGeszohZ2f0UJznofHCBycO/Slt8s6ztahE13RGuiLxs
0LP7552QREEjHJyniGeGoyq7IXozs0v//RtsPNVc4kO2lq3o9me4ljAmUmp5XLQ+DjORKA2cT3DU
lfGkze4g3uKtbcEnzjQq8e4pGgpCp1b6aHGQmocwRxgJWB1KAnrfwqGtMnazv0KcD7COCjeouy90
7jCFRPK5URsXZwFXjKa09umXPG5hEIeBJ910kjIivMWwZ8tEIcWr7xmvWwIbWdaDDGWFeevjDvE9
Ic1AiTebaJLZl6pv7pZQem+vTJbFG+qebwTcUt/zOEIMUeTUbcgAuBCZdrcQ59E3Goydb3vl4WVa
0rZQbO0RbuKGgFh5qaq0SbWHzu6UfH+uB9qFFzHry9jBl6rdw0OQv3bcKTl3C7m5vTNs9cY2FMRM
E0dbaYHZDch0yEg+m3eD/7oMXjNc+k07u0ruFRet/B4GvThpY5enLP5XC3H4MS3UGL1hboa1JRIv
mWbatSmIaDLIeyH7LVtq181M4AOzyiUtdTvAVoVIw50uz5TAcMvafWCvUe5NVmEUKENhiPNaQWVQ
jSEs2DOEqbnfZBiMl7NKIkbG4VVz4biJsdOi/2sS9scT5umhOmv+caixFtQnsHB5pMPC3Ni2btf2
3y4EIJPTp8wZPxhQ9bZTxSlXyNPxW50t7HPu1bM7YvQNBwxPd8E+4mxnUz4Z3hEZ9zlTg0tJX33B
798XDTn8TGc/PtMDL4Ur8G2kNZ4TPaicSjKErXCwRVkQBN5vKncH4in/05keYBekO3fod4VxhgLK
Qgk3MVITb1peZxfHRZZt13eLSJupa5+e2tN1Y3qKOESuJlSPriMh9xk3GnVrVGnQYDTHO9vCRTiJ
ocljF7AdNF7fYmzq/YgaxsRhChoiRRiQLYhnud6uh4EhV37INxtr8XfgybPCFYOUL9HDIztFZTsV
45T8zDP13RbeNy39qi5KDcdVBBDwloj9tR40oc625qdLF5+2x+eLCTmKNA5GjsFetroSUHC2iADu
uFN+NAH1v4kf8cU2SByt7cw7ZkaYqGMj9OaREHy8V/cQno6f0IjTF0IFkvKP9F1zoxby2zee7CrZ
fgoSQ9TgGorlYvIUB+grqleZxN4RNRmaz3fACEzfqgniJFXzxpJFjYtiECmDfnd7BGwyVRTLkwM3
xaElGWBBU2Ml7QxWOxMdmSIK4LtuvhiuMvKzWI2TqbkZln10CuHs5wQ+1gALhNwy7lWsq86VeFp4
l4yviq5BNhCWCcD291LMj0gXNJRpjwi2gRQaKk7nB729CJM+tlQ6JLMgU3EryalL8h8oFM6Zo3lw
1rhBoB7Xmiz6+ObhxuPNA6uJuC1g1WxTGBsIvqGi8qt5LZE1Rea2j6Nh4+o3UD0uTpxTz+586uMn
r6rX+EMFN56VDeoNfCs0NXvgv1hBsm2V+ZbeyS6OZdelfLK0AN+KmtN07ScAS28QGIPfUL66UCXY
uJnfxaCzciYYJEC3IsNBRio0bCXg4iS0U5xpjb/2X6DTbjSE65FCoQ/cuODfHuOl49EHN3dyOxWs
9SaeaJxmZ3wcv6hjKrIgPM393H9Yph8T9KAqioHGP8ag3YY6iSQ0oiQIGIrI8EjVTVg5ARwCpBeJ
9Me1pMwq1+QUzvItGmifmH5Bg3zJlmNT0s8FIFUPm2bnt50XQLBkx1mehpnQw+G8VBVqzW66dtfs
CGTE21CkNctm0RHXSwaH1KjOTEmDjCkHh1qQe8a89QkjmwgnDvLGl9DNtoYdpAPkgBHZEFRVhRsl
UVUylGUNB49E6WvLy8x6ijpH55eDgzDrWTZCxgEJnTxNOFjdz84RQOMHJFIMQ7M1RUbzWMrRYEHK
fjEjrn9w6W2HwSRq7+5dNa/sWqm2+RDM+oto9qOgT9LqBARAZ6ZBwdxPpus3G3CAfjyXX1LwGLRw
TOhn9bYwYak1Gv6nPN64+VB2tWVVCsWy168Js8n4rDe8tpxe0n6JxfzO4y8EgxciFihKK6rpcKx8
0R5+k1KK9IS25S53aEOmDvmd+2UEnjCpBklj+rx3K4QryV/hh2Dmnv9l069G8cxb/iD1lBhVLrOp
BcgD0RdPwyYxDf4KQzDqrZSs/vbIc08ZX+yEEr93bcNR/RBmigp9kkeyt0KymN4iT/9zvSdZ7dC0
tsSyT9BNUYPfmk52fOCbjH1JwFAQeRXGFmmu0MDxzg+1juMeJXeGOUt6NwPwq/73oTILt+IPzpCY
mEEkJEtzYXQDGLeilYyPrPK6Gp4stIvtzqbByNpI3P1IBzXRMjhwiX6CmfPX7bVaRp9fAp+KmKR7
+hm5y7CGXXjFA5rI4/ayls4q6vA9FLqvQMorDLM5Ab4sq+H/nQxfeATGDbgtdkpfs7invcQQMUiK
H9HA8fXs5MgpslOpwMZXyuCwaWpGP29P3i2GlnJ7/uywTXku6kTiCQi350zSH9A/sd4ehlzXBqyT
l2FpyKaImb6Qqz5xqxRN0LyWEHEgScBfHP+JWwDUfDgu3VgyPQYKOoPn1AdK6Z+UBb6k2RpyLIyT
12u1LM5WztmFL9XZy2unms1arAsgg0Ox93I3EugOc/Vq47usqrD50Ed/6uPpVUXMv3RZEq6Wh98Y
c6XmZFXWVAEHZ51MI5yywenRLmSQ8RXEOApBBu5YqLqEDK0o7u6fS3och+1Rw0mpMwoydQda9FTv
/xHcIpkQqG3SXS3xBZQudPjiaJiICwXDV5RKg25//Tp2yU5hm9B2v/cUSk0L5h4b1XdElcqD+zQ0
mxRQybXMVmZ4cNF/MlVHg6pdaBSSL6YR9NQPVt1K+xuC75xt0B1DjTWBC43UbrJkBHrk6BPNsh39
QmYio2B6aXZFf5OQhQHHTT0CHqFS5iDxidiAQk4kvvut4ULvrGy/jI/VCGzcTvxF8m+3RsNQ0k+h
fPEXS44hm29sn9oXt5D9r2lEADNI1PuVW10zMu/8niI3asDEDCjKuTkNZfTY1JY97rrcyOAOMAbd
S5/tuRz2pEJyUWcG8tdzSmjHwCyJNmp8ZhffVy5ue4SxZsDQ60XSGipY2eZ+0KXh7+3+89rIgIQi
VSlIZthX9PHM8z48lHWTpTQor4SA0JchaoAFJk2c2sVktvfp59uYZDLarn4vfQTXXs7gZvahZhmH
YHU5uzpSUobDRHIIFvtN37dEH7msiVQWyNHU6xOVjQ1IqbNtqSO2of5QdKmK0QNmTCvj2LBY0IRt
JQEFF2twNwR8QQLCSKNriKEkGkAepxedKGBBxnohCTA4pJVAnRPaaOsO8BJPdwAkUAhr2MqR8CF3
qzuYpKonIE2PAehzDUvszh4CfNt1E60HrIuWxGr0Lz6bSaVe87btL3J8HIPrr4U1t5HcuzOOEUzZ
G57etbdeqpBO6NQdrL7itUyNcAPoaRoHRd3VQMEXNvmbpFmayI1FHttCHylu5R1Lv6xfZqTquBAu
fAPVybOdnWf5wk9YMeKTq+mCTYLQtHP81gm6/nSSTcGwTEfD2lcDBwmdkgLI39PBeQyHUn54n6Qk
De4J5FybrqYXFgIVzQ73c85qhHzvV26HdnxVjjePYMiWot1ZajxNqBQtyuV7XeUind5AAFs+mo8m
eVa2x3I01N+/p8AENdhf4FGYu4yBgRfH6EK+Qaz51LKbl2OCqUG2hDK9xLoZmmuUfThtDthoN0dR
iapPwhfB5yWJxVL8gyVdcNXcp9c2jzGafk2a6CYUkxZ98IkXa8iPbICBNBnlzAYvlXVwmSetRhxS
i3Tw2gkc2GlRA2yxd82jxd8b6gLs86AuQ4ATCa/rYv410/+eRAai3vUvLbMlXUjvxxL/cTyyt7So
SaVRy+I7HD5daT0WYrfVUc17EXB3cZUvDR8x2QrtT9ltRGS6j5Jqk/SHdBVYUZbGzAMaRyuIQe21
G5pYY7viQJ5UHMjvgcYhZc3j95sFkhspvGnEn+ofGpT8046dyP6QMIfMAaglpi0aC/mj+ZOkxkYA
UkHm+GuVAlQIi+jt6nfY8kHcbuYx/kGDa+5lQ1TWpjUtgOTqKiVPZjHnENRtnAjSRIfh23duzjQI
JkcVfK1TNBYdMjhYAi/QdWJab6+aASY6SzHE19J5xYhZgOETqlLXFOSXrhP7v90g7SinF0cXGlbK
gsJuVUOBihT9XtqvyvfG0OsA0Ax3uugCRLuPQrLKeIdv+REwTUddMecc8ZIpcsSIEZk3Ghi/oX9r
VCQSL88iGj59LS8Y2Oztj3X15WnZ1QdZwzyaueAZctX73+f1oIgvLZ4ZpQqlxhTvLQecDR0jX+o8
nja6Gu6Thsz4UviC4m5YS1JtE/0K+FTxAL8jlaPrTQihzN8hP9cv4fagvt3cElQX0WpHI5iY4o8K
ULum3ZaPBfUITQjia7/Am4vY0EbJpRtPfYWa8T1wrDo5ApDfuA7uhDTP6dWFcFCtaZHOuJYasb2H
YsrucnrgOglwmye3fJZv9M477XwPHPFgajtg484ztqkrYNvD3s8vyzNrAliGku+c1oa7895Rb22U
BWzFVEiNMUG8JyEHFrf3oY/MMhkfQ6lRm38AcVK4CsDd9qbzMnsmT3SffRQkINPdJK9hWykTHsZz
PWpaFEtXIItjjEQNjiE+gXeXWK9mneGh3KFbbNprOGKnei95K7KFC1hz1GYsJApa8ttJQ6RtlEyB
NnsRPwti23VFKda9AwNpoK7/nLy9l4amb93S6Ljz35dSm6Pm1Dr3uv42eNh7HmYF5KD5Cu9z+4/w
w4wEzjCHaM86wHsBcPY2pyQ5Ft2hDVOg8x0xFwDC5Yd5J5fPFBIHYN70qiiEPE1yQEQ0c7ZPFnDE
JYHEatClqRMwWKOP9DiZmhSdqclgD7Kd+HzZK+1IP2VPlyT/RJR1eaWgezwcQUch0EARk8acFnIb
I4x3JmwLmqF6qKwhcVanpUXQXsz1HQXC5RnmF+LL5l0LjHvXLKUhM0nAAinoevpx+uwkQJyZQ2eF
cGWu1xK5pegRbH7PWs8lurLhKqL5jn6K9uTS64ttKb0ukDJmCK5VfqF4DxcfkE682aa0Ks2eBm9m
bdA2J+XJUgm/7CrXgaYvDjFOyud7EFP2HmsLD1MZzaXBU6TEg1GqB6oJ4eiw9F/AIOXuB1tj/xnh
AgeYgqcFiYmoE4i8Gn6WLC1AhuclDVo69lzDRDqw61gawLeOiZ/HR7G6i6MPZRoFjVC41g0oMShH
7+78GiAsc38/pTO+MLWLF0/q2XHpesyiwTttjePHfrDoCpUoB16622RDonQvHQ/ow3bXwsrM1Qeg
c/9iiDRPhWLsl8jGeeGRvhpjSiOEIREiC+wcy/QGpVN71SydvLuA1JQ6y00PmF6CT13oo8XhfdLs
RiRMIwuxUy01IJDcuymVZ9eAM00g7asLsMf7nBMvKaB7AJenMPCv7H/zuCojo0FSRy8aRTGB0DmF
eBfWahR5obUI78DDs4Qxlu+W+BbE/H+iX7Ln9Sp0dIPrXPEcG6WNP1+JS7Ht3QckbrOEiK+gOBp2
TNr4swYRdZXfh+vyYASEn7z0h6cGJObFMG96kNVOsuoHM4uq5NpMnJkQKFz+aIVq0uaR3/kFVKBP
NbetEKPQWZmgpQ/nkAcj6mOi9ss7vRgL3zpXN/OTvNSyI5h3951hyDpX7aCX9WVVTZUlecOaLGmt
GskD0oiUWfdOU1NRFlNZNjKm6HrQyZDgwCgFckWrttxHvEzyo56/Y+f5DUZH2sXMRAWL6QhpiJYU
lV8sXDd1Hcx3hqBc6F/tFZG1q7JpwytzRcgrV4SLgeKL33oMoZ78HFWsmM5c94j+ZrvYTJiDRIiW
qjUfIxNL3bIHGMDZYwexNXv8dGW7KMDwC/5dusGdn3//IPJqsd8EAOptawXC0I6QVXFg8gLpQSmf
KtDw1fRHGrl5Dpn/AyHgpm5t01mWLyrS1uVAXAFjnq3ho3VInaNGMX8Jm3PhAkoLYm8xqCp+yje3
xW32SV7A7SoBfxpzg/bSktTnnHYm5ftu9zYLQwR3QU+y5oqW8E6MsAu6Cidl6fwjUCuFFoSjQwZ3
blfbNhWszahTDQxiL/E4WUa6Ujy4wlXlJ58MM8Z1KV3u6rySFWYqsc00E2u6s44ZorBr9oDNMX44
ke3vFWQz3SQX/bEpKT0B9U7ytkt+PniTbt+PKvmQ0Q4wpAYUwO4NLTQzk4oUyTD1lEn8BPnGzcv5
Ymws7rij9CNhBqu7p7XdGIe7tBUPyGPuSYZZNps75DyDlEm6LOidd5mzzMp63FtQ4EpNNgmbDky+
WszpqPk57FUi0TLw1ZnWt4B3XVQZiO53SEhYd6edpCv12DL6t2qIeL86HcCFQ/ZhPLeZDfoawNqf
ipu8fJTZCQwTLhY8+N4fcs142QiT0sm88Axa0XIArJHtmFj2WcD92dMUYVH42mWogBD/7LLQHiWF
2+MeSpFj8bYd0yzo/CfWJIfsMDMeb47HS0dMC4HqHFYLoe/rM45O8hUVZC0NwuE5IGpaoxdT9C3C
GnIntiYsN3s/zA7FGyKm20/VgxMTOSwjbEWaCDPsnpq0SgZmRW/XruIAIqdxZVOBPD1W7HJiTYKu
dUg+vthkzw6RTvhKXTViNr1aDcmNBX4FmdHqSkEzx3vRD1RhI2SWoetgRkg2IZPnI0G+gYIUBTMv
ZxDLUoU8DwatqntDujBaeYJxr/QhFUMFVLCOmSTk9ANVM+9QM1ZsEp3IAX5anYpVBX3vdKeTGT3t
ntWDijVO14br3QZk+oY7BK11HDqI8qnBm3wnA3puF239UJzKeJJ6AVgQjbyJ4xttJDRYPpNKXYtV
wUwP1aGGJc6fWLfzPjXC9HrE+HPcqLLVorqQlXb2xS2/lN91q627b9rILowgh0TZJIBxhQo1hAUq
Rjnd0JunRJifx96FG19/q2Q6hpTwWYvp0oE5ptf5VkSeNVAkzVlxk6K3TnkNNvZacyEy2fMVgi8R
jIHN8p6x6gL9gCIlZUyEDgDuM0VEEjiHDRz4cqdM+QKQ0f5XlsplBStd8ZYfkGoL9KY6S4Dy95eA
T/ZRWif98KVb+KUgM9sRmATA4SBMTsSLguAE72kJolKV3+qyIqIrYHn4I8iuatp/FytW3e5qqDcF
kKnDxgathmFGCz1LJAqC+b8DRmTh6j3db72/+uH55P7obS0OYlLs/xXpayTuEOuoN4uwi4Eqsjpw
sRf55Gw2KGHmFwo3fFQ44ceJknzEV4uJpB+qtRrjN/tnLjsrWZNIcqUQDsLuuxO/6P6615T1Z+Bq
8yrm7CXXEO8s6HVz0C06XDPttmr40ZCdUpnQyZs6iNJvGuo6CDv60ARHBrokyxlxoOJ51jbnzh9D
CdxRR1lpKoBAQTkj6iqTqi1Kr9jzr/wf5Lp0yxv9YyeyTgw2Tc2Ee/JVY6ag3LjjDp+YoAoSQjbL
USFyo/byUCK6gJbRb1tX9+86KEtAyVV/AQgmH2CLvAHRMt8jyyg0NMir0ClW3KgFgFhDH8iiXRMY
S7UxvnPrkIhF9UDUPNp5gBrTb1xlNLpfW5n/gl0UxgSEI8YVIibxX2UubphXXrgludklSmIEX1W+
DT379LDDnnNiwc4uBRjgCABEiM7Lgpco6HAM4dqaOcLCI0sSQaCn6iAasBp1kCIw3Z3UNynE9JYP
8nAe1fcycoDFZOaE/nyx6K3rYgD+WXFLd9TcpwG72GRggEs8C1vKiHJPWpd86KQu5qiesWjC4gki
5zsIQmtpn1CqCrrcbi4VmupEYw2hFnOrp015Vfls3I6U5M+amuZoanrdTjrk9sPvGa934YL+QtUj
9CBPq97RuUJhb+z6UBf/bQBcDfDAYl3T1Syypj+w2yoiKW+drBhr82kpj2vXDhayuhoG4aZTM/dj
2+6Om3JoVIaidwdjBNRYtKtuF2FGJXdIXYRNSjrVQpclOGatuEoxkS98/AKSwCI3MM7sNJUFj4n4
1PJhn/2wYPXifNR7RPH+kw/e+dBSnlklFEzshpzdJ8BF6oPBvDBzSvuyHCaunFX/PM8g4m1hVba7
4C0AQ/6xHRx3560pECRh4ZpUj2Kpp9lQ0CQqFX/+I7J5SqrVz/Vi6Ugsxf+0Ft1nJCnzLxX7IvEL
4AewtGF4Gmit2eLSWQaeIzH1x7qxHI0gofosaXoW9fV322EUctlUzAwSoxics+LOiT4ikQid7ktJ
W/tpT5sCPVxu7gLQii+T2UcMBX3BN6zudurQfz6GTrQZx0gqINmNF7UvR/F69k1eqMNxBYYwbFhB
NpFKkoOpPgW4PXD48+R58TJ3VkTZdyv4w8IP7Op4RoDqmao1AL7iZUjijPoUzaNUH5Tziblg4cJi
P0hcwiapsca5F6SE4e1WrcY2OSizp5COHvPfr6bE1Yyh/AObvofKSa0cUXrMUjyfpkN5s5bBjzmq
R+Rso8XkCFNOwz4hQCF+Vgw94aQnCJgkr9GH/OaZv4/TMNxnStOAWa6MvwCCs91x1DbTQMyC9jYv
YEEIYzTaoYZUL8G0UHwRaJtOdnYNfwkzylJIXCyJW3QlqEnKreundHaf6LRjG3K36qk2Npq7K9zB
e6Z0RduT2wZqmteG3q+z5XRtlrTwXdzR/tzqGGcS9/Gx5i9liXdhulYVW3NRmx1CDTkztQz4My4p
iRfPmIdWLLyqHfdj1+J1IonXqp4Afj7zr4D1l9yakySA7lFe62fD2g0Ye6c+aLYw6LHxfXhCtqJM
pWds+jkM4OIJJUKtmQkfraOnXuDk/6r8jnN/3LyDjNiOPr7bHlbgvYadj1+41Wlu3vryjX13qEmk
7UOwI32vCfya4P4mlrMMDIL4D5NB8qvDAYSaGmWlhskmz4c1Oir6ukF3kGbIzkvtcLX2Yw+/nQms
7+EkaTiqAcj/Cmy8POCGs8J8A/vej5Ua/AG+tnIf3of1Kp+/BXiOsCIT4A2+RDEvpvSKmmniPCpZ
irTczFLRHwT1H8MiW6BVLrYSYfoCTQ7j2uhfovyQITUNP2jBcl36HGIgp0o6CIKfiobN3n7uDOgw
YQsXEGIMsjSO4G+/0Pfv0/CwfXs9EkVqCdPMVamYXTsbg7h/OA6P29UZ1+OMtbHQTod6+UQpjMOt
XUNEDTM+qgsCT8WrbMCjJF9/xcSLaVm303whCJtrSYPDLAdUXquybfEzzjD5dhBZP7q9S92Vzl7P
3eu1fZdJ7idOwtkcTQ6nAgDbhxIxxibhp8tq3NNGAjpLXvu4dtTH0ixvAkGZJCb93ny6SHg2J/l9
VD4yKozJNiXMZLfMhRPRiOP7vpDRwT3uDAfRM1YkYdd713fdf0zmyy+O74U/A1CQ/NMjbRtPvUCj
jy+Ppaz3cgWpNYLJPAUp0TriRmOWAWxqkdrHlq8MW2tXjZzgiQLOc4IgldpIOl75R3bmokLQcDIx
QDIDmOhb7pIQCS/QGxiolfcPgziX6YSWpB3z8/4ekuxnbLd14pKgOmF/bjx+v2v73KaPhk61ccTp
jg0G5hp0hnOcCghd28drKLwp2+ZVajWWTRVtp7KnbhyH6xbF9ekuPY4+rz6SksrRAFHRU215lAXj
A8FyAlFDP5w+2MkTcvQqOAfpsUyBBooaozXDgbnHNY0tGYPfIebaa0uwa/84W+4+lgsoWrO3JqHJ
icCrzWzrSU+YKgYnBa70NUNC1CU+DD1KYFd9d7alwNhFJz2PsBhIX7tXtfVyJSZtPcijgXNCxeIV
Yml6+pddnZ9ol1fsOLRC8VIC4bPAVxt3Dt+ADG0VHhujIykMvEekckHs8kVYmXBsb7EkErH0iE6W
7Lv3m8PjLNw3NGleeZ5JVQxVeehb3gUQVmguD2OmShjiTIfvfh+gjWrM+CZOX4Z9iTmaHJ6Evl7A
/+uQafkSay6jlnFnn0ZdQncDxDi0in2o2nLpPVnLfwB/nTjmavxcEk1eoBeiaL6UuRvyoK73Jvcp
3nSkeXL2UhjIlNob9gca8aDvYbYVImmSmfMz/Jl0dbYpI9XYxbCDade05+OoqPo591IYWPMv4FUI
nCcFLVowzW1q41SpTICOzopDqIioNO9KBtwJqQgrf+qmUk7MlUkg87y/8OaMStaNMHvo0vryF/Bl
xKLy5xoTAvD2fAITGvPkszv+2nBd0DdJPueUI60Vvtv4KNvCbOwn9hSgEXa4h1iLG+0GLrPpYO4r
PQCSJo2EyXSCQ7ZqJyJp8bOStf4znzCUa4+pJIarvq0F3YwMTZleb4uf8xGwZ2va/GLup/EPuZ2C
QVNIxrqyWo0NCTdjb/jCo8y50bKZ0SW2I3GrUPbCcz//j98fMOE7OamRVPb7iRo/wbRU9xOpYYFC
01RO2bxMDYq+0n+X6I5zrmFOhspQSOZfl12lLvNeI2io5YEBP3xGjpZ4BpFMaSUi0MQTAtVhZ4WI
JS895FAXMLxGLudwjbi3156D7dg0+TMdMPI8umlgKPEr8G5kKEFILeixbRQXSSHoi0AeWBgwsWDl
nxswqz4vjJ2QwGc7RDneiqWujVt4GhO4YAXGD7I95p7WBN0By430awq73H+1VJjmQVl2UvbpCepi
QRGNu2Ny16eY+cjoNLONPHPvFrg6Uppt28r/tDLD/WcvRlbtO1wPCT05FggzLWPwtR90WCJqwOtW
Twwm4beMN9U5gv8tH2x7aESt26RqfIpI/W9DNNOPm+GfedNppm1FEUXqx8U1/KFxnJdTh37A7q3x
bMFds52/Xip/qjvItv2KTafdAJpFN22A/NRjizKYgOXfWxiIYHIEsFIcdqMBIgTYD3i65pSKeSUh
2EZGtBD956XghmaRkKgJxBiwF+5DxDBTxfgjM0Eqev70783vRfCC4i7prBhbNzJnFVSLzD8pa+y5
vUE4404pZwZUbOX8/WK7+yw/OX9ucplcA4IoOVYpM2paKgUR3Rz5Aqfo4S19syUN2mI17Z2fHHUl
S8xO9Q9WK3IHovGS10MEX3nR+XaItrw821gkc+1VSxTOZr5+t7lYTdek9A+ZgX1/3lGyPNCOANPU
C+vjRfhmv8MgKtaI3JlrgVEymv+DRwdzRxfWVwnA7zlavJgZvL4FJ71dZDa3nTzu+6TS0CTqU+JU
Yufub8pJ5AO1fqGJd80JfP3r7ii8jzBjgOe4hBjhouDp6t7e8MfXa3q0TTvqxcVHX2v3ka2VGVi7
x7qwMYQel/FWglvEXE9zjMb33IqO55XPYXGO1lcLJlrh3CTsYXFjOdRtDX+sXaJe6vmGdOgIN+JC
Rf4c87JfyFVkCTwgun85aj3D4KdqURriteMhBeqhgu4T1+WwIYg/uNI9yO8GYqukuY7COII4kSV3
JRVSzFEBtMc9mPDz7jzcVedBTAiqCyayFaKqEZ3HZNNH0Px37c18KGfh5DwjYJB3sqyJ2x7ZsuUG
GhcTkjvkE5hyoEK9uoiEHA2+BIuEYdxtOkE5ei4dO2p3ebV6oB0aYxFAYL5+3G+idoS0KCvxOR+v
DBJ+B38q2dBF4zUU8YY1f5j4XQWWYYroZOdCn6WnC2UN50NvPhwoQSra6DeDS3nGRmcgUH3vSjX9
/WujIsWNUS6644XojbAmOjU690X8O63bBckY1mNyeDPjmJTND/49ol+SlVF7Dm8J5S5u2jn50++e
vYL8LNfm4ez2Qm8I23iLw01YmOewAkF2RFvYW9uIS1Kz/DGdp0GOSL0SAM8iRkrOE3JPHuIrWJS3
Rz5V4LanfYVKFHlt2JvUriGYusl8Vhn5vy/HiehZQbn0HCECpbM7+vXDVUSDd5v4FXi6uVd6+pxz
U3DHhqeBrU2jUCByYT6Id7vkPQ+1RDBF8zrZn19Xg0uycA/sp6PXoR5/BLHSPnvZtMmOBSua/X5N
iwcFd23WVTjH3e/Wk10T1wUKgoE9rnrERK84O3eOdRKpfhCXxzz6ohBj9f7xy/j09/pCEkr9Bt6p
Vk/Bi2EC7NHVfTI6Ydkbq6nq2V4bNK8RFBr2KD0vb5jKfA5bIffu8NtHdj+4D+I2feYtzLAZs6zh
D1iS5hqJ9MNJBg4P1ZQ7tods4vPuTJFRIy9Z/DE4/buaNkNghF1BPRZH+bRk/dsIjXGzIoMJYAX6
bwZj+HEgeaS8Iykz2KH82qqXAIRE08ge1s9zm0tZWLTx9b7Yy6gC2wUX3gOaotqpP6F5RfbPbgDE
TPCxxG/PxIpi+01F4EDotevldadOgY0edht8JB0Yt6poFK69CO3YJtU+Dvf84YMatyPP70ZBDtuF
1oCt7Va69DGQwxThlkwqaG7TrXCJehs7TIBrmdx22uAu0LI+mrOIhvBRpb5PsQHkktdsn+VjNkO3
k8ta1eZOy1VoyHZ+642TJNFIpyo/fr5Ho57PLGeQiVuHjoeQZ/ZXinVfz948PZwSpFIKZBBxNDKy
NACDEwsGpxn8m/hJRRGyOr/WIitQPCA1H/hq+YJ2jAOy1nZucM15emmiqnKSUayZppSouVzUCL8h
tPMkIp9VhFZc8r6cYI45GjnTn1Q5m+r5kbofXoIzB+zNgK/X4GJRAlTMkAADfb2pVOp7iQND5B1u
ntKeR1eWrp1Sx7cv2rU485zar+vleOY2YzWBdfRY6TPvYSqRkfI6zSYfZaiY79su+fmBrwr7TqLC
nDGl+WHzmL8eB0TuSCGOoLIdrxKSLlgS23dwiUwIM8jEoaLe+SRg0hK09uuZXzTW8T5hTbT3GxdD
GAW7mQkyYzq4WL/fEXWz5LrMjl+TSB/cs8ZE9tO8hxL2+iyQHuiMHoEWZDRNLwg0szYccllxwZm8
UG2AGgvoPsV8wDCSe+HDDAwjaktlc9N/ybGIAPk6+jTxdKee5QSvRnOU4bmugwPUmKzpqbDF2OFe
aym/Hcpo43CtJlbeUwIkxaI5pGfleojYC/X8oPJQW0wWxxl4RGcqE/4+xpUHdMU69j3e94T6p5E1
B0IHPHivH+tcPtGHId4Yi3FPCX8ty+vHWWPj0KBnxIR/Ue1axcCdWJQQD7RSC3JNMvsCA2TFsz69
U8Tq9NP1yiSnNeTq3ijx7h+loiagTXjP+UoQOto3xQMhIn+pusojjZGRNwLivb/rdtIoW9EpYTwL
cWQtur2NadchCCYANnEqwB8ZI0XFJmoc1Maxvays/PqKr33BYAWI2YB0Y8iwWSne6xzlFU5s/SDD
Z8qcAla5qf/gZMVJJafM1my7uCHT+lIgHTyXkQkRkOEODxga9WNQKvyGsOX0p9vX+mp/rr7Wt+9f
6EtzFkTI+uTvml49n4oZd2XNoeuUjO6u76ca2j6fOL4S23Vv6DjHy24L3d4ZiO6leqKSM02Kuwne
AslySFvwzQSZRINihzs6uVPT9kBkj8jo2U/kxS7tEA7+GCzoGZzl7eSOAuwPxKykiMwkk9B1gPAi
Exke3mi9LsHibEO/ZtL9mhMVtSGyncFd2dWnXxlE2JDnskFUHrhYk+V9T05VVfMG13EpfJ5MGyRP
QJgxzyi6rgenjyfqKNpaHC4KMcgvB1xQJIUHQ17JNxLHzQL1/F+vFlhke7VhmFRIb0YIxAhlnJa+
JtLWppjsRnRVi07EBRaeKXapTwTYaWZQBVILY3tK2vQO+oKObgWZL6i3wH1YzXCXUAK7OEylqlCB
WNieJiZmINr91K0cEh3WClSpu4hKzWmOrzdUFyBiIDmq3PWhHhq+7HZgn52cqEU56hbzkWz6LQA/
dSbxyvwFs9o4MQBDmmSsnX0iC9VGnDQmFuhqY1ikIk+pVbv9TXQwlyF1fDOSmemjKZla/kQmhXqZ
IOYEMq7g98ArfqBEHw9DetS4i/DPxIH4UlKw0X3wl84VPPj75JXet3+gHyB9tjbeHqoiH3sk63RY
jL5tU7UmEbMovg0ghNmaUtC1zHin+Q/2C7wlPxvQkvB8qTCs+0t5WW2fEYZPgrgom4whpcVHuKFS
aL4GxqofvlpGBzGjwdH1GB4sGfrBtnq36GaT5L7O0H3dmgiAoaz1xFD0zb6JRTU6iwAlw2/ujk22
gXHBKLPr2qlmGUodqpZA+UtWQHsQt1f+SSWyDCnVUJk77cI+ddGBbL01lUfL5F4HgB7iSyKRWMT5
uYeuYfy+i1KfCOBRY3/UuCaMHcvLNfxmuXYAlCOzxCXAFA2wcaGZnMJqRYuuCyVENAkkPP+/FTf2
yaGkaW7l4y8zWgp1pUTPZzAY7I7l/FWV+8umjyU2/Yq22xEygugl/Tx6+8E6Sz9JV39RbxdRlDWG
zOAtGwKiRQvjxVqlbWXtqImSBcm7p3spqdALQ3hgDIfXeVP2hcPNZZCmxu8sep1U/XQn8a+DwLY8
O0MpzReB8VvLoOFntBjK6dcmtJIhVTTFn6GkVccsVwqmfFqIb+x4WGnMpt6gKFOwcwZApCuktnby
VEexgc/hmFREgDu1TDCR0SLZl+jD455+8pVCzlttslOHbJKsRPnmfpAbl8wcJPaZUflG+sSNBm/G
XY+gUMnW6bvgiY3kqjOlvKiFNURkpvsDxrv1l4V8sx1QXGKAuDJryabPhORhZogS87vVKEmy/VhO
4VqYDdw/gnVd+72uBdiaxiwVedmK04o59a6OaSmcd415WEYdkNF7UcwQ4R7CuolMGblEYKCP8ZkT
I1tOoFjT1gsB1iN0avQsKUNeew0bv9tbqUHtwaC5vC+OAbvXpMy93YbtLu2NQIvJlesHrmx8mmGD
yWRtjRNZLUWCMaP/zC+4lqRxOe98V64htWDw6pHoNX+zO6eqI+J9gIH2zQG4Kl4U6UhzxBqUSysN
dmnncHraUyBnzXv5CzcsjOu9G4SDgllaWTwKIB+syiiTVGnPe4KA6UmoQye/aNwPzljFeOtfusCe
W45IgQ9NM3u5BpiXiwbGahSHn+2ryRRTHJ3gAR3bAWqbiWOvObUDESK0lPkPyYj9ZnD5ETpe5Jjf
GvZGBSE8xaDysClcTG4QzZEEfQIxPeOgGHLqFOrObt3VX+hPO0Zn3mHc8VTWaZZtKrEkmqxFZ/Jw
y+H/uZdGu/qqsC61obYUHETQ47rCuZ1Qyw77Rx9f24fluJCgBkY5WJUNXuwhPtBqfKw9FzRQ4A1v
wpNSxrsTVOlZU34eGUnGhI0BPOKsF+pHOSIVWb/D9EYP/6y5IIsLnn2hG4JqQHexnTetTMRwmLrq
llZypK/De+ThIAuyPsoy0Rcn3WK2yhQgmLTLjCVJRDV6qjL4/m6grN/ibC1QoBIvi0WvFOR1+lbv
HQL74YUCmNCaxDszbfzFfkVE1sPy8+eyNiKYP8J13y+6hlPi1EkNHsz6RlV7N7ywnx9x7ZXXpF2X
+hfeToFpVr9ABPkYpd/LZPJjyYhhh3gXCr2FYP0LukPntjk0JcB5dQbDxDj62fOmiiX8ooZHaktq
pG8/IeLvCM8VITkbN+MOSKkx25GIfxl/Paa8tBSMaO+BSzGtHAdz/gkVv5oh6CGLB8GwF0cAUi40
hCVOK3gDwHicPZZLfWHTPDmmrOJUvwjvyw9maqXrDme4fq/DVBYwpnqeLmkWuyDC8m64cOHWsRBf
sqkn6UUd4/N2EXc6Lau6ExBGy1ZhDlHo+kJlgxCSDJVGrCtd15bkP8ADdEF/pf6OIzajyW9T+ODs
M9PEpKdSiawCKJb/MIZuK7/28Te/zAFO1fVLUemRzaIga2QL37H+nZlgPDjklWHgdX/jfYybr9Y4
yqV9tBspVEhDxcwSjhpz97tiiOJwO3nkCeGD/zCbksvNCqt2X+kOn8ejpAKYP/mDcSEE7+wRzoOB
sGfWvt4R8Aceuqy1esnQzmvqEjQJfiaTJ83vHbaMN6VYF02Da7Naz3jeFcXWoI0Un0AQC4nsawS1
YoQ90N0/dhyGlQxbWa/psLWDtiDT9So9WBzwrhy8wKz9yAT24K/2qmvKUDAEnGfsrayu8c6XGlPQ
Ehsy9aZbuRIKW/2ZnnJ1+E8VIiD8pUG6ty9HW3J9RsxSBCBfCQlm/qDxqSTp0IjWCp7Fjku+wqUE
y9vLLJeqk1W+DpinmFDpTzUa4vV+Yzgp44sA8UKoFlKj/Dhu41s2Jm0Mn9YT05t2F4ldzRnSisZ5
/H+GkFBf4j0eHxz1r0AJkNjOiBDlZDlCRvqAW6+RgrmIZf3IgkE3vyyyrCp6HwAvrUwamKLLnEzD
F69wj4SzqkZFDiCcoDE8qgcpr6e6wtCtt+qu4+HDIHImUFUJ8oS0uFy7nnlSJOy+tsNmdT1TVxhM
LO62JDzHFNGTHXc9TVQYpxlqXLauFMZtMb6iMXT+enVAQT4AhyQLNAZHgSD0bL1Bhu5qPMWvkwJ2
wj/yI2T4hjmzQDPpvOYU/kl6/NhtftMbLZfDetPWsXacxwC7YcXfKR9r+/aFcojU6CQgvBcQuSk4
dQY7AYQUzdVhs+Tp54mXzyZhZn2w9R/E0F2+vYjuFouQZuEpQFe2lz/SwRE8BdAK9gFYEKT/C7Bv
gnxQk08Gfor1t2jH7YJoOSYbTOHaeRss2jGXUd/UvpufNZ/s3gzSZMhScCZOthToZbGEhIWGMhUH
C0eKo8lYJh9lPTARmWbcVMVCfH/dXyq0KxKPNmJwYFJXh6B0a5vLpFjk7H4FYe97YwjVLRjvmCsx
SYZtBSviZIplx2CkeZri/Na2o0Jb3ztnsZCrXhV4WQyChH7Buu7PTbvKNpd2i9j37Qe4jodaIxHr
jh5/GzF6L5Y0Ew+v0Q4wjenvMYfXTNEw1sEmDq7C3bFStOrDbNG5W1DobO7Ax+4piJpC1xxbGK20
rugPnbeIi/oCwJmIV8x8OSUqBIFQrh3IRDpqSnzesWdHjjKLPn5sQ86OALJ0gkwnIA9dQqjOu3XK
rvM68DARl5TvhAD1fmQgpPyyd8o4R6F4DHhNuBHHDBl2kzxY8jOcCDXuF9tDfT+BM06jUDOtU2X4
pnHFBBskjw2aKwewO3vJSWrwI7K73dcJkZICc23Dbl5XOZi3RRPWIoheY7a0mKTPK/7yb03LgDNo
f3z5U1QqkjQqi6RZ8onNlK2lw52B5Q88yuGMn0vgD3OMH1SCk8cJZYlcCGZrsaAwp9y+we18cBhn
vlPcl6JRq3vcx5vORqij/Z79vIKyIuj5lBmldwg8TW0nUMkplJcN4dMHZX9nHt/DFSVGkyQxFtQ/
ruWyKSwHhQ4Xun4kSZHnbqIr8CMeOtR2l4vhrPSKg4cLZ9NrhUh8W7AJBsm/onDVLoTR1i5tFfQe
jJJt5XktoTQ2RIwSq1lG4QRm+1NdUAOC1ne0y8s48qY/Y1JPe/T69LPUuyYREq5E6rBUvEbIGjI2
cf5hOv/3QlaZDaSzzCidSLZ0SrtlytqIl1pFsAJuHmt26yxeUblLtKJ2YHj8GJPEwYY9KbhpLl6s
S9ATN8cDMh53cZ3zC565UJSY241u4CWgqVjSGFfqNr2DiAhBBsyuSV8DDZR5kV8u8dAeNTu8yvga
79uCUp8WE3CVaL7JpIv/HXwSdUSbZKw/KHTqZCJQku7Hf7kXukeOES1VWNKzBLK1nfbDJjTlnqj4
6rQ+hBKyiul5rIIdokCj1oiUp5otKDrDjJO5oHaSluVXWc65YOm275JAppD58q+SHVQiLV14KUyP
Cns+xXNdgkvWoQ+p+Sza523oTLNt2xplXJqPtCj2CxRAOkgBujYYxoxAqEiCAoTryMiTuaUZL6u8
+Zf560MSwi441stD/l8N7vtHxH0ZFjaMNaISGv4kqbVZFpeb0OvRiA5237wdL4cvZhPIhItAbKmI
wRq6xHsvFShOU84c2HQGdvVDnwTh71t4xJiWfLR6jhV1dTFvc7GvZIMYCSDe0GHovx+q8q5r2ljh
o4/jc4K/yj0jbQNohrRFncLBesaPOtWOioyxxm0sauvrY5hPd15gt6gZLBz7d1H03T8Nb+UL/+8V
8I8mFXWjt1rANaU+TULbcWhbNfD1bcKsqiuEjVJMznYG9qeHRW2wF2Fv43EdIUWkUgvTyt9F77LZ
pDzGCXez1COdMZ2yz23bH7suwa51MnD1qhK9KeDnpVqYgvoZ+NM+0cj6tw+YclwcN6SW7WjZWOr0
W57J8B8xoJT3wXJVGEgyX9BqaQKsQ5XnWO69Tw0pbb8Pf8y3eIUEDr98XeDgh3z8rO89baHMMSVW
TMW4RszziTesLwQNoMnOMrDuQcnHi5CzPsgfV0HJbHlAmGvNqpu4D671pYiQp81eHOsvhe8DRZ+t
zPQqHSWP64eHaWE3A7Q8p27MuIUmGM7D+yxooCeq5DNrGdC+Cvc8g/x45QFEl3B+D7zTOD2+zOlc
Zd/QFJ0Im4xfeihVFajrcOyiRD4GhgU4hokoIq+LEksA2MHApOirGaIIUut1pfZuIAiX7ZxelzXK
AwMCUu3UB/mo1Z8k7vDIXrI3pz/VUUWFJ01X9sh3l5fm4elhrTfA7XgPGmOg0GPqro8ALyjIdmjT
ItfwnnycVhmplsRsKQw/uZFgy9LgDSw3cz00GtFj2NUN1KsXiz54CP7vwC0+T2hZtkTqdITmBySF
LVUtnuGqJK/rrcsryn1smL9kgRMTCRY64E4a1rCGftVcsSh5ExG+7jtsenmZf3fgo3bObCAu3625
M8njg1rNZx92/vPUZWBeg2E5IPWGY3IOtHrVznB7nD4h2TpXgbN0rzak9YxvagOb35gJa9CJ7c8u
X8sOnREX9AkZ6sfe+pmaxP00RPytcWpYW+Db5i0IadTr6oBbALcOiwKLzuOsmL5GFyy4uBJM3iQD
WKQvWc7bHGFaQqlIyRVc5DeA0aMQZFuyuZAx/FBR+v8t5tt9Sg0t0CuMO2m/N/zT4X9AHZcmyb0V
SO1bql70A+Uf9pvWXZuQkdg+wLo/egek1iJiqD/eq4XI5fh5WquPKz5cbSy4y+iotMyBxtEqYZdO
MwumH+KHBJj6/XHk6Bjzu5YOtCybV75+fEWZKgiqvy1dHWJ9QQ1KUHLZ0RM+3hfo9IdxvV3DvO1n
93DYn/TID+eqs0ODj//RkPquxBG8lr9AYHtMXlHA0ATUwzxAdv1EAlWOIZ6GurwGoKJNpejvqmbe
jdrvhspNmqhbkolY/HF8sVbs3m/+mfavwCOedHW2ZxEQHEZr36iaSEc2ZJ8Vcg8xickbWeW8qFbx
E+FH09wuU8nw//iNisdzgXsUsBDgCIxA99p3njMOUlxDQHSawMxY7GvlLS5kJI3D4Qx8OV4LNVfb
Rxezg2IL7wkU8SK7WzsYCbazzj7JUMT6yXUDIQkX/EV8MQL746YPX/yz9/9tmjROUK71394lUIxK
GWAmqvn6dK38rbRpmzVpfiszSsZxnCAb5osuWluPz3TzNPB9sN2WSC6npYjsjWZJ8ciIzX4S4mBP
VfFiS20duMsackohMhZNvKgyYa4sV0IjNfeB6oae/vdZHlK9zAhFstM+9NWnZCCfAy7jpQavB12I
7lvp81x1Cf9U67cYzqLDNcZMacLCiese9nPfLaxwp8kQPkWFexH+NYKKipt58KZrw9KGRw9Pk0aQ
Zt6M0FbbKvTrcTClLz5Yf6Lt9fX5d+T+MJbnHU4FtNACIDHud9gcMonnkBzzeXZpFYrHLYbGZmUu
rHpPKBNG0Jr7CUavqm6UUknA1tIBhzCOFOMhiK5kJAISdWh1vvdC/dk7/Bto/Kmfo5AlaTnN6GfL
baVV2JBFnuUfWh3aInezPx3WvnU7A2KjG+7c6hcMiVDFs3yDqWIPq1bA4KGOW49ktP6NGSj9Phh2
FgNK+3W9/odk78ND1498hRXTQ5rMp5JrzCpLPjb8k4f9Jj1/9bQCawYAuhFgU7Got3/cpiShdATz
ZherUHnm3ic4A4RECSeOLHyPkxafFtVrMpGwm83T+15R2fVM+5++Yk0qHKA48yTb2SP1OTMHaIP/
xzURjPwyPgMzcuWsq+FxTUOESvfyb/7hMbBbEEHgnmYvS5UY0g9en+vsz+8dNra4JD1fwR3v7AGZ
qTYylSwnxnN9d6XK6mr6f+D/TR66lyDRChAV91HpVnpUrn6d8KxnygO4B62ZwjIrLvUv+eIgv/d6
zpU3FJyz6+IR+colncumYKVfQaNxJ/a4DMWu23b2m+v8R7FPyNliSpKfcOX/mDAF0YIh3R5HvmfY
s/ouUJ/YJ3W2B/UYoaPDZnbHKlsfDUnIFBZJtUXv3uHTVdQ6q8D5W13rahGP2btChFeEAqaIslxf
vs5A9ep/GFZShnylVSPHvAh19h65fa29aZBM8+V2SZ07bJ2O04n4g7Lpotk++/jUSjgpIYexGTfO
X243lCT9C2sI2dj+LyarTvFbYxeH1I59+n/5fGV0co47PxJjPNOQHhoDxDVLMEdU5OjS3Tm5yf0F
F4RkVxO7Ko1/rH0oYn2SZ1+4zkCR0cpIcpsEUrv1+R53j+0rQWEccLf2JA3ePWPsSrVxfySVyahm
i7/Li3Yu0SXc01xkZCS1ddvbq2DIJu2RhaC6jYhZehfLWhpJfBn1uiBlFUx5ru7hwNlSFul0Qra0
URlM22PEB6l3cY4fQ0W4ulVHVcSwhoTbBXoDgqgsYuJnBRBomOphiR2MqvOZhqmgdZ5vLC83Pwux
AfitaRfl9Bs+uI6moPzW3Xh88aZ8OD/t+rKRTZZ+ADWPMEfOqA3I3dwKKawXfz5D0uhyn7k2iIru
mypihmacdKRJy4ZV2c0YUBVytevsCLmWHRQ0g8eZCt5ODteT9dnGu49YffDIeE1jVIaQqTO1rPTu
JoV6HFOMx6OqxhdBX2miqfiELRLHipZPZr51UYVQKV9cU4e0DqYjW+KyW21EIgpsENgjigVqug5d
QKqNQim3xk5emjJpe0DB23kr04gRgYNNNvOcPzW4zV29coy4icSqvEukagj+3POHGJfaMA7Yi6GZ
R7RHG8fDhVprdDTggsccIdzlLdfwVkVczNeMqpQfPyAlQ0/LCwLhzW/lDZ8lm1JkT8F9MSpP7f50
N/E7aTIossphVuiDre+u4Zm0r9oCzEvHM4EXxSrStWmSQaAotfFbifhkKSzaF2NJHdTexrjMNO9v
Zi6gJGiVcVsC+cao4Qle9mCuvX4CiyMtVrw3FoKTe+7wvxemreSy/j3EghhzSLWe/42R07DrANOX
/e53O+RGFO4vGu4Mz1WJ96fbYGTwVFUzynsRV25HBjBtXyf19ZIJ39VwfvgDYun3kt+oa9U+Pc42
l/OxeIXlqNZ7P0WSLxULnakGntdgm9+bXLycNRb1JOGrK9Ytd6vqB+oEJK4wSFwB2S3CxDI2uH/I
rXHpqy2vZxCiTzwPt7YJra90+px5W3QE7RHaFvUw0VuzCxaz9E8aFCk535rIbIzZdHq2IvkM7PoE
w2drLUtfN5FpAoS0owvV/trVl9wrRfc5xHpQaAeVWCBWHQECZGBQ4hPvtx4h4k0iMch061bnrgs9
tZ+ZadJUgJIuSGk5gcP9O9clWc5sGLVqEtVmiUY/cf87bT2ro4HQ4nt5SSdJ15TCt6AsZbXGJg0D
DDc4lgXhHVZF+Cs08uOkhv75IhuxePVpmhrPOA0Wl/tZmhUgznbegKATFIXhC0SN+WNKS0fefqZe
0CAPXRxJ0TTCCn2JW2Cuo20QIn3Pix4e7BSrkNwjDGy+CzXHD1KkNTaX2lJaV2vPohlWfnBHKAVy
1A2p8MEPSBhG3cc5kUN3Uu6KkG2R9Vc4IGptfuIRpYEUJS5KipvyM4p8qB1EUVUJ0FfJfPwrS/ag
hORpxWTuBdEkfG5fhOP3cvpC8hfemnBFw595zyxhKtJWgx0aCnwMdhOC+/pA2TE6WkoWVh+e9VYc
PPHxHy62hvFzBrbnlkNEr3+6YBQz6mZi6CP/KpEUICdGFlSajsFkGMYFriUVjIgYEvrN7uKRf7lU
Fp0i+sTBUL/Vw68NkOY+oapCO6zC09ufQKGzswXN7NizRRTHCRX4uNW5SrL3BHW7uLhYuJs+uS4W
9ecIcCjBevJjPQhl7ZOC3vlwlMKA6LwFjeLnm06szs5yTl6nDev/m6l6ifGLAWa34HcaYhnvHSnq
+ufrSdrIQpzB0AR0wbQ2k8MxRbuXseXI+cSBR1DTdGNOkIBrn84M+vhQb+hQwexlqFxfbdNl3rQD
4hyG+CZUAbf82LttvvaXJTwTVbYNFpCu7k4I01BymLpsaJ4Zz6NxUOLRdvgXIDhRBSvaPuzMN6UU
bCwjgu/BY6fPNZvVfKX3njwDzwA8nYKkeS7ojpeDELd0f2uc560w2fRzFDrFM91UiTtVW3mfMM1X
RBgB2XR7jS/SQF0yKgBtL+AcTte7f9GhO0T9OV3O1ijAy9hf8J1NWJk45yPRLmEp7bDRr99Hci+h
BgWShAUIKTTz+n3OF5lplLyOknGnnpjXWaBcrnK/5m/kc3rQW/kyX/RizKXmr6JQ4lt6YraS4BcX
M26ocHJM7scB0UKY5MVp9U++tqhnHfNxzNd/5kKs0K9wXimnXcHIZ05wazv0uH5rRW7JwGAJiDPG
qwfTs1dScgpQ2qeaMzQx/vrd/bR9JCn0UCsN50/7IB61HH4VkpGcQiIkSXlq+9TxAOL8Ct7u9avA
7QAkCeX9EnQb1SAmf66QKArKpEdc+d+TlyBN3D4FezrnaYZ3qGT5xHItwJ2tS/i0yAf9Lp9rqNXJ
4lA1Xhuzm/MS3Bp+KdTSezTwws0tHnLhObCXzMsYHhI2wpCsX8bZxAMsUeQUnQ7zI3oCPoYcFMmN
VXhXlVOjoZRKe+F1XTRL4V/nZyujIQklP0RyhXk9GrnAPQf30Q7CEMOtJSxv5BNPwWtUKdtUWpJ3
dk3ie+vlTpoaLkEcqGcTWzI5cCX3RUqXHPfe8jEDRYL5hj4hHg8ndbU3ijEj32QwSEl0ThWwueKI
XN2pfg/aQkrnCwu1Y7ySorcyzYaPL/KCOE6avkFoNj7kQAqgu/cGXoIPO59zmdK64dDDXe5uiyVv
Y6OLLazD+o45yEQDATKZlOQhtpXk7+fjfrEraYT0FaDFj/FfC9dplX2UtodGV5jxgc0OMffftaM0
f7CrleBp3A3pu6rsErc6po3XGRQ7hof69GcCsRzoX9SvEXQ/A3E1yL3/SsJJxK4e82YrqRqIobWb
q+vNsQ0243j3ympjLUFyBMqnR6dILY3OQ0yMMvjh0zYXWomdVMVMnIEhmw5eNsY5Jq97JtLx2ZcP
I3MLo6oCQMcv8TX3iVUBpqZFe5y0/vWq1/PcoQVwJjkuO89vPHiV2CTG1N7vbSf3dVTpXbsDE1ln
SeZKyBx8FOyrpTCLqicLITwQHnvcvS8Y4RnoqDEQLG66ZSmYlBM2cHDxGyVj525txoFg/59/hiKQ
EZOnXn1b+yQ/0qTuzCVJ8OXV7DZWTIahCLky8yuNYOsl0ZOOBuRp2Of26/Sg8EkVEIuMUTWcsRe5
9FP3RDkitXd2JoyKJtOt3z1EWEq1FIRpDbR59/NMl4G3/6c0FH+IPO21KJ0E5x/EGL+O2kaVu1NE
Z6dyHbKHTOMlwXWHVdQk7uftKxOuRB+kDJSZ5UZRYDKbK/aQNxWocbmCXATX0kCzxRDNHFNXdzC9
DIO5hR0eNY0sQzfECXZ1slyxhyvLbk//HhrzODlS/UapxnublPJh/psWRHAWfPM4RIYGEK227Alt
m3AsVs9BM3yHzzgoArRiulCVsEiGSdprLSQxr09vg3zGk9+jWLBe5O9FZrFvFyKWU70c0uaaBMz/
kxnNX69xv2xO23wqjZ5RwFxzOFNXSxdWBsGO1a2KU5TyYcExMZSIvmSfFjXXtFxXczDltN6Y3l4s
h1OVOe8PP1I0FG3T555uehQq837oJg5PfLMEOeCv45IEzf7PxvLfePoqtqVcnmaFLh6m64lUSKk5
ePVPk/dZcSNZJESSIU7z+KQ1VSrAlsbMKF89nrvZYMcHvzjOEfIOTALG8/MCOj4Lm3eTRsuUODdL
/gGa5Yu2bFL2+DrRw9uWYpt6PZCaSeLgQeokBTWDFhFb6XrNFiy6XaFM7oNxMs2V9vfsGQZbzyec
VlBVKTsTij3cutZQUItf0Nx7VX2z92javva0NTt4IFwFXKH/Qb9eCXJlQC93Ob359wev6rxrnrBU
nDWVunIEIJiLmBCvtIql8HlVaDB042wcxlM3+Rv38UUZHjHdUCZfaC4/XuI6+Sfm6+hWpIzWqjH0
3uU84ojBRa1e9vHEGNHsuDiQzPNTe08wR9ixNURZTqzeZqfUQdHfazbLceMKhII78KvFdAzM5MX4
0SaqTAh1OjbjhMrccilyTovSgFAvutqMmYwHHewCfq2zYrs0VHmSzCnOiENWXsesJprueJ02PT/R
mVwAEWm6odKzvxhyyGyt91/O/0xx7hBzrJ5a2z9f7fT05n9B6xN1Ak0/iTEHRb2imy4AAa4otGYY
fDINoGnk4csumPM0eDs4pHtvrTUQDR9BjXkGwRmn7Uzka0X+k6wHeLgt7aL+RtHbmIOYVxi2SZr7
my/AtYXPNxytwtZGMpFEW35/Wvc+P07NRsc8XjxPrpGTF5wT8yCWbmq7L5vlkMizVzIU8BJEO8Ei
Cswo8lFE+yVeCgdVYr4hpRnFhXOYSaWI3LhwXL6qy1piyDYuwGPHOdU7IdsWz/U/OnL0HQgChiM6
kZTH18QRPyvT5rwhD+KQbjFt/xgbh35odoC3KyUdeovCCbSUTBi3O7gfuYEqZeEI6KI4fcxID8sn
dhKJeq9z+KPSJzcZBG9E3HMr4he85gC43gNuGS1/vrShQvgpJIg2KjFGTrtftTZdSonBh+82JsqJ
WN/Grtd8mvM1np52XIp/owa3Xn0ZBaseYEupIC1Bk9d1htYkQC8mOCbaR2CQ0Ffkh6uZG4mglQjg
k0hfllVaavU16qNKyKqUCJc+AepEsgydgnGNmY+XXVr1sRDzfew7cYd/AEc2vK1uFPbuL1vLvd3q
lzD3c2NvO1ltaemNBnSlX0Qa/zCam+nTl/fR07u5rm1YDqYJ4qfl+qtPiE+Pb+JKwWV6fURDjCAN
WwL5yx/4Q2sYKY/H4WWvyhdeShiYfWCqYDwnobt9qkRzIKgJ9meL8NM92lAIygKC+j4XtlrEXO4D
yEuhzWeMA9Y91kaG4aKp8ZeKB0FSqom/dWCej4BD4obKYNv1UG099o/USpEHiiNE4Ksg3FuaR93S
OJpF+PuQtbElztWXaj3Jd8dn94gkf5sxsU2dzlds0tEkG0OXiuzzYhc8OzNyKNkkw3b5qXh5mNgI
gcAJsfvkasllKdEFBNXRs5DRlNVAFuAukfLN7cWuhS7GfiGzHodIvmWJrrqtY9W0vB/H15a2TgVO
YZ995R43+eFU9e2iFEdYyzs62/u/7peGlSqZaKog2nEOeiTggPyhZkGAsNPVQ6OSIEQx5dvwSMYa
wTjysipVX6BF5SGXu8oWaqvyOqUr3QyGsJW2zrl+9Z22oWS+7KHcDuZETUFiFynax0GSo4dcqW0H
CdPmJnJO8swsctAI+wq5JddefoOHWLb6saIAIx2tRvPEFwheKjrc8hAAD0KzQATTm2unUboIEW1x
breVEMH3oSpbE45OJGzpT/YwBCO3mt3rM2SN96Hooee5Ppfcu5JQYZ1O8sPYTvbG16X0IKuerMpw
EIIGlfTSAr3hoXCX/JObxVz2XAn4DSDYtPkxA/NIoJ1RdYBVYzxmste8gLii1I1YqeWdNSV8mMC/
ycgAN/Qm8Ph0ekcXkMYSxKscB/3EvOc4w7IcR528dj0oAACpogOi3DGy+ttEMSQ+kUXjOpMSYx1T
oZzfdJ5LWNDVmEah5fKaWaHS8pKmShYHE8Ef+BO/So3oIBkNzCZrZIbJdlnrbSqmiPe+7Pz8wt3J
taidcwyaW136L+TlbM7uaI+sTePWHoc1lTF+CEE12p8MJ4HGBKLbmTkLFWJ+JWgstj2C0ezcwWLY
KXYdqFa96gBvMy2RWOwvssRBJOOSBX/YHq+e0r36RrjAwaIui+O3nSvKbrZ4mxrDawFskBLYZHkh
55hiQL9EtiNAj3YaSa3Mv83YFIVSs+Bq/eDhAvmeccGXSJMPOJATCMQWHpsDXZ9U2NU758dNfTaG
s/BE0TlXp1e1w8seTCjVpwQMofyZmaWVRz26Kzsx3C0ziNWgjiUslhtK33PLYctWa51zTDd1xs09
XoPTSF051vlse0IsQ+FQf2YUI7qtjFjo1P2XUBxmacvSIWD6ceUWxXoWNsbgLs/EOUePS/Xz0wnW
x/jrtiwOAzLwLolU/9RqVxvaYyqIxSBIzd6df4H6eitd2RjDetMzEk/xA09QKT+hlw2rhHBf/c14
aFtDmp9JphG6VQyekHRvSfW5rmFHqc5hcy0NySpOH/pM9RaNMPoJD5VqE35nuNUmvy5j/jiA/Bmf
bAFW6HM9q7XXjrtxzdiMg/haTYb2NEtVSCag838BA7xOqqPuBs2IQu7F/XcF1vNY8utDQrWWxbTt
6FSgwXIvA5YBiyE7jRScBEcFdHBf/sqaw4o28enxw89orq5wQYPSb8KvwPoDtlsoveH1q+WiU3cg
U8ib4F3KhPTuQ3orBena0tCMS2wrwhDx/ZVaWgsocxsCGKeUUPWEfItbvYC/19IXqrZOQB2TXlRQ
wl26E3CfFbnj0ESI101jhkN06ehyY1uKt3VdHMFGCY6rucMgpEj0ogwIo8BEVarnUdEgbYo+infe
MWYXdW7mAlXA/i+KkbEpF4lBbR4pkE0386sbnt5aewyPR8FwKEcurxDl70SglnhYLf3BLhMiBX4x
qYfwwK2MNCXldHGSTDg9xMEfB/kdbyH8WQ+qnUAfXXJcTlDYRQM4+wTSRv9I5mwlwMjoFZCHxES0
Alz0bxC1d/rQ8kYxYGKQ6daGqQBH8CwaHTUvBR5MDduNmYMYfjWfgE9Ay8l3K0Zn/v0/u62+OlHT
vqSYXeK+5WKvxuDl+Px9DroC2SSNEXsU+9y62GyvwWrs6qehLDOzpF8clAvSYEMoDVgmh1ismqwV
ScwnwxfF1bM2hPUlO7i7D5qh4Tv4UENcXLOtn01YNIzXfhnYAZ3lwvtCoYGKkK/y5wS5jmgFtFY6
xrUmYHgeNelk2+E53aicySKuhU2MwSgwI9f4H2nXLDAFrp4Erj4bhIEvaZwCbuQeBUwoV1GYTv8r
eliUu2ePCzjqVZHRR8I7u6oAjfhBrvYXHWelfmkmZhOsKB6l0NUniEOPxcOTBs0p1ywhV9GObCD1
C/CO6ubYFHIXMqPTy5etD9AV4jMNc+IO9R3lYNMXrzcKjRrOxL4/uwhXix8MzZ5WWotmYbRiDcz/
i/wWXoJKwFvBzMhIeB7xEstdIHWDwz9vYXjw4ocwwip31Dhuay5Cad3jcM8CkgrrMF5SG44JKYrs
eE2MBL0C7/123YGEw3Xqg41cZQOsjecxHlZ/AsrscdjjsdYpm21GoFJoaevOKwFarMAFrOuf0uuD
AYuQuNToHznFqGd02LbWQHKUlgj+wQ83Jad4L28aUPuN1q3ylXGE2IDxkSHfzsd2KHFkq8R8PyhF
/Wl1VmgVe4b6dNRTH8lsUQzEqferRINV40XnzZ8+maBbzoV54lH9C5cQASCooAOrACbDe6VYiM+F
+38PcbhmsPG3I0IQ6Dz4f2Soxgtbs9NNGF94pfrByGMqs2jKnmisj7AbdFH05DVbpnjKBRni0TWX
76L2OcjcbsGlOukGRxDqHOONzyHX7zEWRnTJUH9A/oYg/5jBZxKjOKU1lO1hdCqinda+jaKjOOlO
H2PK0Vl704IVpo/kDEXRhMpksBXFTZtsFbWBrmXmCdk3OwVpRDxOiTrqe6gN9EtNPjENlw57rlrN
hf3YFPhFzTD+Q9cCm7iu/Y4RmSBjjSWPqWrK617jRoFS0I+JHqCpFqnVtEkpLeqDb69yvS3iMuGG
TO4jNJdshJWdJ28NzHytR3jPSHcnvsbWoIthuyJdqZ2jRUHpZAF3rvDH+acxcrnt8qo/ysHXgLb+
9lvljw0L8ar5KphojGMFUna6oVVFxrPIq91FVUqEs6/3EOYiPcnhm+CvKr1aScUqBp+zJrJ8BShZ
+Stf6d1pr0+Z0g8czwjsUAiq2aq2bThVbC9TmsSVXMtl8/p05xPpfnLerWb297bKjUjFizZHwQl/
qTxKCwXau14v6+VIxNXH2br/Fvm7zOidfRBV041xP8SjCUf7pmpppunGjKMu5HmxMy5pUE32hSTX
C2HmnUT1fXHuMUiYERf2Q/5N+GpAUyyaKFzDg0B+vVNRPOaYmFg7WrnZjE03AnkH/oAPR/pvkVA0
eAJQCOmBiJwzBHSZbBg0Id3O7DkBnrZz0J/CSsqPbwVkqIDn/lNoi+SofOpkHmFLnTJS5w0MtsVh
D+sj13DyvSAHdeWKtgQlOwMUWOBwmwC4wHAXrkZ5a8bHdocxKcds0jIKGP9DYNjNedBESQfMmlGi
FGBbVBuevBJ6AkeZtHlMgn+fJsyhrYUTAO67/HNVGtWWrpvoeJUlkhE20vTmfyz9DvC+kyIh2Z5o
pK/fjAvAklvMIrkoVZUUtJbiQkB83TomEqzxG/X9a/fDkxvlDFq6rnZVZKmBx2LlKyoWmFfNi2Mn
41S3CXnZtbaFqnpmBJL4LwB2eyz6XkT5k88P7Jx6D5ok69U5a1ImvD6B+NMMufYMR79LDscxhl1M
P7YR3DxObqTc8Fi7En6PUiXmkHKGxDRIWOk1expEcGdCewLo9e4os24g2wf0XylMO3z30W0E3yJQ
1T/Jx7Ts2d1k1WWSDmkXlXt1z1nmDBp+QEXJNnPBsVjd+r2BjCzsgs/vUpkEMsM+BhcOgUBX5mrY
CKzlEWZR+FjqY455mWfUcHmjeMgEcT75Q+cniFRwZ+B18AO8EHy3Ym7VOp/4D2duqCax48FYQpCQ
y+nZ0jBeDssvvEZsC7/58EThWiqZRzo3g4I/QM/5c3OmzW04Ozm1NHHq5+FSkYOi2AQp3ygeGH2D
fzTj39/kTT81GlZlMAb2AJadFbX3VSV+ZA/o0L1uX0/pxgF01zQ3yWRoasBrKIh8Lq0uu/UGtOZ2
0vDnknj1GLOzLjiaDkWx3nQYGnLQ7THMdTZRz0a11jwPnQE9o/N7NE7FkkIDbctCU4YLRpV8Jg9p
Yv2g5hX8S6xqSewGZD6NGarpC/p1JhWRKmEGjsOJ0KuOeT0tHGaEAoW66X2HUlcOqlDRZHfSZddS
0vR5Q4zLvdjpZ0Aaj/nZbGCzFDk/6Ck9gq3wfCYEAvArOkh770ZUAUTud1gbUy2bYtGs/zOhnbpR
eaNg78LBTfljxuE7hVM7YXAssD9rPdjy5QitMRRqQbNiKETKw1vXg8Ry85Z4pH0Gij7uzGvIZOYn
kmMBl9RknDiHzg4OeEoPlYtt/hm8HHnPNdhXlXBQa1O0Fk+b0TskMbLek9wZqGPbwgjaX9WqG0kI
X75MjWGXCFL+3y30rigTRmAtyRzAqF581Z4pLNOUPHhpBOb22XS8qkm3vI/Tra40wGz8jScLEFfB
npDBWNIWBcX8wStWMKiKth/bE7encSJfGf3gem8ThyseMJOHWApt6DcedvNAbMES+kB15LzUJao7
VCwiz+ahtEHUVM6ktFUePF1KVL0vg1bR/2lPzBgngtkKCcbfFtCUMXRuDdO0ujZz38znT59zJW6J
Rfb/OfVNMh6M6LjxClWmvelbWx7NAzqM19MERyDX/3GFkL24vj7FkIdzMSESsz/YUP99xvtcT0x6
kYiTYCrRoNN+qKFvgxQfqFXxnhFthI1vho5lbMV4ZGidAOgk4uxn0DaRu1Kbk1fl1dbVySRCpSMU
fDlzdeGosmesswHX2c/o3ER0sJVmUCVn/EX2ob5tlHhumOhgFw1DU1E9wonsQkSj56OjQC4sTMRf
8xPhXSjQnB76YaSQIfvQr9fHfM/XvOkWA+ykFEfm5Re1ky+sCjfdShofnYKrXKv6zwc4hiGxI08m
jffR2JvaQfMjac3gedo8ru8tYiGcwjugG6qBljk32/dEi0cZjvBiZpd3BJPs/K8eqFVCteg0QhRQ
38c8sioE9uZytTeUFOHOeg1vpGPh8otiKgQKP1SV19pZhzkDsgtctq/rZkeVId1IP3f9+4Goyro5
CC/TJpslQ4pQgUbQuVUWMK45ampthC/3DJHoKV7s2OWDut/lR1tkkxdWmwwHUM0ZOxz2dMP3J+TC
4e5SnLxnHjyeSxAev4eyZE1cZO4ZgAAOycZvkqpmnCB9tHWmD6B1F/rL/c58o3pGBAtnARUycrwV
RjHBYlT1SIu2belK0Z4BAqv8FLr59DNxtcHrOdRy+qD1gQ6LKf3ionA9lDxCRwOCQh0wxPYLto5t
n62H5NI7QvEDNVgh+gVq2kCNmvu2t9GutpaYA5r4JS2P3DH26rm5GTCJXEoflaEkcdR+hS+OXTle
CaBDVjyOHm10vWUEb3TJ9FdDDI3N1ph0xFyVleFRsRo+DtGwI97rYEg/Z0KruSyWWI5uxgJQPvT6
qCjMuNfKxD0cLprgsCl1f7CjKqMMPXL7zzFOSWa5ojkH404HrGviwl6iN41+80qam5rFG4+JboNF
a7n3gZKO6TYQqtKG3RyjMnwolEjYqlxm0IvDXrWKksDox1ZfOJYOWu9b2NdnfU7sSRR9xIlSaRHD
L7NJFz/Yof/z9baXt3AKoltFtth3DaHlkahbrkDOJRdVsPfcHk+0RggsUfr5pfbh394iK0SN0EbN
weOqiDy5Pq8koeLv6rRex0AXehIRxowaDQQvbWt7nJxYTqSsoCdLJ8YsN2OBJ3Y9SdA4aqdWSwMG
gWhGUOvLDS5maYM6rXW+NTvadLgaL1MHsVxv6v9kuX+k4SSDKGy/yO1utYPWx3sOlu2Ge57I+VYv
ycalTu2R7r1VF13iNsU4Ey9zhQm9IWNQCH0sDmdl4Sl/MyHz0bv4QxgoKRRHvYc697iN+XaH/X6K
kuKhuBBrD1oTlUuCIMipbN4sRUEAZL37PUlgkJXbs8nQzQE4Hp0+Krzb6U0QQgqFhJBLaVNd34F4
OZibqWfwBnMAZIDfyPbCAryG1AVu+EbVfMfaqsopMSDmnLrPOhHgx9V/OnM4jC27aOFem9nJB8me
LRgLTYx5xzM575Z08QxOAbf1/5ZR2ad0qSnXkizn3CSuFaEm/28tKTPKcLXMTaFwsmTLG8VrPwUy
8fds4L1VgZ8gjYdlNWUyfVrqKVZv5ncgvXX12Yo06S9HV/uWMYs3BDnQeHZIByBVN6zAjRZ+kzOV
L/5OBF9Z40ghKtBtYXGZeEeF8XV4tVrB2fmbD3vxuiENyznm6OJOt8Vm08YviX9qmXFKyN8E4yJw
+wauiuyILAOTDagU1hgoOe2Um6b3w0+328Bif6B0owm328De0Pt0yq4HwiaLSmMhLrt5EePl/puK
19Ps9V0oqkg0WzSr1+8Z4LmE+ljAy3FbdT0z9TRlAqWcnJhS72nWBiukyF/Tm0tr+ju/ZawFKyhm
S46DPs/KgN8Bhbr3Sg/rJGUD/lEur2/9KiM9B+vPtf5sTwG0D/F3qDDTfXrXINFOAuCR1NBAqjg1
6XeCAH7ffU0R7c7ZXQSpFiKqFabqhJ1qGzxcJlXTmDzrvTHVxgavkntHHmOwQ3Z/ZWYbZy9W+9MD
D8YueVy4WpCDVOywLgAURAmbdbcyZQc27z5b7KWYiIXyGvS+o6xSt+W7N3ZVZ5KRWWy9DjIhhPpg
jYVwKCa1iW1EwB0dCGI4ftaiIGeIUfU0dtDYUM0T3LDTop3JDTwjeLfmq4dtYZ9iOJkUYTTujTqj
rMYENlaWFd3wQHvXbRwWvPxWi8T5nzJLX1TLljZLYZ/pDiGnpq+BPot7Qn6rTy3A4WTmOmsE6mzH
uG/HVvNZqml6mRuJh7RiCZC+PO+oMcHWX+BcOSpNs9g8wYpLlMpdb3urnKZshcnUoIqLQD+56OX1
DXN4mcJ3HXB3AxYGjtG2mooHdcBz4Q6Aup0QLRTY10RrQLXTfKwo2Wpb1Cw7KMraVnbSm3TCrwVx
1Wz5DKjfMNZ5gRT488n5sv9ANw63yDqgngQcEk/vkYg09aTDx64m2Jq8mBjwZO5MHR8GqRFw3zpD
RTuG0PqgYDITNGDk72/edD2pG1391xZ2ukM/9JwFid2GQIRkYyBSTbcl3IIg75OmXZuCDuxzvRIj
TSQEqnR3159EsqfvUPhBhuts6lefH29agKrpHBNQkK2B39lqWSrAeBmXHbD1BGBiJ2/6QdK3sQAF
/Xalu40KdXad+h343R07oZmGBqMtsVQo2gQnUjh0bFxqMueGEv45mbQXo72z2DzB6ZFCzOGLY+B9
h4epnXL2mhcABSo9n/Bvi99lK21hUUpzadd55wqV7drRh7RZVV0bJkArkwqCmgUSyH/8sxaDImnb
uDk3pZ9sHjnR4BGGXEcjLIvCBRseJEUC273qR2mQ1sJzII4kXafGZBkMPqhEJ/W2BEA6dT6apAgg
poMJxFHQcKi2kl9LxaZtobKaDKE9+7byIZac/DJiAKzWsTOwJXG4oyeSaIyTLVakBHN6wmUPcr4E
IasGsQVmVlM4mxdDU0CWZGYnlZvlfkcJvBgywIR2EcZlRo/Y6W2gm0oUE/1SMXjlEIytKDOFMsCp
INuaRghU4vfKjbtF9J8h18eP9lvNDqMG5vJIUdoo8Tp8VjA85g6NAdPF4+ppwujeP2NDgfDtrdKM
SVCeK6jsuaZCYKTssXI/alBA2Y1jx8JyYGK261BmJgth2/CWDSWBr0ihnOJ3cNxauxnxXkxAH8GP
r6FPZ79XSkyQlfkGZHZhEu2KIYzmGpO4TqAI4mXleZDNJ1XK99kp/8WtHujHRoPuK24Pbm4JKYmj
Dld0W4MQUzjNlAnCxNgd/iivMnFMGVB1LTUzEyIij5uQhYsaOxX43qTeDnIhSC/2qNtN2LbzrTUH
iz/Xhl5R1M7VaEWXIiGlUaHJx0HrIUUmr4lxSI7Ccyi/6nG0TXmZErceqD6l+VVdzDGKmmWepRme
4/Oa7M4Ouu3sDt98TgSaZZ7AzhZEAjwNWVAoZQPOgdMVWbSSE3lu9EyI1/fG0F4scv/FAbKCtVVW
+0UHc+xIxD1FSF9FSzv8gf25ub9l/IVCFeSSajJ2P29ODrkHCtZsWkjGCyLh6xAJKFc4+Wkfkkic
cfnDKktmdKuX5vaUmlXxyYDCMOukdFdKVdmkCP2gHRZYm1Z+evIOzEeHpa7IXC8gQXeRYuxDQgsE
XTCD8A0eM6lfcx+724nadx5JkxEu0e/vsngvezeEcVQ3HBc/rIY6mlR6Hcb3hCA0hau/XNLkSroS
/knHGhKJ8/XrCRmgQAQ7cOGxczr1sxQirBb6+JsjrRX1kDgQfwkOdfSMGJyn87Z02HoqlvnMDxDq
MTxjMi0JmoNsp0iD0Nfk8TRBt7zv1GvBfYqxSD67Y1t6U9s456MRiSYuPvTQrYO9jFsYe6NWXjT6
VIiB/62rOdqrmxQToEp5HH/hEEHyxjVsx5ZQYAIXJDSp+exDZqxUpe3cCuD7+a6YFOqSKbLLzd+i
hnFkdVmx9tkO/2FtJgADA4Pf13Q5YP+XuaxtozN+JkscayhnOMf1CRer4tHj89sucOsQnNd19zXx
4YoYefQCwRr3jtjnIo8rPXzRExUXZYSD+gMgpfDRX0eWMPOg/ekgXOWwm+YxeQZm6DsH257XhIeL
V9TT2OOg/zUpFSSCxAHEhNK82Hoskw2crmLd4o8/YQLfIhUVMPdqtEfqOVFw12Tc4gIac/okdyth
lEX/0+Hm679I4QSJL8O8sU+LbnaKGn7YjvqmKqDgoKqmyaCI9vKSaBULuBmzu2W8j/gaREKrpRxl
3pF80XtmJn3k3jbpLlQI3Kho29FWlkfXTEC3XGSdzIZLqSXPGFim7iDJepgvthR7z6Wgv3/ErTkO
o5XwTnOWamb/KrTkWWWn7e++YGLc+e9v60RwX4Da8hNfOPgsespKNSj63QvkfIHX+4rXDrTDAZSJ
pz7oRLzumzP9OQff5P44xJLtpC7aPPZ7oclFMobJLbpPhoI3L03VNREd8l8/Y2dzz+2bD/DGpEIv
sq8M5Dvy4z8SpgrNcevun/UigrBcqp7E29LsMaLcXEStAk+3WDD2WowMuxpk2Qy0lJpC+Qm3xy+y
e5bs0ikwdRrndXzxfdjOmQ+10BUnNdD5ZNtR0WC+d7g0VyVAb0ftVscufiLMgXweZ/ivUs9mKLC/
FJaKU4fN2T8EPXl9PPAdaPZfpwbG+I9iKS8JikA/unno/ZixYmbYJFwFuA9LyWXrh4xM4aCYurnX
Yvs7upqra1uaL8HAdxPf53N9gUrfcnvxktjqlueILQCmCmVHYQ083NiaJc/ginLkyTNvYOIvEJmZ
U6dwPp6liqquGjIvhl6JvKEP5QGr3ZWjsZYKUrgfnKrwxnehmdCP4SzILkpCZ1Ltwrq9YBTU48z6
1rXNodDaN3q56eOYbw0X8xTJuldC0E+oUEJBtpAWaWRBHgeevu+dp/FPJ9vFHAaP8PtjedwcLIIh
b6NRglJWoc5uPGCsNyi4YELmvDedugTdzHqqM3KMg/VrSgeMYgYYFofBE0j79XIdFGBFrf+IMWug
bSe0Gj9wmTGZoNgDKxkv7j6SXCiqF37ln8Bm5rsbs3pA7vTuvVgUC8aFlIXtRCts/giR5Z3Jwm4e
o0L2ZMNStYzkWF7Vzvnsa7cmRe7agJ+6EnT82AjXoGXhoSYobYW5VN+X5qnQwFXdNaw1eJa2kG40
GU/cnxM32GHvftAqnaJjf/6CKLpicshIRycZvwquGVJWqxVRxNUj+jyaxIzFPwc0u8xXs7YbGk4x
DBqq6LEYsd3Axwp7IFbChwC7yFgOv0zUYGN6qRAtz8YquqxlWLzwK5bBBOpzEQirg8974mcFNk2u
mKpokW5dR8PY69778IkLxzpQ5Qc7/bI6XZwDKy8cD7D+rWBnJpnXszz7ZhV+HCS29+waJRkGr4XD
6dlbZLJ5zgXGCJK3vdWxATi85PQfxuK/uGj5L/b9hcwieO0r9I4BwDQrXekl0fexGe3b+95m+fFp
PmDrGnuHTO05Qtu+iMrhHb6bXP7MR7jEIvSuR1qp4YoOvnC7u9MbWbJUkfCLdS8rNt0xvZ7Fn0ZH
7coShLk+gLi/ejQpzqxVlDBxLWqHwlNZdROp0xgOz+2ilQ7f2iV1eAaYoy6QBdZTQsifj2VGWLAg
FH2xVbn3AYr4jgozewSRNSi00VniiXdPEh8d42NMmBN6dAqyfqSJRAPeloUteMDPBAMZbDSnNPxh
4ciAXwYR6p+H+DPJUlk9BfhD3GtYt1i0o1K9vA6lXKyZ6/dP+r9bwztApRFks4oN6j1Vs277XXfE
GWpyy/mYffpSp0yLTo13I1zKPafZDvq3xX4T1AeBtGroT0mUwzuUDvnQBW1w39JqdpprzSKhFOFh
CQCKY8FjFj7A9a84u1NinAsV1B/gianJLtQR3S+6dWNMd+eNvxqLRkOKupgcyMqlp6NVozins2UY
Wanc9vxpqhkvvPUc5QTpCXuuiGM8KgeTRRCek4IfdLNbT9CALmNM8PDJB4vXWXZtE+hCJGff2m07
B8jcNpO+gyK2FWp9eQwS1xT1/SispXNUIIGrhTm/tQFByw1jgJ2/McVUYFn30ShhR2kFQDDgFiuo
lEIJmRvNdrImskyFO63YnA+wQy1PuY8hWPBhLkZ1VLnQHhbHZNB9EuRRiC5FRJmQPfG61bjNRhzD
vq6BoYKQSeV8CyoeYj8praDU2vpCmRAcelEm0rxmyUJ04IjGVK8yks/PI8maNgEQpeYmhf+re83E
Yzk5m4n8Ji9g7IW7osWWCDb9LnyyabsIC1NYMTN8H226giMcbOJVFUVi7cbYQkqo6anDq73d9fcK
Y77Tx+VH9/eGuf2H29z7LiaJUeGRbD/E69aXtIbJIwJAXuphZgl5vabyfI9s9k9IXOym6/zaE2S/
/mgBy2f5qjMCHQzbVjpKtyg8g+oCR+HEMcfNNMmCGc8IeCl7wUsMDOagBBNdjfFjt3ZfUXRrBG2Q
xFHBGF/PMAyS5JxC6+bSrIUU5QAwUs53j4sYPO2PTtP4UIAqbQcrNBQMTePMw+p33O8Eg6QzxOzD
E3aIgZu1LVvO4S7JeK2WgB7H+XsOzTKXZ/Zn4lhgyg+pHjch3dFIOSDziw1QwPo0UOAiXAV18hiy
CaqGAA5I2GImh8nYi7hKEb+N6b8krE3Vx+voS2zaS+QvoYOPwHCfMo97Kw5P7O3E1pCefMPdSWS2
BaNiR6RUl2MZca8jSvZoJkm1hUueScYFT8Om5ieP6ZbCLClUeG+az40nGImCyEyVI1CJgfP3UuZ1
dvzOHDIyzybZFTv5gE7y7f+AF/GovGtRQtgeHp3Ag3e7dEcWLvoSF3ZIPO3Q5lCzdipl/AVhhrzB
R41dqtYMftuqadHoPToHHasWyp3Ql3+pvzz6XUTJwAztHERVHBv0iMPe1/T3gNBnfVRmQmQrxalf
sD5FRGgOduEyIb4NCzo+PPoQJzbDMs5u/NCz9ICZoeNhgzr2+cRTlwm5K7oOLtTTC/NG0Vd9OcDU
UdTnze8clYvfUQiN62bh5BV0inAy9p4KHauYNfXKxrjjruz/qAS4Y2VAFP95Kvh8JokzoGDTGLfG
ZzyFH8nwRFthbUgDoDIG65bOC1wO6SGKOLxvyYZ7onMsHsbnZza9pIek1rqCV9BLOQ+S29lJG+93
AzoWN8dIMrQdDykkbwE2shUiAwFAhyeG71NK+0erf44G0pRCPkG+l9Iz3ZDLWZalYiUBNGP3BSXR
EAGFDg8ph0TSJs+hPkSnaaE/u2HbawFhYuElNOD3ciGa3/EHIzMAQJRiLR9rDBsI7paV+ptEjJfR
ziAutxVZHRPLIRDiRHmX/+fqIfn1rJiZQ0VIH5B9kbJUsekfAI5b9dKmHzIBb9PFNm3oyvLjjrcy
O4GlBSX0mds0g6X9VzLwIJtd9Y+Q8dzJ2KJAYafV1BllsVDRjpJrGoSCXSpr4VUotvoOuUP5YjuQ
fUBuSeTYxPDFzVUipI2VQI4sM/g+vCJg+LhYFZMyIyPVcuHOGAjDO3akCOUDIWoPgSF1BcQvua9m
BmRQaWRKWYJxk9D4XncL6VBs2mmu3PJOss+Qh3UOvLznd4WpSZ+Xk/bneInJllwfmwUhle2ZviiO
D7oJZyZvS+/DEGzFKimMfAiI+astuhE9E/cuzkBkuH1u98V3zDFCwVvEhZ8bDz6yP2OCZ8gxifJ4
uftyzvpWECCGp3GCjeUTG2Hzgdbk2sxQ/GRfs8z9jXGfwf5BZ5VTU5S+6r8i6m6+u55HUIaVjldH
wijUBNeIGEJCuQBkC3nh0GrsCcwbURQy7dIws972CC/vkqP94oFTSYNWzZSMwSuOS2CdIOmebHb4
57xjf7JH0mo4xcF+TLJOURdcdW4G2cbKQdmVvj3laLC2mYOzFQt0JK6XIvq5ih2d2B14dBK3fhaV
7/xQXoV9zTgsA2RW9qeMBKV6psxx9341LjY3OPdVoL0zkbFSEHFVXmFXSSEnC5bm0HyGP3e9jqHo
eBiu5PDXMPYXc9vZ493Z5FJ9ZmNb1XpY0FYtKq83QfqNwU6on5NLqnSNkmSSvxLad5jcFBDDtymF
3rxzJBkzVKcpoMi56tS5yYarI8acqnDAF3ocib+3dmcs07yQCOq5L9RmLECEv+DWuP1KDqFIDsF9
JZ6VZPSi26Yp8YtUwbNWQK5n1gIu+YA84P2cVW+5r8X7aqLL+J4pFab7mD+8El0vRsWLRb2n1Fw3
j5EM+DquGo/cJdVs8Q4tJqjwIBU2PYlakEvzdc+p0Wr4MI8yM9A0Pf2uHjdWNfanxIaQW6xJjpsz
QQbzTruefeiz8aSGlowE/23AUJ8I/YXnJYYrfrcpUYk7cUncQaJNf5sF2Ps8eDnbSnfw+qTLdT96
BpuKcmhw6zTl0b88qUzSl+MolEwZ9RL+U0TQdfPRA9PeA+psqqU2K27sPzRul7sxg4/LKWKRc2O/
0u+tEsnoUq5lp8D74kzWB1Ojv0bmrGuj6t0T/m6ksWTyhCp+/SIS/wuK3HveQaoUTVKlE6a6viqD
aAFPCRBv1AYt6hfl1togO2JltwG1k0tlGMY7ccE9Zlnj4M1Rg8VF7z8abx/fQfP/OaQqk+W4ai6s
FGyS32KZPcFsqRtLL4LcyjwAwOobHugzAIm/Sb11suS8/QqMi8QccGbKL3IYWo6jm0kuXjP3tVDd
ptm85utVHauBCwAYz+JCKwVGDzZ3+lBto4XhEyUJWzO7DDjM+OqmxoKFMynnJSJDatqpaHV3fZpP
3VDn3VpStx7i6K/Ysdi/YQ3Xu1xS9Vx/lJKxz7sRNU66gs0gEpOWpBrXmL//08NNYgRuuWkoXB0h
asJlzDLoUhD0BqV8TB+jpJcGtcIwSpIn82b7Q0nu8WzX5EX7qhjSdUY4VxB5nU+AoXI0lns+KFYu
upTGCqjHUPnzC8HAK2lL8EhpVGCQDQBLeVdvTCwxqg/gA3iAPaJSgf4EvGl5r7H9V1PxUCL8Mf7c
g5b5wowBJlwuPztkVYji0VUlLHGiBBWY6CR0JARziwbdzcqh8zxz4fnO1USCDb5dAlR0Q7rlCrT0
gWhdGAwg0yLISk0XxnA7irlhUCxyFG+BZE17GwuqWuuZRL3gG+A7OzD4X+rtlS/Yv4Jx7Dyx42Mv
A4rol9Gn03lU5T/2qSnpMXAQdHFeaaNBFcwwElzJZnovAm/ABaNoBIODrF6joD5w/IGsLVOuu8fI
il6WesDPDOgV1iECwPLlhTmHupcInLEWiIerzP8FKYTOmyTXTW+SX+uWAPz+Vy8XGtgxuSHlyqdN
0rDhitiQjD16iBAj+yEGeqpAQAadIuMEVGd6NxccWBTk7+LBeFYfUxFiw9+8ZzZ16YmxUX6WCUCP
LdGc+riRtqrVeAkq+MQwWGmTlibzYKsey+1mwHdDaedLF7cE7GPylcWyp28Y+iXDxJBvecTSkeB3
Zo1Q7G+fbiKRiQLp/ZJQ8CvCM3MRriSUOZ73o+Ztw60LGsJlrzqok79MrGmnqJ5HrU8Tz7hbCUW4
3vPJyjdyq8q8kL43xIYd5g/J3bRincu7kMHS11DBkQLqvvEdnovoWbR7F9a9u/m9+sMfzTCgBfMo
8syGyIH06JN1zo8pOe7PZa8JGEBL8AH12uWUwHxFo6EMGk0LU202A4r9tFzb/6JNymoM6507rctV
cg8JXDlVGEm/XapOCoy9foTc+FKTAGFG16Ht6cB8ZUf3yjcpfyqxJ6/7/s+PC5PtZVd0m1fYAiZz
gP3XgzKjeWrdRirhf8iG7MHWz+FZK162BBeNZtfKeqLaAE3XMBMsCXkNjwTmAVf/CqfCLklH8IaE
WDIimlO8GYKjDLdq88rA9zMiHbnVn5Gwyzw3F2s42F4cTVKL6NcUVvVdiCGRdgfBUeDil9UiqhLh
KsWo9UbCFrcAD3jH8X9WGwoGBJ7Jlanc+bPhg2RuOwmGJlHHEtsJLeVXhERcp69P0k/TpMan8tzS
xMYKL4rIQWs4ZE/ejvkuc7vMjQXJRcZGgfs5xBbIV55F6Zq4KkZ/1LLrBS15v3KEbH2YHo2e3eu8
9Vv/gZoD7tdIVlLbt2vjwWuZBApKwVEUR0I9zcIuecTmbojxTjCLtAzYzmlFAcjJVe1C70LLXARQ
SoS78UnfurJWzRRKwlDtSzaqS++/lUL9HfhE38ZhdUy70Nsxu/5jcPGq4R9pU/BIx3ukWuYbEg+b
ayl0g1NaWFBHk6ZpWNfLWDv08GfYUBBy8nQi1r3mVSc+YplZZOnOn34tVUM0P1trikWsyi4HwySX
dNcyG5HDM7GqlVloDnKUnDKilNlNpy+tr3IxIHh+TtjKZHC8zSxXJPuUCFoJ/SW7dmY4KLlZzF8P
9NaxI+Ry14PddXFqMoB+M1IY/BbLMz2UzAQyzWuOAuAk630Yta4M49PXZLckPHv+j9q2dHh6pI3F
/dJFhTpeC7YXo+K0vo98Nqbs6gSj+bZG7tjKKiuMEiitVlUJTHNwHkFso2/HsD9Cnv4RtGnm0jF9
WA1EZV0UNnX98ZeMXGQaibF3AiZuBnOmlWlPqgYcU+DAtEGLrC6IQOJmLaFcUN4Jo7p/o/ruq4uS
MShhPjxw9tk+QsQo+/Jzu7rCQGNaZok2299l03XY+6mAwVq8JOkbH3AFEwFeso/mtrEq5c70BwjT
gpO6db5VXHXv4G+Y2fj56ZFPhW8hyExUxbN2+uPFrHGV5O5wMKPWnp7dI8FUM48qKEIhC4gQHJ4r
gC8gz/EdH2S5Vcur3snArSBwkrA3t0L56TtIMjP+pcvfeyCGlo5Ga6BwlJv1HgxchpJaErsanpw9
XMpNhymXZ2XPBBuhmqSookY10oZXSZvocr7qrXplwvHSAQ78zrb7c4sj82jRMFBm4jrw+rSP8Olp
nj1Y2U2tMHHxH8Mq/YR7XjEK5TJ3YKEq3jXKmIjddqMxePgcGuGQt5LdFMr+Ypn7pJ4zb8ZeRWJw
2wOrlPdsWFnUqCZMDe0X+39bATUqC6u5BCCJJ6RU36al4lgqeo3NftlA4IfwYuz36MG5ZJZfogC0
yhu7KDc8ZYI9IahISn+lQJJKKNveE1ZECcu+xfIkqWtg/6OVQDEeMFMyTeyAUoAfPklIbamzF0U4
ovdBuCKURK0A2pubGd/RZabGupuN0kc70ScYp568aXDuBINylSvAgumBxGf+9I+tr+27ZtdyyWkX
LfuuE2BDwbbctkYCfdi0I6tZDxYgI2ooFkIh4l1BNBuxfBhmmeiLF/EZ4YEmgbAgYlZJtt8Gok73
6bXf57T/zL+lJ2ykIHWyNbeIJPzk6t/qTxXvSR8TmJGZKWnvaSVZNl0YO9TU0WIND2lxDK8Eslcd
uM/jwfaon16HDKRSPIX+tHvx/BJ14/ElVl27mhCnXKsuiLiqmmy0VN61WkhEjjP0R3jhwoKOBWwz
ypPPJ6zoON8HXRE4lPIPktfjtcYp1t8faorm5s1PXRaEO4RtF4uQdsU4l+z/kefM/jrYF2BE389+
PlUriUlryl2Hk03+mzfrvkL44THa0+TeuHODFduv3uo1SOMdvjZEwoJdXO1mlGmzAY52HikYY83A
57qa01em2HWqFSOOGo07fm3ZYSE3nRWZ3UYZO87VOPtuE0HTUbVthFp40QOzfM6xGzs2FHmi9eJ9
LNW2mbM0OCPlfzDhH69VrooprGxCKfpL+9KWrRaDYCMzCIL56FYOJHTMi9pPEK2Lpoh/kDVxpfKV
KQ0L0DErSLXN2VFO7jnqQaLbzrBHT77SskMPGzs6kXQW24TxG2lDU3BnuT7ZGlVkj9GJCFBg9woE
I92FW1z+wGay6mA0llSVQdKcRswpq9QDBWnc+b0qg8LzOd/yumzUKOhb8GxqCBk0kz6+Z4jfcCch
N6YNVMb0j2qW8P9RJCw3T08uTq/RUILnFLFI6fGEvIJVSFq3igbGodOWNUDnkKNZR2/CtkwRkUxV
8GxZuuWHPrYGymdatv8IjM+9ddMbAeCWoQKq/xOT7fbeosThU0fHnI9/uP0y0lmB2K9TykFuqGx6
f2C/+nN+yYOf1FtpXFXOtvIOIAa9E9b1Pg7WZDTPwFoyEw4EegfPtR3akBl+uTJ86Z1jyE5MBap7
/SQJa577RuTg8oGAGRF0g1kNI+j3lDpxtA3ct3eTqLuxqX1VAe0yeRYUzRLW1Jux/1zfelQJ77HE
3a5z6uwNOMCAGkzYU1COT8aSgzK8UdDUGj+vihGVliw5Jt13szavSgeUc8wC7jEFdB4omfbA1iuK
WCTUlgMbP66AOA/ju7oT9vz3rDxMnknidBFJYJWjMH4Ruz1GOg1zob3HSwTky14hnbyehnTugMU6
faX/M2cRDhcP2LM3iEabHnBkdCFsDFQcKdLMto+0LpGbdYdlovlkH25A1g+uXjW+mqlb5yJohT2m
7lgJnzSgvjWOGMMQPfXlk7yItyxUSylDVVSyiEocXjM9+aEUJs9CeVWKJa5iEYwkacz0bcsKOvFl
t1aGh8f0W+CpHM92f/kTXnOig2u9VOysYi5IHDf3SuE5n2AdAJS0g+rsS7VAvZYoprNs7YHItl8F
bPrX8cyotXzFw4GBaih8fjXKEFC3qRAdYdIdyi3/ndpq/RRKrBjixYY938j398ALfPS34vKDK/lP
mjdpx7csaAuv5a2mTrqqH3a+3BmXeUd3zDgLNssa/OOCQ9GusF9+BNILpvHzsp8IYyuWyCjFQ9rc
cQQvHYgudtNzK404srMBV3Pp7xgsT82jaUTdhqS/VQnN6bTH+DaR5JQEAaaMpuOnluCe3LPD9Jrm
uq3FMCqJ3z31mD/gSrz4bNIG06qj4DvKDN95KIuYozZVAYuIC7eSCtw77Zfwon1gR5iGo+KbEWPt
P+XUsYNf1RcSVTsLKuhnfLcehUcIlFcjLADgCvEL+vf4128Oi8w9fLBZbk/cdu/agESb5CQzLg8v
398wqixPoOAeVw/AwkGGtfP7HvIQm7lSbbhjWmO/DDAwchCplfGqXxMzzVCo9Inq4WWrcRNDj/Ek
KYaSO66st/kb9OsraUsUDCqiB9mZ8ZzCwvc+ZGyYod7yoxxRQrjm9/9e/Anbj+AlCch0EQVk/6rJ
rFKbwsdWBFbdsLlyCvQj9wfJZkqmFursS8258jjE1cuovzk6/d0ATyGSmXdcKtegI0+T/qppfDIQ
dIFalq8j3Dw6CrmOAua6giP3WsC5CwaW8bdO9igl6dfZXljIB+rxIMnVDgnUeJO4+zO9EIeMM8m+
H8v6fKqk8xhh+zcxkE7k+T0wmeqVYO7swNgoahNvNWUoCK5Z8nzdk/k9ZVP5+F+XHfwRCdfWkaXg
avfOI7+82TF7GokYSvnEsGiF0C46IELXJmhrUbR3zNvAnWP0etnKOVSVIf25bsRX2nXKZlYie8yz
7a6j42COmghcjqKRAYP8zeBdOLvi/WCeplT49nHNGTkESn2e7CXwUYJ/NpnRN1SITcIbsZRyJV67
MjbEs9P9V7LPpdNf6P37tpe05+xvI/ui27qhJVGqRVDqtYfHatFptddrCkMawycHxWFOBOPPZj7k
1O4fs7Vzv2qRQFl3EvKf5S4bZJfmLnOefc96uwkOw1CQXBgG13Ztt14cIHPNf6v50Za8FUJw+6cW
ty+HOuBtB2+mgaFvkDDljLiVnqsYI0k+wT0SJzAChqMJ8Cz0QSmWpYteqJd2lzOtCYWY+noniKWS
L+A7I8US0tl7uKUA18Bt4YZcjzjVd6ZSgqLNW1/gKt5Y9qWa8sDpbP7O3MnfYY6DU7gj+imPThO/
ke9xFneq3Tz1+5/eDo79lLxy/B71wyYchC1D+OCti4AfAWUb3P+AIvIvXq1CIPRT/rfk4HFFyAQB
luAmXF6ntiOxkWfuh23vveZSp3ujKYyw65htcjEecODh1mdiVoBCTsjSB5aOaX2qafjQrj85KIm3
lY+edAqlL0cKjUn1i6Th9qOwwddq5zePZSjqeduw4S9x2HQ7RH3kSr26ZSa6yiv+RMggLEDe+3Mo
xK1tfz5mruxU5EZb49F7VVgeZMvtR0Y/68Mf06//7aV82wCWwJybfyxlYCpPf5Cjt+cd3Pg0RlGG
OdWPdfFZAgGSQu5QhJuyAOgF38wlq1qzC1YtcG+iVUP0cxfVvTK+Izm05so9ly2YPRFgU0tAeO/G
ixQsJ5ChA6Q/EVlX/jHTP6wTC4jhP5uGUvVuwB3PHqFDqV/tT5SA2PEEtu6/+WLjuOp3I2fK1Tze
QotlzMaW136GWgbRCYyDWwyshmqK4be7YzXzt1bsOmSkTNGHoz0YA01pB7PGXQ4dLYR6taEOKQXq
4cPHCd2YLIVPhb/MShSwfBqIFDLeLNL9dTrN/rZSSRhoAVLxtBATuf7IiPpcRlZMLWdWuvH9l/a9
X2nrxe6Z+GJJhRFTBHKjPu/DcTWbfv0iBd6O2tNae+WCY1cK8IRTVdzn3mVZRwahKWd8l4YaZRNP
GESJ9RYoCpmKiVvB/kjonnx+F3pWh5lg3JKDx9K1ggZXQ/G1TLBv9tR5PI0iFrH0gO5LPV/nm861
DKSN2j50ltiZwI5/oDtAyl/gyV0dWmBd3LJCQjx3GnJBkd0co6oS5HSHxTMi/ccnhKFXlQj4/omo
WbwaYolN9ocw1gUg4UzpiEeLlMTuqMViGOGzvnDN+jGZEQA8hwb/9QJ0ATZ/Kb9XdJTifupPlJex
zkd7pOZMZQna35rfeoh7Csy2T63l9b/q7Oz5lG44eJnxzhB6kpYAqcQty31PeU3f+Au9f2oqmAeK
CqPYH3D630nt+U4BQySSs9bmGFxQ67+x3+P+XDvn9MbW2TtbvyrbjP1ULePUbAEXo5mgA2GcvsWG
WWkilhTC2YpGHuePeehqdAYVs7rgYSnPjWE+3O8OD1QMUz2EiYs7obSmdTF36uySDHTm9WKkojOj
xDbuYnlFXnqQTGAMOdgdJqPuFyYKqE5SLsDQ2s4AWlu2xV/nFLlAAmX8jTHLCz24M/l2dakT1dfH
iJpMcAdT1PbkKHX8Lf6r2Mr3z8/MfB8ot/XOdMBI+IdnG0jfKioHh3H8t6EZfWKDqSQhEz9M/IGO
rcCCnZFJW4Ycy0YPHk0JmK+OckMaupmb51vD5gpEGCNTDPB4IeiwtS4/xK2ImbklvDgz96yAJ/8D
Blc/OjWkDGiNCA0AtOmnQFePRzWdwF9V16qY46Gp87pDYLUQ5plYDOzwtaxXI5gwspR96IUYOeuD
+TfTfz4WzS8wMb/SY1lAdudg/YBedYvU0F3dJNbaLfri0l2tm8gy55zTrbWGd4imiGRKUOWyMwqL
+vmfzhegeshGjQLt8vcUYegbSl8/kUqV8xvj7VEOGwIcOy/z+jThcBEk/CyjCTFVNyEgVrH9Pp31
9dPNN/GqRdQTwLw+h8O1hews+wtKxkm0PPOG/4vxkKhqEZD9V4Kg94Nv6aOJxYC6bzPGI1Iy+8E4
gjTZciLDKmRLJa3ljwY5d5txhj02WX6YUwRxDhIWF1m0oM+qOZ3k/uUPSYUFhJk2fGCgYLpH55h8
fxxAVnJVgh4bl32j0XQFDyOeXmry9dZ3bOfyr0WpQHEV03CqM7JUCefTyqsS4G1XU2BapgPd8ep3
1UXV9ZTMPgOr2xn9GYNmPCpoiwYWH7LLZNzUC8KAMa1lJSLt2dsGT97FY7VMn9mu2CXDSIuKsBig
/vL6zi5kknlQKxqmXgkmqGR+yUTYvhvKdvmC5rTgJ4fE+jAVMud8vAcuFTi+Aq0sI0cM2WCDcmoA
QhFIbZGH3TN2mYGu1bHAvrcZGgIE38hUvrBqznypkGc52D/7evAxWzkt7PrnAFimFqDFNUQ7IMpm
2E+4Jo4Jb8S8kk+QVEeeGzzupzPXOdBZlCv7G8kIdYaow6+//VU16GnAaqTzdSn+Rf3XTrXtzQIo
X27ymlWdw83NQcWe3HmApzPaEBjTaWrBz7cBgYB88p17IqNZU6EFELoHQ1If/7HKNxnzuPx+tnA0
aMjbtoarH+Zb3Dor9BEYv79V5689m48E71Csj5wsta5BFPmHn6PZ7C1XPccelGxjvb2snZSf2CTU
QPdqntngJUbetAzwxvkUtsUT9l/Y40EYKN1AHDoB0MwdKrzk4BByYxqahlM3lHBpXQ3PksdG2GL6
dVW2hDIZTF78pz96MP2KVTqC8Gt5ygRoLUhD0u/xyHCKuVafPgybVbpjR+jxY/3mVV0pvXUV/AVu
MpOinjM9eeCGySs7EzBaQTBCdusU8cOdroYE9oOmbWx0AyA5JSf56eKE3rFbi4NOMFEoxcnCpFkj
UIsEo8Dy61Wk6qFtfrw5D2qj/MIZ3In7TVp81W30ZgG9rs3WM8ZjaMX1vdd1TkcxBwLM4+RjuUqS
OSQmzVKbuM7q8ThAvO+B8SjNx/V6OI5/9r380n2+8tgJQfgrOLUXEwtPL+x36gjcasrG7adNt+7P
fO2s0IIbO5iF2GIz00GpOP1KARjLLne1Bgq8jx2JcWgdo/jbpM9kZxsjM6GXWGhAyoOkBUzyZpl8
SJ0GRZqU5gsvlaq2X9RBJdLdVvCZttm6RYdnL09QFy/UYLp3La/UBOqHLlEbn3GjR0fgrGmA9T9Q
0C85gwQgulBsndTlgNVpCg0ry/duk4Bjrj4MLMqlgT3ocH6DVLoggTFZ4RYJcaENt6z0HdEhTLoo
gw6e3GDqiAFWWaK0IwWcKtxQfvYfpFN1ckvkFX05YWCMV5VGSVguOBGqgzl872Riq7OKeNAmyHda
zAUqjio9jJ9rnIrDoHDp7zOIaFG9oRPkt4tN45smLN7mXEOKfS7PzkaapPn3iUgXvVBdJFqXi4Eb
W74pcSFSmHIin+FXUhC0IiISRuIcz2exKadM3Xk7So5jsXO1LJuWchhUl/6lJzRuKoqqBLJLVwzx
gQJRR3F6hnUgA/ra8Hn3LMz4hFDyDxwgdsoAF5xR/idypYbAiqs265KKOwXV9pO6P7dsDhbXR9Fi
Fm0UVwuXPlCRuyXJmYgAfVFOC3ojakwfKR6xPZUnyVzsulJaQCwF9W0QxLB51Xw71KV3PMWgu/h4
ZFeNBJpJvT4xwV4AzvDL28Ret43EfA+sql0veJ4fqiRcbloyN3lZVm4iDTKC+SFtMmMiYslGlk8M
epRoFl/+q2EaAuOffyKy2FGfgR08u4XCdAUtfnohoXoNDMGefVUx36LF2OQg6vWIWEb5tgXwSY8s
1DXeDn+SOGD/DH560ywZUmHmdvnbEsk3Tqy86BrfJOwCpeg8B5Cser6cfq2eMrnfNFbdtA3kSKJ3
hlQRmum1ghb0CUm2s2AJmHJRunP9hwVIPF5t9p07PLEc2ThK4BCTIVF5pKs1ZmaKmMpug7QxLwMl
3z9VMe6FMDf/IZ2HXdQs/KOc1NNp6F78bjNe41zoEP1BRAnPO0OMNdALed1f8f7VEy+l97aQmAdx
bSKLDy+/R+lG9ejJJhVgjBVI1PcXROJU7SFeQCccyPZDVRYTPRiqUxCQJA/glRShkFD7olVT6IHa
SmzLyRBS1gdql3EwhtflwYRr1JrEPXSvJ9WupFPnzcr1EFe/5uGBgfYFkOMAlAlQgEWvK+Cwd0pY
6aJG1tnH7AdQfscrLPXD82yZRXAlEV8MN0acU02rkaPLxxDAhzT8bRh+TRpoiyoOBD2BnHwK6EJX
Z1ZIAZQSmXBP/mn8omliX3+mAyiZIOZVf0wGQwYis41jzeKKgS95YqVhjUZrPYBR8w3LkmT8Zzyr
yXfxkdkN0iJstoB3U8d6FCKDL3ZFO1RsQFHD3ipDYLRW+8ULe+8ah1RsJbCuof7TyEvqJv0hnCnE
CPoYqEVToznHCnnTKYuCflSYaO/o5Wh92MqZgoiE4qfUG/LAnyfdl63Ow6HgAaPQt942UrRtas+j
Fz1PFCzj6eM7i7DGqG5rpoeIj0+FsoUO51cxpAs06xXWezRgmK8BZIJiWO++Y3I3zh51kkhZLzdq
B4B1PJA+SH7wdVSZDwR4n6RJOprFLF+jIXkpJwjswkgqz/aqqMpuEBPi4z8LUdPCmSVLg9gU5vSA
zb9lChlMJeoVmVJh9WQg+a1iTbDOy+06TP8VBraOYybChEOwqM/yH6/yawM/QbxYj2qHchmSXpyb
+cLIoyS8LIgx8dA3TPqw2+bl8e7PSS+3aJ9GfPJFre3DOFf9UNJ4y1tDxttPOOWPZV7AGfN8LSJc
Cpq/FHvJ7gueJT9PC2Qb/NOZU16v1dmb6by1Tw1MhCmlJ+WkbzIzxoaeXBFPbTbCkH8nGuQ4WExj
u6YRcjHg8wd+higQNfxSYJf4Rgxv1WPOb5TGl/ubZJZ9ERngcBuY95NJEk2HdsybHgCXM5Dn3agw
lVUg6T/EY7CPEoFmzOAJMj25M3WD0qjyrSCiwE+lkFg+CTmnV0WcocoJ8aIG71/Nz2DjeqejGvLS
Hp2ez2q/Qur+j4FMAvfBmkjWIpyW4Owqe6ufwkWwNQb7Hg2WRX6ZwrXBBjuWjPZ93epUOLwYSKwW
BZatwtVJJfcSNiNDQ3r576gZov608CVAAdLI7Oqw6p7dpW3k0WPwKKrRFq2A0jHtm4qxa4mS/OFZ
g6zOpfooMqkVjKpynXeF9ey0JGaBQ9ciKdz1aVuZxl74ThcCyogwqI07rkMeST5CaHPH1nU78bm6
7KjJkOjwJhzw78sFPiNxpRbUwh3ywHQi08/oH2v5PN4HY255rN3NZTf+Ur8nQp55vV/SwoHatIN9
cln35vOr2R8e22QJdorsZlQHb+6Ya/HcvCiR8phrbsEt1QmpYBbJOuBVuQmIQOOr2mhNSG0GO7fZ
4yQ+P6hPB0JmIuDqnSsrUnRcNmIKCXsNmpG2gIOAl7fepYMkV94H5PNM11nMI/gyh7zI9+UU95Ub
LiToi0JPs+2LpA2/KIU4Vk4/bEJ2/0C4OtzFvJK7i0AvL2VSfU4zeb5ZqtYJN50vSJoohwB5II1U
Ix1jZRI6wU1LrZyUXNbLAOvBPMAuFbTrbCaYT04OcopQx04czOeeGu+txanbo/UgSEtrINsmG15+
q1eH6zjOBRu1whELe3Vvn3K7tlmgLAzERE1RGghb12YjlwmVyKr6lph4Q/Pfvgtp8nOvkIWyabvA
GHYSBOhMM0Z9FDkyCeMnPqkhLJVnRotOoAAAkK1XxFmleWr6PfTSVdpv9sZdRexHllCXaYNrGZMq
saVwUFbevz/6CRDlzGeJ890Kj3Eh4sdSSkUpWgcEuPnEznNEA+1AL7ES0GPscRuPEEVZGsoUyn9h
tqF8rctMdbWp7UXSKDTYWSfmHz0G6H6fzoZKANttWEFZYtjLtKRvc9USTJCfrI7IePduQQKugQPL
2d3ZIzHAcRcbH5AVIhX2eomMcoFNe/oUZUoNgRdX1nCpdfOQtydSdxz+NEtOzbP1O8Q01TCfD6Q5
ngtEXSlsUo+7wRzEjNufGZ83qNNarn+bZjSPkDivS7ncprmpmj+OUOJ6hDGi446EBAhptD8I7Az0
EVIjHUGGnynsCo0q5R+4U6WQqMiAmSvz19GtFCkxuzUE0KzIcRLqu7AKFdeLRPMN8i1HfBI89RCP
/nYeGHr/weAK95dZlak3bHa9EEY0xVkiKodkVv/4+LaukSpms4Sbl4OefeOpV+p3PlwRN6pS+rHU
GNAtKyE9ywDJGe5ZjaJNjf50xMMroG3M/GT1Bio12iYv55Cxxan8d8CqzrnkpebV8gIBhZKzOjaS
nSDJ3JhIBJDGr/3w01LwGtSPIJkHUF5ZBuqwlq3MngWBpyjXDT0in/jrDVd7xU0yeZy1576sBovX
Warz3tGaHbeVFwtVu6fXwsdvvBOHUv3W/0njhKMJVacHPpk2dgD0BiJPRWW6AfxiJivzszBV6xin
Xl55ch0RM2ARlqca9K+zcy0ZzNl34bXRuDPbq2ZKRxQhMF1BUli8MdPiobXWGPveRMYpwWTOLaW5
AmM78ATEfDOQxUREQIa/JGXRl3kQ314yaetXcu6ppKxsNq7TZF9xtZQMVXx5IePuborPCZcHdfm8
eJqJ6cMi2X5m9esrpbszZKtabWOhXotiYLuAhC2oxjRfbtaiYY4OVuuJYHpn8mGWp+ecQf89fauM
SRwIpRgcpDIK2aTnfYwPzyU72jIsbxMqHaU03RfU9JJxsele5/gEi816smVXjeTCVWCla6/voKJf
V4XCFUPexD0iRuV0tHU8c9AdQJ3HYbwyrZJXlgNkLIga17WaFTOuYcUX5RKM+qi4Qn/JTGzyQkF0
QiTfUpPh11wf8ZgaEf2kM0J7I2z4GU/gx6Uke21ogpBLMJGA/GGzBx1OWTE/N3NHQ6UlrGkf2aYC
v4e71c4h9beyg21qAbWQrZefiQh/jxRawAYrRQ+ICYmRBRwZA+k5/h8w4XzRZljRcG9iDI0AYKvb
Ze1oEfGPgL7/37Wo9G3H7spqNEyngo1Ud59Fo314uo+DwVdSC02mEHoH1O/emyux5dCiKKrU7yMW
R9oPu4G7Br8evmjgSIjvtwFBfIA2x2VMsFGDt/BBUXQge9TkPtL0G0akWtF5hWI4x//fmcLXY6p7
Xecez3oaBfH/BxPQHFXPfYQTfOOOcrhr/PkCADc3k3Kk2OHkDMHC9YAFZyPyhiZkXgnXbl+lBE7a
OPJ8MMRVo7rS4ua3QbCszdjcK3QWmLFT7TzJrPUVVclDSyyNzaxc5QeVU1r7+mW6gb0o4/ZNOYPN
GolQJrfxSoUJsUK0sIEDV+4HOT5XrM4p+f4Y/Wjw3BRWr6MVVFOxtH1/08TF2AiPfaH91lDAsrEx
rQaEhQ6bCM9AHExyG603uG1JsZZJ0sUL5iX1fnnjQEmM87YF7RK3Z8il6l9e/enovRqUWFY3/UWq
1ETcBGKzWBN+adPLEqX1XT+yWYJBO2UKh/XDOT8gNeFYIxVl5MGa7Hws97clmbXVnBLAJDvq/0R1
gQpoOSV/krqGoyu1JrR8Q+ks0bWvJv9j51Zy5UelNaCOGlorVpfQwUkS2zwwRm+uxKy14ZKe20aV
c+5BhZr05trxaCqk2f87Q4cJqy2+JuhyrVHGZ/g046iee6vcaMq+gaXfPY20sgazOaD1SeUZ7/Pr
OfAUPkLmC437+4mkOFy5BywIdBve9416xyZKXyutdkk8Wcb3bCs8ZOTRni3XF4GhBs0jvw/thh7n
uoNO4cH0rnTDkpSL92+lIVfAoepH6XZOQFjpQFKdbgIb68HFOO45rVNXpbDKgX+21UpdklQfO9+y
4aEFL3wgLSiOBzENMvOWxynvaTqrKQQkUFx3zXlvnbCplQo99wn1BHH5F5S3GROPCSiLAJHuiuPh
UrwBxZ4xskJUQo6Zpurs38Ef8gJisVHk0Q+fHojZw+7oPuVB8ubt9bruPpRw++xEMQ+nQrriqBMr
oRoqb/hkd8YeNrQyvKKxN7lEBkR5haslf5PADMGwYsL0svm2ctqBjIpYWM5yEkDWBSF2sbRuVWNc
IivKHoJCDjdj1O9PHvaXUC2rspmGVUditsIoO7NrZL+n2QmgJgj9SYrgWekJOqBENrKJyrflXoOj
9sNaPoMDkSb5YU+cKC7bCuqnjLBDMRKxUgl8tFWeNQU3PQtcBdzd6o51T6usErOaQdsL317MVd0L
gopKNtqa6Fa1qGm/FMN0h9QgyNTBKFgmMQikPUSfgNcginLmVCBy6ERz4urSI1l/twcjdxgByTnk
uF6KndyyaPXz2SEUYRhI9S00sWYhTu/op/Y+snub6i5cW2d5vKcs0fSGTY2knDQzA+kcSZ7krJRJ
EwjdNkSNQ+oqqP9PwUgXOKvALPmbSBIMtA5GBTC0PfWHbbMJ6RyhoI1VGDQe3SM82ex8hAjP6y2j
xqFjAu0Rljv/7tSbJ17d/LqsczWSrb25xamJtGAoerxjX792an3jvX+xncXqhsa47rM83So6SW37
Z3fRXTw3YOFtJkl2pMzENmvVHvQCjFjT9lzd0BScuY79kSuaZ/xtHt6JPJsXHXj7AlLAlmLonMah
GVPtqsMGrhALRMfAytTRmGXbEL6brhQueAKkXN7DvXbYJSeoWkAAN8rnwGAjv2hFDK9NWoS6QkxK
e3gTZ5vfcYPPOuODRlQA+xMkkCD6TKcH3dt8gjS3S3z4JbQtPjZXiID8vjWOF6nGJ36V2uv8RaiD
sFmZKShb1bx/BUfL7asDge08eBTnoR+BLmqy+H/PXSjswNyxKQfhYQEsWYVJPI/YO2QRWnsMx5UP
3a37TVzW8xeWkOe1tJzAs16ibK3adiZ1ZT8npF/uF/UI0Pt3Z5nPlkxYEGubC1ObKgQHF+SBsn3K
fVLNNswSa8UlC5xWgO38pwprk5hfSLB0dre54zFMzWniYXnU20nt3tqSHMCu6SX7oswpfPOA/I0h
4BL6VXoEBZ6MBMMn3oUjnbCeB4md0EUGnFQnvQ6uEuZH68u3DfWwdTL4mZGw2gE7zGG72/GzM/QN
Z2xBNTV7iJrxiyPoIKWLUutXtq+EQMcZK94s3Jtklx2pfArpGCaOr16O6JQQLXjexi42UjuDZsab
h3/W54HBIgwRIyXzTua1km+yWRD3cioaX1AIpAubysthT3EfYwwgCy4ZAtSL5KL9gQAmlzzoItUU
++FQZBoNOftXQYdmgzpi/7djFf703l+OJcBz8l8Rme9LiSyMs3ex8I2QHmi5S+91ZlJg6ihm2aew
r1HDZpFnt5rCPfomU8To8imLuleUwKeZ49DfLbmGuyR50o0u1OdO+br7EBurUo59kYhZWcbh/MQH
6AhChw/Ez0Igo0DyX6J9zF1HVaOO+xLG/1Cff6EHURkRtMAF7J/klTvatUiPxqNFSnvLT0JV2cDB
qLrWu5euqu0IEeyC9HiVx4wn+PZI4ne7eXuF5ai4XfOK338t+Tuadrab1EC2++DYDUayLQ4R+Gmd
ga+HF9wEeepBj0dwOhByP8FJw0roX0PGqxPIW1Sj4jMVnFkpDS1rB6cF40PjADs3Vp30g+PhYMo2
gh0ibyQpWgICPxbbAPsjw83dIIQ/LQNwdxEX30ixZawAnbBOcm7x+jx5xCYuRdh9FSwBhPE4Ybsd
OfpyNzDeVBgQ5UjQQSJxmotqd+OvRCRie2f8C8B09kGcWLrcc2ZHA2/nRxgRSVGlGmCAPVVbxC79
BtwXb/UwgtOR8L3vzt/zBiTBHZ61kxLA4zLyBRiZcmjRa1B35U7efVDMKR6w95gW34Agzs8iAkG5
U89wg5kkL60qXeMmCVsQDkBYZTEGEHyo7VgzlrYZd0R2q5tayMA7kM1bZSUBDdikwAc52JkbSGeJ
DOzr8rwIORcOUBGz6P6gT8+VpSRhoIei521kKCFbXvAyIMVoTLwxPE2xw4tB/Qki9fiFLq8JgIL0
LSplRf3piUKlUV5U+b9zq7R8Z4eovMhe30Wlnle1CE9hKTAePTT/Jnw6/pSJ/xcU2fNwWqCacTLG
HwzT7ifFd7NzPzIz1s6O8tWOIvv6Z2PPR6P8zpuBU+hUqCt126eNJ81+vTHwp+TvPkjYMw/JQSxc
xPIC2SecfnkbKwZvGoS3u5wKFbBobZMgo3w3LqHmaWKQIKmsnuF4bnLCe6xPL+JA3INTnlCHqyMD
2Ts+yRiCSy1hzYiZ13NV5EFbNJE9QL5XW3A1CJkDr7FzCVxJq0w20/f1hHT28mIQyKO4RNo77X6e
IQF0MijD7fpj9/rKA+hSi2iVcEEfApSuURz25pvf2oy9H7fhJrdr/LQa9ETXZPqrWCbENKnCOT7P
6RK75KUYw7AJszlP2gvSmth4C6FBNfGW3rrQgqUUR09cJUpL6IDXZjD8ML47VMHyZdjXZly2Q8I1
DVDjp4LCPybPd/CqPelLXZd7GDbswf7nwQo2QQaeNJqS4C3rJh/+BnkxkrC3DHFZ/u3cxCM6pOup
zZLm+1eA5JK2fO0zILmSGSI/wSduPqVh8Tt7NEssrFDNVc+21dZhlWzwvA/KnCV3MYflEQBdgI4l
Iupear/OyTv9RI/ThP2EMKW1WCHplOmzPWq0A/nYSDIt2vEAJMcphB1zwzYs5sxYt+pZHB7dWQgE
4k2Pl3ODcaqzfYHwg3ry795aL5Yt33M3ngU9+lQSRjYXQnxVcLaA+zWukWEwhtjvu3EgACw5G7is
JusDn96NCTVu5Ydl/bjIcGVhDToGZUae4p1XrIpmR9Qmk3y2HW9erkxEWc5pQeOAe2ibA91lwGeY
GZIDbKQ7Isxb9I3H/Cs3lwAIE+OQuLszpI8bWbklqO9Ed426zRalwDM3xiUrtFu0Ozy0vIeKwfLa
ypBt9+v2iEWyxtr3O+o2HsRb2Yreb58AOypSEMqVFhA9J/8OU2/ekrXQBXl8f9ZZhQGcUrtwb8Vc
ucHNUba4sUjng5HsfOhAHyum6SQBfTXNHJT7MHKKx2SksDpVL8YLQy8BpFrcmNh1/1qkXG4AQxIN
kooHyRtYrwu3+RJiTok+QIQ+siPnL/M7Y/PLKF0lZM1TRlOISHmgpuR6e1ZOnjaBQeob5BuM8OGS
qsM0hXmB9AM5xCSl33g69Lk5tFrDmLiNQqURET70fnKfyKcIDt6A36PDa4u53w2WCdVGQmZdpSo2
wm2r7I1ghIq/g4a8eIgA2p786cJ6TD1hnul809LNl5HDvoc2HybvkcfYukOW3V7LTqcfDZ6ucPXe
9Clk+BNMNi/VGOiUVARrmjE2Ddqe48aVLWKKfsebEosGBQwaVEyssaQwrjS0aH06DXTpvkKpadEh
br257lxBCeUburKrcNxYvBFkxgCR2RK8ua02JgAjTaQowfPvCwaNkZ1XbX9rx4s1RN3cF9Q2CIET
fejoBV2bbDn5j6eWRxOaVE3C42mNxhBuz5YDPLgSjT5d3Z7tLR6y2khi1IWksEosNfclyAHg3ko6
kyLlYMbVq3D4yP5VadLiXd20VKx2SbcDBNDPMgbNOsD1ULKUTfVh2DBtdoekdnNiOjWQF2SDxysf
O8oeKAbbyKvhoBzfcy2n/A2Gij8zVJNSZThPZdo9Say4TiHPRKaG8DbGZdrnqjZ4pFC1Sy1/Bv86
lKHrbuW9NIEv6yww4ZJZwh7s63J09O1qZF7/7rM5zGd2mfcjD2eyI5yvV+BWvr6iNoNLUbV0XJAo
8OqLlr7WXV7SWTucTbJY7vQU5OMCRDAj3OMyCXQtYx+LpNTzQbwj9bfjJtGOY9Z9jlDYzx/YKkrv
XyQOIXWBP8MiU0ZUtl4IaO/ywypE2SJMrat6WvXzHTmGirqUFR/Fvf4y3qMAkxNQVw9nEVyNIISj
gMTnkgCy/6vy6njvbxIbaxwQ0x16LQ/Dk4VYNV5zbdAvPsX3pXNJgfXHbh3GSAEBSqN5WRW76Rwb
1SxZNJQwjLJ/A5aGNXogdWq2VG76yeMmfzDouzXaHQNgttbsKTZZhJfrZ5TRUE4x6ju2QdU9iUYl
KZ3OhpdjxKTTcj/ZxXP0bqYdI2vHq4gVKFdjTfXdBGhH4bMRFO9KBvNoOn3DaP4GRePSQUoPczmt
h1GgMIIHYUXeScvbBm5Eow5ExpCAH78qR14uzf5BXmb1OfcgN5MMBBBZC6ywGAZ4MChkdNLr+euP
QT5omceDaltEFU3WzYmYSFohx18jVuUsXxnC9qkpCmFrB+ZJX0ICVFN4fYTYcxZYAU3Wr/jg8ISz
50WNU+P7+Gkiuc58CRKmVWci2jN7PNYyhZ6sYdGZ18Uq4ucl+owI4EHJY/v6KltVPQqRzv0sj/xM
bERyuCAH5l0cGvZud32C8M2cAvS0Rp3u35x2FjpTSkKRSpk8+LE3Kyyoge9EUMFsGmY272G1MVNb
qSF2fNpp97at6C7nGlrg8lPrBkeREnWIDU53fCfpNur/zemZTMrCxkPMme33kf1UmkQ3UEGpPiiC
YsHq6+lV3dbowFwc/G3BSOUuCaEub5wsmE0MseEs1DBiiUhLe7jxN2fZ1JGNX2SVYeJ0ISll6i0Y
Rsz4lx+aUF0PjsGVQ3VUF6r6FGzB+FVoOHzLW1B7V5/BS/fP+hW+5RhAXPoRwAo+s/awfrH1BANP
PJfNvFoOdh6tZqE0/MTl6L6SR5k0v5YFsz6lfTiFSL/4FSesxdme2ajyL0nFZtyv6/9IYHj3DjWB
7ifu/MyNL5XKVoZqEfVhVKr2QRT7Gvrzfouqh+Qt9CQT7bYRYcxGHChUCXvkyo7sgV4wqtZfNzq+
DYuI66J/O4uybLbMkzyRsRoj79jgCjEqC93tByBY6g8/lV5QfPdRmqO9COZpfW7sNCagecM/Sddu
9xR1VrRlpCysd4GJ5sfiMup1fWXIpY2ZHzI1WZnN0mD72zTPKq8A/Py/f7i64b2mMMPPynHggXnI
8x0XjBSmqAYHsnzNJ4aHxxiumjdQztbt3ofeZnXMCxQtdK4umXRYhEHg0VIXnbh1lUDi2SnWs3Fa
YouKc0K1vJcGT6a29vh5IcUqd7RzIACfiSMdLGHwHTTAtynoBn36+9UGHDtCbwNzu6lVZ9LXhwou
8lFh1Dyou7vr9J6JmuY1/yVIk+0DKX6KyLuXJEBBPbywKTu+Ngw42fAdfVI9dxmnYO8KAXq8Pxnt
kiXxKIyhTQ86ZoTuhjN1wFIlf+7sbimEtZuupYopEa74Jh6/9aT5TPb/9yBdm1KEZTDeIDkFfbLc
t0EHKy9gqla5FSzSE6w6oRx05u+H2hLaumVJe6iYmxkIe8qvp2B4TEaUnlT6Dmphd3OGKixuMbCq
gLj2nyylWutpB0I2xUZO/tc/GhKcg8mBE5H/kC1d58GgIN7dZuI1WGDkxIob67JxMtZi36Fuc7Gz
t+1CJrMfHDGyq1HSYzLjAw3g7N5IY041gDqK1jWSWi5Qz03MIuxxe4bHiP/HZdhGujrkzYX5NmpR
KuJK6nGbi2HsRqq8VoZmtcn18zbbTyq2opFGJ1Yp6WyMmPBcZRhHvNLRG68uctJs6naVdTASs2X5
7MhqGZB9ePA/HzRRgAXE9ScSOcPQtiMQeb9HCGQaM24Y0lQDnG7NSwUcBM5bdb0z+kxkUpQn0L3R
i2iF4tsH5m92t7B8GMyQaRuYdIj0Xlt8VaL5N/wdrMcTM2BRnHi5un4ac64H1muLk7x8SJBwUvt+
tuizaaJ1emv1NNh/dvMstz8boISlyKWPW5w12fcErUgzsQCSQgioHvukuIsY4Rj6bqmi+aqG8Db1
jZWIb/gG9u3IjfHfjVfQg2dZyGxCkEftV8DVTbHlQMziEx7zwCaYYowWv1x7Wq4W+UUqQc299hdA
4jidIjELDRmQkoI1d01rgzPOaDt5L2gzl+LVxvmChCxIJ6aKRvzvR3VQ4HhcffteiuKBTZY4lLDw
o38T0qzX+AaBPfjyhb5m6RwUoLXY9N42PVTPY5rOROy5k6K44Qd2HKnIms3hwnCL5uNcvnaQj9jI
0vmbsVFQUcI51mgNeeKEV+NA2BZ8drMcb8pNwkJgobUr3QDlAVLeTPFHkdR4bVAe48j/O9tiN91O
fUX2WBpvuS3pZXbrmBxRygXEyxv6oSPOUl8fzranDjqs0z0C0D3MPIZnGD4DwbsLxXcIYoM170Bv
AziJvMCJhAkaHrczwLwBWyk56NS0iM8YGG8LeABhRsj4J34KWEAFKSr8S8XR5gj6JGT5R3VV3j7U
cHPZymScLBxiUL/lblIpIvzAQwDbOu1gfvdMHqPDLVeP0IjaEgzfvsbmHbfOtGOlD9WewHm/rXHg
J9Jd5rsuvJdwje8F8RncthHUqUH+oQLhm9cnT4OKDfGQ3LW6wwHcY78B9sDkmBpKQUw12GorZcNe
adlytl1ORXON86JaMMlQNfxKPNm6b0F8+/skBGKDXRbgDZ8u0qBMqezSqbBu/503y78v0/eF0iuu
3sM074NBnjIh02Ah5TSZ9PcPBG846qC1XQ5AiXboAf1EHUPdJDHCGHfNm4Pe9ILiEnbKbtpEZvbv
2eRWQedsme/Q7syHkqm/44PV0jpZRsndMMohdLnA2ENdywYOmrv8kIWsr4Y0H6o/oPAEXR6mUvSH
0jqN4XVupI/F8oAm8fnYc3fFtn4qF6caAiyAo03JYQ/BNR/raDII9WvtY/1IiJnKCBZs8cLsyjbv
TZnwZXN5mzEd1gEBWwSDdBGi4yWzt7iW8nnyoODvBk/e/eQmDGcx06fKe+RQt4Op5O5Ekr43SbGd
4Ws/ohrjXBmhLDpIrnVNfXLNThjnik5/lM9ZFjGZqMfhvRS/tb8IQmJZp9pF3hSn/S1yhI10gnUz
EPtHLa/Zr2DlVoCBcmGIZj6C2cYU7tbXJ3QaiRtQC/lDvDntYZsEs9qBbRHaGyMvwQ4hAJpa8vYL
vtRh2JpKCa2zFuPCkGnSZbrf706eM6wdwNNiiBjjF4Nbun+CtQksLytfMicZnL7rfr3lDaVcbCFV
07T6BAqJuhZ2/7ejwI0XcBujGYtQrratH+qIOydlXHGHy4zV3qGy9RvDR+HzA6GCYZOLWRbHtOpA
SzNGNUCFjuVXyu5Rdv1mSG9P+CVMgB3ZgW4kAtCJNA9M1joSMz9TPtpMO7A+nDfTRyM9Mk5ywKAX
6/29gH43jyLtzAbUeV4FKew4RW1NQ0A6CgFGPBv4miip3BtBpthuyfIhFLc+kKkuecg7l1ncqKOn
KpL9exWRVP+8vch48Asqr/nF66kFzkVwMZ6twzXavRBnLaXYL60a8CF/PF0qizxHwSgyRbAZMF/Y
2qMUkZHqq/iCOZhUTr2Tet8Dww91hlW5ANTzNUIgAWaHM1EfrTbez7XE3CXc9s7nY2YvN8oZpvVx
MSYiiWBpw4e/kvrNKz7FcxG/Rj5z2hMF3cB/GBpBT3aYdYicVacWLya9FULvPZmItCIwKmDyWXE6
odqr91btYoNvEZIctqJlSBhyd2GSBnxyf4rAnporzbe7qEpF6baYz8xMw9+wAqNYHpM59tal+EeV
eYn7QSwUWxfjxk6oy92RAfAZGXGtKsswFuiQJ9B2ri0OHmwFRvDhMlgq+Aq61O+3zH9DpBixgI+v
E8Q37856kW7l8J58/p7I6G0GBY7W6rsb7Vd1Nabjrft6NDqiFPOPHMjKde6qChpsgZ2EIrFy4jnW
a43eu4LNE8gSuFo7/013SK3dvK/pTgoT2+njoakGoXAiUR9wK1I9nhimBSuzTx9yCOAWOe5jXa5N
6mcG0Fr4A7syih/cgxpPZ1xMapgVowkArjrNVwsXXexbdCw2jy35ot7QKRxKkKIihoZMiXbn3h3G
abbgiv9CZ3X+n3fCJTKeLJEE0UbMFT5+qAQEgxFMx6Eml55Uau6yZtQlUn2eGo+gwWdaH0Fptejf
OGthUiHutcKuXQwlAw/wkExouC85LtEZzv4ctkz7T+70pMd2LPUPEUb0nGiTpZ0I/5eAB5ANtNCL
vOSfedOjqfaiO8TNR4QGH92paPnIMHCGnlXN61yzYZrtEhBBELtOxzEbDCrmHoZHL18k04NFNT7d
ofocojLpeB9V3gR5tWH0CbzFLg1qEuVTs4dliWX2QoZyaANxRysHJHqRhKvKW3wHnkLOhXrEnJBG
uw0kzTcm9r2KGlwsFHWqR3gZvxPK9K0RNKuI/EFRlrrrI70nKSUEt2KYlN/9vrz1ySloTnE2H0H3
D4DyqAP+C/Mh3XvqK3IxotHtJhOUry6xxR418WMt5zUecnBgmYXMyJSXVMLyxs5I7iZLFOFU2/hB
2w0ArshbvFzJqCp9AhSx910CiFI1/7faY6lUfKjbmiQITQxolW3PKWaAt44Lc1HCcH4iNFVsBO9h
JJLEV9Gszt33cG1HLZsxOACqN9LhDjOSHr8b40fJ2Q+ZvKBcvwKbSPahEWC122UICQXcXOb5La1q
4/+RHGHvjwKgcukAQVibiIVq/YG0zkwbD/aBKkH+ewRwmY/NHukAuY63r+4gkvChSsRssr5npyrN
VDllNUXhbG9kB/pb7GlNoIrFWxiIsKq0BhbrrxMPxSsufOqcjdLWrBDFqMw6UGlQSmM4t7wuSpbl
5YKh1jQbuMKfS1OecB1fFTQssR3exNTmV25OgnPHMY5bGzn7/weI8hvf//UELLnWqcUyc7peQ1XQ
EWdMxJCS5fDXxJv5muf+9imjNwRIkAAA5E+Zm7YG0OIIWDFdy9nVQIzuUY99Z8AsI74oG8PiSoL7
jLjCuV5JXO0F9mZ0llidutw1OLxXTmKrr0qiV3bOgLJGDEmpUVVfILn7PFGnpMjuj57jcUJ4039O
zKoB/GM0b3vcHrN5Q7E1qNZiGjzKTjA+VvzetjS3hOd/+7jRrESptRU38qhCp9KyI6xzcbQcEQx/
qZpJYA1tDtoDpLaCSq661h81HFZKjbuUnTXuGS2o7zWmavLClqXDhGhlV8KZ8dL+7Jg7X/wK/Cls
QMVH3szUue6Cqq4cwtq6fNsoYnK5f1vtnD4BDffh5Yh6AqIbdJfKUp4bdUV/UixzaOyYe4OXz5z8
0vF6NFkozQvOl7QLqGGPfOH7j7q/kdLDfyq/oxYymtYVCpdLTwDUf1Z/viUvHJXooG4Mj8Ghlz95
F+72f9P7THK0Dr1dzesYddDrS7ZVylXfacEAQ+DKlV51/F0uFpHtgAY+Q2jIG3uYR84xXc7ij9GO
BVEmSkwDlrcLIfcyy8uWEgtk/+X5Km01+Tr/EUNT9xwbEXJiKcHzgZUUcZIHxtRds53hp4+DrkLb
FapP7rHKvvDV9Y+JhqSmRxnQmZiSNrE5eoLSZZS2L3y6st6Xr7SbWq2etr/CpAfVDvNrABUsRO+7
/yPSTLTJFmwvqxpn0OFK5zcjLSpqUopi1N/Yj0wCA4qkwgQ9xQNF0KUnhSa/mfTjfLvo0fUTzDXh
pUzRRSZPQv7utWNIxFz7uQ1wm2rN7Ap2HjFiUYzeti5h/XM6QgRuetiPWAxXzuDZ3BHwussIZ50R
OTWmDgXFijruBZe4CH0ZX4YPG6Es+GRmpXTxYiYgkx3hRQXyq0OPbbf3E1li4EQmIcWVm+7lgVK4
lEO64PV+cXZ4juKPsJCRvGUEcq0YABzIgaSUpsO7kZoRoMTAL5jQB4Ao+2rIxS5DYYMoo+ooO2y+
vLTpMVXB9LnJ9RglnYHBhp8dJUd2bjzWAbcvlNuDR234zQnIefCAYUzyC+5zSNuW52kRgMk0eprU
Dx8WypgY6Bji5CpMUXBygkI3KFpi49n6ihcSuPizI40fJJ53uYq3rW6isJPKZsMuMLfjABlFW3FF
YO8wDc3UVUFrq/UqpcTZ2REHmy2BGyxmQrzaT61jM2SLO1FiEtojAgO18Uy+bSvyuF4dHDYNVLBB
eQBl0zusbW8f9+pAP81OZQiUens20S18QAwAcTAJTiYkxhGLxdbwRDwqW9/VaWAMB4DQgSv1JK9N
V1iGAjoXLRnhE+Oq5YoxDqIxlu711eyZFXJjRzrycwr0ktmSnJs+NF1jCRlODuETDN5+onCk1hEk
Ct1ISk8RN41IF/AnE0lf/KwC0ttnx2r9yg574TqutBWbrVZHIWB2onxw2qa1TJVUPekks+GWZ3L2
VdZNgq4r3cuRJwRLAxrrq+1N4Oyv4EoANnJpPuuoBDiPpRLoEUaCKdCqTJ+5RiCbe1i7ksbnvmZy
uRRW4s76yLcklyDyl9YI9zRpglV8KZfLWiLhcVkACGLCQonE9e0EvDpIZxk/DKR3bsxkdl8mvV7Q
whvWM8+dpjXLhS6OJGDhL+ht0ns8YX3gnYl/NPfJOLf+paCxI5IDJwW6GpnOOz2KmHeLj5xPAwar
mv6uhcGvvzec/ayRN8dk9lMMzrBou8Hqfb6ZknaPqlnHRs995qto/xxMSYPpmRvQ5wsYLoCetpts
5PUxJUiTEjXbgNyGgjh+EO5VJwQ9jG2ctG4lLJfm7TMv+yaSINCQtgcHa4fpgT1BOWRAEWXAC/po
56MEPym6FbhWNNlVhSUKyDsl5ffP5ZbvyGH2mc9o2fx2empt4J+VhNtddOwcuoQBQLjNUJMhCJIz
Yo+rp17mgLGJVH5kGtFiScHKsdlOtHlqDTwyL2nG6rtDypK2Uig+Pn4LcfhG/jHnwBh4DskPGmEs
uNmfZTPsiqun5qNbvVZE5GM+p4Hr8J6fIXYivB7GcBTaIM8cyek/QcKnrRC50mB8i44Oc5nk7VyD
NiAvgegiUWO/gpTfhvmJxMSl0dnLv7LZDKP8FP/O5sbhwSiVpIkaV9kP+nbyLTsfI5Jg5JYlP6Sp
c7CBKBkgV3MQfN7ANBNn9PxdE9jQZYabpoEjARgeMFpeg5Ljz9+PeJoo2/+8Hl6uN/nTgzFxZwCt
S3U7+t2QWXJr3mGoj2MuQmU76mSqMW44bUibmZGNDevGpo7N0c6MYBXMnOC57aJ6e5uSxFc7zaIf
eRx7tG37oLtwmaUDHX2RiusYKpryGa3IuhElt0nzouhprRC/74HOtounwMn45TXeEss/xEMi3dJB
tlHLMnRmVLhA8hv3vepnjln2Hox+DawepF4rHmTjNysd4ORtnUkTW52MB0cHDMlA6D3i0CHlMAea
izjOx9398KtO0rkCcHUyJ3vB8vSMNYv6yNGQQE9n/aH4g0xHowRPIKp4ToqxyWQNAsCDH5P7E01u
0iuuAeHA4+z5hELdOeaxho41mkoCVNtTBIIIGoIi0TBCw5t8iaqx/A6Wtnb1+6Hda2ddAkPsz2zN
iygHCNWUEWYJ5hfwYvAaQvj5DVuWDTdofKTh5XwT5amkAH7svDWl77gQjdMC+br4bd/Wg9zz52sd
lXe0VIUg2Iy2rTnoPRHa7rRGRUvphYvZ4cgI8pCrznphqMwekQxrrL+8OXCYrjPUw9gNK8xEUyGx
6IbWMBIBWFKTOarjw+hPRPiRlHm/cEy45lj3b8HhotlWHDTmJRmPuaJc0zfYDDVl25i0w9ZDWxbE
n11UysEaYp3e11fPnY+VEEz1SNTWtlA+7hgW3hhdKnDNHbhZKl2uJuaHXWyTI6ffLuLicogQtOhm
Nem9RaJtMjE/eifwbGKBSZqROpZWr/1C2Lgrpq7OYPpn+MdSFeh4C2jhO9nrl6H32Zl7FApEz/32
cFJEyR80cXT5KXGCYKmrDmkp5Q+0LDEhN4f9AHvLVw/XgXoO7ZryPb9aJOT/Af0HB5RvP2Nn24yu
JfSfcTfEE8Bk4mSzqDNXv3atFV4PXAK3ZrQqyu2PLMEXH7h+WpIG9cQdWFO9PwJXbNozrtZUlD+K
86cGaktrGNB+OzFxmbYJ6ZN7wxTVAOSrF8/fuP0IKpevyITsmQvJs5mMdW1+NLm2/cZNgLgfD0F4
eBWRqELcQwDs1zFZn/1zwYeQYwaWUJoTlR/LxsMT4gMAvKz6tQdCF5b1khLMiphh9U0fksZq9Jlm
d2GxNtb4abw+GRUmSPZZxJd6ZFmJUognXddWuWBy7NRswQSjziU/M3NxwgZYtfqFeqkTuH83hA9s
Lze0wvm89FjGwWyBkDz/y2NctCxKM/NM1BMYg5RuzEnSKESG3YgjmsqvkKz/ugTkRQGUIIuIp/T5
nEz1/3SSxVz4hQx5b3PVGC0WqWqRBehO4QKHowQR3I6neRE/GkDHAH9R1+I53RQXMCJhUPAV+37h
3leQCR6s6H6VXGdh7ufJU4/poLzMrmRr7KEYnyPj8gaCdBnyUTSCzbqippdFrsIF1lbOsPnj+0S2
Nfvusal/wrF5TIS/daRmKs8EirUFoB80blWRf+Uvl6p/1Kpd/9KLPXFT3utbWU4ZOgFeWS0MngDs
6sV4XP0vM9ax5+yWTRDAbQPYTicQazso8eyjukp1/WVj40uBeHThCqySfJ39Q+vukK2BwCNBSe7r
DZAtsKEQ86pUyNlidT8b1rvin+jQwQP7fJpORqt8JgV+9nGjniEAbwbHW4nS6ePocZbUa2vOQuym
yRzwKiXPM9ylKqLAC/zG8/gC2OiMXBa/Bgaikmil+odtxq78+XOcPnbMvllYghUwJIU4RXdfC4mA
TyDfFPprtr8+xh3mRqmuTE59p6LN711Z0F+uXZuK376vjoxC0QHQtO8JlihvmPwulmdd4v0aCrgF
oYJYYIAOPz2tQoSD8i1csBTgQwMukYbQAh90Yt2iRY1DTfTj2rL7Sk1HAv0swcS+i6LIqtAAITI+
mHzQcd8+nmfdF+HcaQlexzQ6kvuvmffGN/s/caJe/sxcBlis6B+VwrMKwsHeFxMOhin/oSa+2vfA
LoT9ulq0jrZ8vIYAkPgZuThpdQdRkRLWUu5Gkr/wxejBxLPpPIsqwOxWkLr552OpjAQ4OpRMkLNo
9gRyBxpANhHyybm97Q+N8YDZQ3gDeuU45pJIiSq285FNmwDFOVrznPF5tyfVVD1tio1w87R5q2Q/
Fg46r5VM7FECdkrphUOqvh55zuW+dijkwIh7O86XwfijUrjZ5/bQltQLntoUhywOB+pf5RkyAXI8
kgc6NU4uQ5kWIC2JeRFnzaSwdMt4vnvKOxY/byaFC/zvisLFA8glnDOVOzG0h9sQTUZ7EeBnOL8g
DErOX4ZhdzgmWQ2qShyGebjLYCOFFoVFjbew36a5yzndUorz2IwvNCtzK+Aqpds+fuHt8tf1yBsA
FdZSJ7CwDBlaqO2NRJuKP1IImaJ5udjmyXN2wRSve0M2uvWvXBW/zK8sy/OLRGtM9QPh0uy2zNre
J7mUvvnlX5e8EeesKJuz8rOBLRR7TNmymJN15G/0M7OWl89jE9luwMWPtAvqlxAxW3tGVIyPv4d+
3GxMqX7BfSzRxQCDJ/2xRFvrOZemJS9AURzh8LGTDbHRiDPjrU0SvR9FNF/v/3G1rb9qpk/rLP+4
OT68y1tXQ+XsAWb4cGyR0VSyrjEmXd6+8vYDqTx8k98xwkYWW6/6ju1brzWq/FsXbbUjW0w3D1VQ
ORpq13tcyESx931iWniS+JbaIdZfe2mPUluCaLyZKev/oJ441pJ4r1aI1qdTXum7/tkQtN9KUQih
cPD4thFJkyI2gEW8FiBDGK9F/3d0TJ/gXL/JxX8yQx69RcygbdoMQcw96nzuXoZFlH+EoydbyiWa
8Dw2hqT6oMtlNpQb9PBvnbmpIsEOfG8wTpl/EUx4cSMxXC0MUT07UKfIkssZ1r25qi4cAMj9bxeA
vEqIk7anAHEot6nVn/eAOcozHNhL04jkxK0Ht9KlU3jghrQ/J952pksGGmrVceR5o/ulV/NZjGDm
ZUrurtYevINuNsQGfYkPA0R2DXnPlhtR8ig8YXe882I/QZ8vF+2cZ4QHTRulSxDibH7j+zDkx/sb
p+w480vRpnIZgQzGgwzdxWkhc1K/tXqSrgwnTdSi3I/Byk/tdr6QE7FVhvbnC9csqlJfO/DyMk88
igkuIVG6gp2NxcGZ0IGfvH+wpjzLk57PIaPGrLl7Vn4kVMPp6dzVNHe3LRximzDh1Z5xCcD/Z4ok
Ih7m84fwQaR/+3Gc21uFf9muhsNwFPijJU3r9jdf+y3hB9yOsDEid66bubHtliY8YTKRyZS8YMoV
H+SQ+/TRlkSJSiSD03JZxDpEqgAfWK9Iyd/0zusgAuQctnQsbft9eCBelyiAaSeiGDBkSjX4yahs
JRty1tt7DyGawTrxpLgHIoQjZwXkkvr/d9jUR8KUDwSX5SZAIHn8eCmpG3cuwkXElf/Q8sAiivig
Cjr1IJxiRiNGK7xZhEeAvNakwm8IDGmbZV9uCefWyMMtZilFMRoBG8qfC3WlJjPZ/QSIGlO7hc7A
YU0RRxaiXoOJwlLINjEcwWMxSQF9UJzOGHbkbKsMBRUF3jyu6L2X/m9DcIJVuOX3u2yCIHircACq
QV2vVv09Yzt6HYpgzbL7INyQbTKOFhC0pqSklfKELRFK0P4/8m9+Pi4voFv8BVh0Xu0UEFVo4Txx
NmAXd0wA8E9iHdV+NB51pq+JsQ3cNs5GCDFlCbw1dcc+eVSmGvThDBmIRYiwW/iBc+LL5XdjSWTW
pgJxxmDHP7lgLqDWIPghPT8afCm2DectwMzuuaiV2z99fpkLu5FmL0XAHJo0v5tmSQqiugSkNXdF
F9V9LQ1KDlSvpg59Vu32pZaH6f4jzTlpYdoqZy46U1DR50mRc7tC5oHEs2Z74oWm5o/hhSYvRQk1
/xKm3yWZunsg/U45VHDOytsY4Kgj5WsT0Qlrf3tZW0ptRwlVpQdySbELhdqlHpOErbOHX3m/Oe2E
JGyUIYYKZs1GsDpb/6zyyXgkf8si9wplO9CLhvmjHcTU3df2aym9+QpoUCD5cuVemS1ucSm9vb9x
RkoVUaMmLFQF/9ZkOU+p/9GQvnBbNypxV38DYLdiCgRu80PBVQTk0bBm8ZtJagNqC7en2crhcXGN
npy92HdYj4CHxCTCaxRsNG96r7mumReLRMHf8JJTdwuu3YLPuk0TrT75ewKkA4kyy86qvR+iMb5e
682ALAd/1bKzCds9226KfoR8Q0HONOl19Vpv6+SB8FtpiNpB6yHwJq3BlVKFqXkJYFbXO9sU/+xB
EghG4ZOA2KGBytsXYILWq2IBMq5WH50S1N/AZHP3AWplz8pnUFaGVJQiihxOEWED0IBmXg46NWbS
vHRoLIsjpcGYMqI2c/ArKOhqoE5rSmWV+LqACGPd16eke18SdqwKgZvCgiiaMVb41Ma9+97yIu2x
zUhQHZ+kGCISjQeY5+Cxy/TGvKfeBlU+zMb/mB1S4AzcZ7f74jLYzmhLvHtaGCuAf2qHJ0I/Gi21
70S9/h8gFhCU3gTUqJEHQk1vbnFijiBUY9Rbe/60B7awhJDEGgqqL57bDsIxsEQxWL/p+noNx862
lBBXR3OsuGR+kyubva2V+mQQQf1dOEE5mDM1O6ij9mj7fSXKcfuAgHBZn++wHoEJcqRCpWULkqgU
L6r0AXZMWEMJaeN4KyxuhlbBnk1tJvLQRsbs5E1cVcnMnIamlT7ftt20jXDge4gKKiDjBODKh4IL
z4rofCCRgv228iywPiMOjI1/tFAqH63BMVHjnkrFJs8k4qJ0xgjvHn/XM53oPPVfPSV8aZevGMTT
zHipSgzRG0JEe/kYr6PP84aI3xZX0KjrZUbmPyNFDx77dRdiunCwhu7kkaHPvuFYSEvgtiM2UH9Y
zQMANNO0lYY8fR1OgAB+iyFmbcqyax/0jyz1ivYqI/eDZyS+6Vvt45lNeDsXCBVQJwB7AOajayun
2Ix0M7PKS3EeITBVLNU6eRppOVgtot2YsKSWePPwW1zdRMGHQ6gmJBzptJQiWUr9205xoC1v9OFM
s17Aq8oCZBl5UmJKlnyX2B29k4cPc2a+LB9CMfk9n1ELv9m97VmPbCTN/Ru8lt5/GpQftNg09y5T
gFVGQsWK3eDkjvSwR8c74WqoNt3Tyjnx6ERfmrnmTL6ozZPWaw005IHlzed69TjP0VRXerTqLlZL
2/8TvZnBiR/XopbsMm9HN5MrNLVB4IX6b+osMnUMojpxaYmCbj30xti3StIt2JoXfbRrYl/4KL9v
8UCcu9AtAmiACh9003G5sH8+Q4BkgMvSeRSXUp/PpJQTDJTwYimgFGv7e4N6UItv2aupY5eW7Gwn
Qyj8AgLxQPEGy/t36NDadZS+mZXKp7XrJFaT9/wpyLEPY2oIZFLifLUK580ufl6XfgMB4gp+q4TS
dHYsaWHqf3cCIunzsw2kNVFzKp9nFkcsKhn+XWuMt/3goGO4ucJf2B+jk6sF4NOzGTzEhl7zZOpg
T7LcRGjLnIA0WhPNhkYNtUeLNN5l+hITqeXUIUgfQsSj/04zK+BHJixa0epjKdMYJYG6Mg//QDXo
4QkAlqXIb1uzLa5iHbm52THv1VBtiQTmgWy0mQU5+cmGmnkq9/Wkr5gm9/8f3Bk3jTVQ9h3SVx7s
wR2PuO889cun9cW/iIQpMzGTaFpXYgAZpT1vPh3d3shn/yc4pc2BSrH9Rxq4W4AuiR9isPQe9ZSF
LrKyfsji7ZqOWRNv1ODW8T8PHR55hvvFvmEaOjoEoyjrLNFxUGAYG7P8a8aAnzkUx99RH6ybZO+2
vgWdkXFh+9mx0fEn84ZpZLwTCzAhE7fhTOooUkFarPuLzEl5uPsZ4ezJQsicm12vZLSdfjNbhZl/
fuZ/vtfk8fSUAKchZDYs//34cithUPWNj1F0dyqYndhRtokdczbcL4Ebaxd36ERSZMxJALPm0Km5
2+aq8roLVmuTHDqMoPyZOgQrmXV8ZA4cIn+GaIdrzDTT7zj296xvdWdPejHCdWgeOGoMDkD3Ooj8
t5WA13QO7dIEuNtOqPyjdXUbw2dj5cOLFNXoDl5R36ikzSozPBgMc7ToS9AQdyy1Daqg2Fu1xcDc
t9xITQoc9ms1Wj+53lzLc2tyM3H9GI4lw0WAq5Pc9dEI3tip70huC6YQzQTPNZ6ihSwZb8mS+RGM
BahIQPZnGXlSjmgZBMsYZy36EMoNnfVEEL/8QeT0TlSZ+ibHrAJn+iArBMNC9ozS+LBHbdUbEK4J
y1WfJTVLuaGxpahFEcrroMx8dQRyPVO+in+rc4ZNoo6fD8MQu/T/gYEBppK4TKO1XbznjJ2RbEoD
Tazl7q0orIr/QDBThLdTMYpQvu25a+C+d/5Ar6xcka7H9o0Lzbdn7WxebDhkQ1JNv0Lw0ISNp69i
YxXxP6L3H9FmttLEcy8Ts5sm+mXveVd162Mv2MqWA3/wA5cEKm6f/exmhpAHtHjuRdle0E3rIhbT
fFVaikUGpK6tJUxkudLn3SmIFQi4XNUIReggvBcfp8fklp4p3Y8aaEG/lkLEMnJO39jJ6xvcwQSx
FvTUP7j8RbJojiVdZ3BO0QXQJ8HWuhVqGBGqK8XPOaRcyqUCwulWpICQDEGlEhl9WYlCSKrhpbHW
rgDy9N+m41ssE6HIyG56HQd4b/KgW09jEE+7GH69X0mxKQ6WaGiSCrw6K5Ybt117oNQVyReRmvIP
ymcOdgXYReRHNW8T1cP4zzjYz74FiFLdsVl0/4N2Yxm32j7qHZLJQHrdfOOleEjzn3D7baESuvCp
AMVZ9xFoe/FgOBItmv56vvknZytStNkA5lXrwlBOiHjYMYnq05W4myZgNwyPljPZlP2srKpzoFfA
3QwQNlmq+YPmGhY77wkbTe5vUnyXapMwur2BdDdmC3A0VxFD2Gp1c7d+jOM3qSyfxh+N2uuEwNbm
P/ltG/bHY4uSnwb9DNmVLERh01Gikv+Va8EfO1FCw5SIHtTGFxgyvqc6ZM62n5Mal/DNlqU0aSoq
+rDou0pxBTE2IrRr4JY5W7CKQ0DWRvEASRaiwZ0p24p27DVHmGgbqO1wDJrHjgNHtST5fi/NEUlZ
KEmlL85KiICUYxnAZiZRHcyPXCWFiz48LtNgc8kHVaEGn+PF0Rg3Hp287WWR72GCKQffB/+1jZPT
Gy695wao1K1yqYA07er89xH8b3tvWubFkARZZvDMaqQq/p5qMKzbwh6m7+i6KJmokDvREf9PYWZt
nG8bGK4+1VgeAE3hMdOZdrOYPqDjzyObmL0jYCNP9p7dwAf7SgphyRPeCcqZUa7sL98KV5BRevUV
DCCchiP2v2+EWQbH17S3ZDVgNPSt4RAKoAJPYI2X8ksuUOSbxg4bPokBE6NWsIwlaYfr6g0YaXeM
ItJrmtupxX6l7WKg3Nnm7FHG+MOLbmSRBnAKmHg3rzTF8REDOq9XPAFXqX4ZwDDvrJhlY/K3T5/t
pOoru9n98h9rzq8X/lbSGhSSgJ8q3dJpvQX/tjDYz2P2Creh5puDW4m4XUMhavDpfaBxMQCCTUyb
vZPUdPeoGIccGl8Y8pVRvLVUW2/7qeb/B4JCpxuj/VkPnANPMjOk9OVTypCgptbSJ5lGzoVxMEs/
HfOZGXA0ee3ShZp6F54+cLMhOSywLZY37Ko85SXCiFxqhbVzysN7qQ/nUetBe0QSNit3nHF2fHQ5
ij7LMaMp51I5loKAv8PqakU8XdPXRpItdtQ9/MA10YP6lFkJ2GyGtX1ZyAb6cY64yyTDD2pPMXLe
V4t0x3GDs14QeanqVA/VhRes8pKkZWndbl3T9asqsnRUUSRAkZLcmHVngCx9O+FiDh9R3d//0YGD
hGHqnmoeA5eRdEHaWCHZDtU8QVYonyAFjbl+NGFJtAvCeC5vXmX9r0E4RAAHL18sAtO1Q20GcgRg
vdnbR7vCrJTAnglRH3XDaD3sJyyRBQ9Gek3YTt6dgysvfSOAuQy3ycXZqiVZdHu4WP22VkVgIqWt
uvgUL4XdaArG3sVBd8grP7lHsqLazb8AgBNVAFcuqmd78rACScMI+TKjB3OPSXNlTE/D8X+A12dp
O83E7wr5UwsgGdUvwzSB5FUxqhttufKNpO8k1aLXMA+rvhXmudQj50zuZae1lnnm6Edx/lz7dQS8
06P3lLUfNymEJOeZZuujLtU4PuTOrQZuQ55d2RtaLltpbUzwIXwnB3/t2MiqA3fvXibA/6LChVGU
ufqtxYXuAkX1JMDBdT5b7XoAbLFEkE/b2T0sXGhVRgZCpjtQLx4yl7ovtMeXVngJqUyllK4BhuRz
iko7PuyAMmIsZqHR5y57BMsPGXsSIxqz9NZq/6iEYWU4krhmfurw4F/QogkO9hHMCkyn2jFl7aL2
MvyYb5UbKz+v/vMCYcRHzf/YGl7NBymYwOO2YPwhyhJcSNTZP9l/A3EMerThoLuLD44swSFMlnvX
Ci1l3vVLlagYivq7pEgsiWWoPFA6Uu1mLxlg3q+/UAPeUrnYz4+q/MbygpArNXMvlEsY+rj4+7FJ
d2UsTegjcpjugwdtinmyZEHTaiT46NhiWDupd9YgW2rJ7Qnfvw2nNeQ4nrucYOVZ+VsT2RLSHbmv
aL88IUHeZgL3C6wBEDDuEP29/6VcejZ6ftMmI5Y/pFM+u6epbquEejPD7OeBNO8Q3wl78k/qllRa
HEmAhVueaz6CpUTTaOjdZbYR1DN5dithVg7sg9qxTbaQQHQ+8lTL/maRXIXeavJi3Wn2FV5TjuU6
fz47CWF1QHRPo4COyapxowDA5p2wGClj8phJ5CiW8BE+td/fZugP8Dw7pkQlPRtxTMGmbcO3u/5V
hGh0gmxKzt1r+NBMbYnuBpEF82iYNyn/8I5yExDlfDRpKLhAw2iEYz0MDws111SHH7MTuyMTtdO2
uvVn9DwLePjjaxYLNilR7F8zoa7pMDn2LLJBySBMT+6bRwUUr61r0ggvvcNzCW4eXPde207Mr3kf
ZMohS9YRkg5f/Kei5M0HBUqwBQWChAal8mMAZUKALSa7hHyt0IcEYsrwUWsg4zXuEC3nkLEBuxIw
HPxWUZemceeg5o4aVNGbBW8gLNZ/m6kkLSI3pS/B/kxR6p7T4LCFpe7Pkc9pPDZPc4X/TX/gCDMy
ugz1ceo2iMTtbF8Ca74UnrrtIg31u+xuVbVBHcXt8n0aykApmaFt2afZan0piFKMoPBmHE76N1T5
4lubnsX6MOEIstnwBLLkfZJX9ifCdbwXp8BERZx+Y8xbyobOFN1YYDy74R5S4VPi0scJ7HxLhPXx
3VXgUT9+Ud6lXKVljOd0XFrtwXFDlA5+V7+XP/cdHN1vZIagcnjefMIJk8QdzysqQGWGVkrljU9c
PedfFVgKjV1J+tG0YPGxfWdyJYdyL4EmN4L4ZaR4Ri6qfA3RuFtPzJZ1ynoxNrvMR20OxT1dBIYq
DtdOmquKklaC+sZTAhl9xUQP48LrubW8iVSXa4SmSaGdUVpjXFIG5aqMZxTAl8Oax6U51FCcpvBv
qB8qas19y0pH8a5qzZNrIehvTE7gyauqYr17BFh+q6229lzHqzvY4Iv1ejd6BK4BiE9QwFSbgukh
vBENcGGMz4+K63IcHIoLRaGFqPzcHpvcVGCqFoL12yIoop32LqW3DlVJSfozmbEVydpLlSrS+tnO
LvljKzwbYdn9r84GOOfP5QABS1o9VuEvP7sfIARFF7HqeGJSQUj459jy/yxDj95zIKSUCJlVwtm/
wvSADS1NF45k2AyTHPJ0z+ocACP9TASq3CyXS8HLjoGuXBEq2gpZG7LQfH8imjp8S9x4pLBDGku+
UmaXIqh9dzzGlPs/DgzjmJAMyF5Nel04jGqvnl89BoptdOYQ1AijzB0ppeNh7oSBxnEvz+xfHyRg
dIV3ciz3Ab1rw0rySCEihmLup8ftVw4RFtVCTHR2jwqH5qm6lOXIgmepIyxUWEAIPQJR1wNG0Hyk
nZ7hKQiyXIyW/3u3vLBVMKSxmBIgGiubmdHAM7u1jcbmOe21nlLvEarJ5H2fjNf8qRmQA/u4We7F
b/fq5RO0LOJh9++fNVEHAeBtgGWzbyDHkOcNY25ifB1KWhIiYvJxY7MoYKB7tBF57eif70ygxUnz
8Gz7kEd6ZT4eBVSbFOySrmIHZ04Zdbg1Id6noeR6Y8cLSRH0r0IauGEoZBMM5ac3kVz+aLANOYqT
/SSQPlKcckPYFOeq4MM7jknSf23D+r7XFP3C9WZgnGUIr9IjbDAI+kQK6AA4ZaSYFHs0XVnRqba1
8XJMijAX9jxe5FhAEgXC+nI1HFmaIQ/dJBn8FrD5SMnJsxOubCNBNX+PVVDuDQzmSVDNyK3AQIsI
t0my2Q9yJcclDFmqflk1Y6ga9zReSJsUnjDxrDF4ovYxgz4zYc06C2xZIwSZTtbFEzaxIAfdHejX
WopHl2c6X/m9Ni/8zSXczv1+81wPR1hB+mIfX32itH4A5NkGA5yrwlUbX6uANlfWehIL2PMUarpE
IRoJHg9zdyZjVmlpj2SoPGESZ6TknQNTIRYEONylpDMCVvgbsUXgbRq/2bpE9OiaITCzVW8sHCjX
rqTyf0d0tnCzK3howqEypmqdxSPrsYAhOcCLG9AK++aUkrVdDdx46ZXHCnQ/RBeptZuDWo8jLhyM
rUWSmxFU+Ag6aZZ3+FC1TnSKOfA6sM9kaUjoDGEkh1D9bt4R2bRVGnenGDdgaAqvYLwjScpHuAMN
1rDxc/7DJBwudO1tj3kNSQXFukoiynLhFEmmxIslwzOutromNlL3JavvcREVeg12Ifs5E1CjvhN3
NKPadCshSptgnK834SfQkq8wVFQp/puVi/8YE5jcSLY9wRNJm+kpCvHPTnu3mt7E2tabLAuR+aj+
ZAiPVDxOo63tv2w12jWmOFXK5prR1DCIe6NK7IydvmwmW6o/Z9mQFqQ3OnD3FRrG2Yo5epUXI8mV
Up0jAfQ36mR+RTm3FLJdONN3t+O7lDpAUTZJOVCuK2wp4VL0wr0iP8Fhen1YZ2lBhtP6sOiNmRdd
aNSFUcPhvMBXjVlGtO0mLKiSIsWEbHTynN9zQzML8fXHM3uliuqaFyHf86ufLrDCfoRrDb19I81w
FuSXnFFVEy5z4S6tdN+SMTo20PNJJAcaf6CWw4LRRdexL0oz3AK7VW7B8w82i47psA+5fN+JiX4y
BylOC6V2RwC4QODJW/2/glE2nVhVXMhdkv9TkbmVq7TDONw8PxUYt5J6v4Q2XeC2AlOERZSuJ8aU
C8VeA+eCI5hKQoojyy8TEZ1Tzl5LgDQQYGyVIIct/0zvtJFaZWybayrUBIvzxwH0ivq3l9Nea4Gt
64t9pEDUFtvgcW+WcFwpjCax4Ecyg9cwPdmdqhdkOhTpIlsBdUAu17vZ35xqcypTmqQf2NYcAOL+
YdgE6irgYvBksqf9zloLu73YYO7b4MAsaTJauBoj0/w1IpFpJQQ1fPf3299xjTyBLtO+L22SHYSt
21pBWHG4fX5/yFU6PPqBxFgUIju2R5SSwcaL+2mLsNNdeqwi642LQ7otEr80jOBBfSYCmBgrTZnE
N/0w1ningOOPo4yfN4NmwNqF2EO0N8Mdkb7lU1F4RI4LykgkDFgl7hnUhXiF/O1jGu0AedFARQhz
nCakCHr+h49V9bkBDi4rQAxiCBxSKhIcxDFiOUuBveF/Efh2EWxU7Kw5w5iyEtKMNu4VJknHBRL2
VnSxjQ1yzQ/B1sCgguJdmElyYFdASnx53n6+wlQ8nyEq4XZ4vQtVuVlniEcjIevItVrL6NyqA28k
VrPEVfMNwu+/B2IzdCc9LZ/NAJVXYFXG0BjRKoUNKE1i4oEBTkXAHmTB2tUkHg0lQhMoy9dh3rWi
lfvbbAikZDVUABcLahj+jr1XzJkAAjbBHSd+/mnztq2ZU6MKuMCLolD58pbXtMgIZuOn7YxBwpiG
f0tDxbXQkNA6g9SwSGEbRt1J++cAN7CfG4ktptOUS7kjAJk1k+0Gc97OeuXmppPZm/G9inXmvWn9
Dlt0ZIyixcXEijYDpthwUiB1HnLpFL6lDT01Kc6+jNs2oxRrY2qjDFe1hHCGYa6yhbfZHMzu+Uvr
ZyDmfmGHALvcOahD7aLGvvcCZNZo+QjSFf0T2wcVZJlN2ukcXfLx7HUW6CLMJOou1d4JDFN0aMyW
7R4ZmK9Ujr8zaQ9CVrZS6ykMErNjr9e9ShX0BafBknKX3+DvTpQwG+3xhz9M0m/wjCU3eazIkcNa
ort5TWv660Y14h8RrNwwKjxoVBK8M6dGPIVDz7D3zh1UeHdqQIwlUzqU8Nl2g9IaqePEqUr4p4ea
Qn5yX3hMl5WqtbxH4xhCHNxyoN001QrONWBMCNsgQsd7hOYgOtw+lFA7BZ1Qiqx20fKbYham9rZb
oXmdFeYVoDfV8xu1unNHYXrhhynaIeefHqav1AwhCuFb91whcOZMhTS322k5Zm30ulAtTa/LZnNs
GMtiZPCO02DYjpqYYhWEC76BQI1Jbu93mzclT652/dHN0Oo0tM65tU9tZL+QyERT3n3gaAFNU93H
Ds86uc3k9x4W7cuv6In+EljCA8L/tF4jGAeAYxhouhsHM5tHyPlMcHGBubpYycdkey9WPFY98dYc
fEMgoxn9lQEdHkq+WCXRLqr3M/QHg7KR/IkamZ7i/yzJWz8L5MCxjyLfgimG1EAyz/Hy2yhgtdCG
oir/M0gYHRBP+uSH72AMTKrXHqgIizVnSTHNYgYlTA5pXAsbeTEUfiWlI3DLFCCX/AbYKM8iTy/V
n/6qi8n/Hh1LblzfU+KrP+fOanObEIe16lNbfqQIgSPxAVVcud+CjPJ/2DN+fwEsXdEeWmtEEETQ
ubCRalfbiPXz4oSi+tHr96b3b6ywJ+VFL+4BxfStDOXuYLMJKPIdX1lcx+7deUpMtBdBTk/V3ep2
DMBwZVKxrbzga83RY3XfdgfhroUU3ZFO87D1UiUyuCuYG3LgNeOXj2ICdidT0cLlngAqTleJt5xQ
dsV+a0TsiXIewC1wqVpKhz/s3zrhxP/AJHdSxZ2SXSemvcarzfhZpIu51K9mNiY/KT9i2dTzVvF/
HgxwaNaNvZA6qk9B/YUTrZyOMgThFzlY8+sHLGqgdDLSk0+tP5x1zSiechDGCuj2evcOHFaA61PM
tf06W3XGCdIJctF24KBavldJQK5GwEKQJMijrBxjTdkllXqLmDDXv8Sc6JCLvuCgOLrk26dFX4GJ
Zxocr4uQCnMj4mXNKdQIje5J+Tj3E51dwpLpZB74bABMjxbFVTdCHXwiYe/Pqz+5VTQ+6jNgjCPW
EYcLRkdKCTqY+/VoH8bit44FADkVzqiXUm+u3/MXNnlPlKua2qj313Js8bJl5DsDML3dIHZO4Hm+
YQvKE73syHL2UDE7zoKiN6NJqzTB085J03OtGIYDh2XulDol7V5O0eDe9AJba9z0uvyin1gTZ8z1
Ve0PNzeL2Vw4Gg2KPbanLQ/SVGpXHMZmMCFGwQd1QJJi6cjYjfWxF72YAwuP2PNiT3N30gpczJV9
q45qnAuXJxWHedVGUMNoM4bWVc0deXwARJxBNMd+mN5Q3+Jmf1ecjKH/UG6P7Jo67ssKyAcy739k
zHGycx3NrijDvBe8IVydWbkeTcD4ww/H3Zbug5IACYi/t9by0vHkaj3zGgCFFlIF0ttnzqZZMfx9
TnBLPg3jhY2qVJOi0V7ES+Yo2y9fRuExv5QTnMZ70usjA73RDn4FQPpAZsPGkPWG1WYlr4l+3rdu
ynClrattEDTI8s/5HSuZ6oJYY7rs2oltvXDDsb7B3HDMEkuWVfn3i8g45L6bQwIR/JKsSBeZoCEe
n9Od8ff+FbEreftK4fGIjoLi4Ubsx7eBfm/29jgQ4kTE4QnUUlFSfUeR08Wk9SgGzhoJwxmPlc6/
z1GS0NSrfNqmljwxIBbORc/uohvsfoiKGOG1XX1UjAQUZcLJM6+7mbeZ0cSj51pE1h2PPevr0NHX
8Os7MQHDMFLTPEz2SjBejsI1oghThwdD8CpCPJuCQnUMz2KsOIqSqGhpqw1on9L90XJbnm3i/xdT
hlmo5Smls5u7233QUwQ0x0JdoVRXVWtgBKPzg5CPu2ug6IcQ8kWTntHwDtfpppSKnmHSsm/00qnC
u08txoPZvdv9MQWRn4Ew/BTVcNzcWOt1KWhHURML3iZ0oSjvPx8IGdikut7lDfWy1QKCvI5eHiL0
QZ8I7cvUJGxD7yExA8khh92fm789FfEeaaACB96Ss0YW6wQ73oraV1pziw2F9f1MC/K7dQoo13hM
IAar3v/zwZaUvKkTMtH8NUvvqzjgP+WceabtSKTuIecNJvPHRm8VKUZkXPelmfoLNw6MESIoiWNG
Wef6vNT/HuRaJ7KEIKNLhKHAvsHLHUmervqA2vr/IGJRSiklYo0F5qvoH/p8q0KIo+vIgdgLrQts
0BN++iLVSN4WeU31Cdelp7Ibz5tXvuW+nekqsx3SOoOyv3k0g3D9B858+CRg2CWeWwKKGH9Mvg0Y
HA+kms5czSPMZfet6NGYMLWZJ/UKyyuxKkHWxy5EsZkES+3o19szt5TNf1haxt+/uOVmOSzmVhyi
nsWquLH23K6Rz73OmyyzpYaT4GaFKmByAtDMOHGpDx3MphP7vjeeniV2pUF/W2d6NkFCwZ7fEcU/
IxwBmPLgXeNLoLWDY1yLV4SOhfB3qBTybxQi0QBsU29jZZ1J+ZlQQJqYKBoMxXeuVB38CMOQUYgQ
q/SVJKicCqmQuYJL2awMwctuYj2TzClvpvtkt91ZbXIxj8bbijPzJ0mKU0UwaWoRtWClWsK3APEp
7BC+r132qTw3NYCoCIgC0j9kklBWxE5l5yyY0qzrQS0J2A8KpqF0nqwy11tmKj2hHMUjW+6JbfTv
UClFgdYIGLYGddVi3cndV/vjkqM79+DKOBmjRONPqDQTYJhMajalPwKLKK8XNTBM2xqyvCgIFLMn
jZa2pSlJDDDDsNw3iipD1TdN0ALC1ewCsvhfrvg9z7hGsRTremmteE/Fw6gcU35rOrtkSSSzx0q9
oWiJvYuSX8d2NV8cN08jjxK/8i7AEUJwvaO9FdUtlFStq+zmPaNPYyxw3+fr1Z329ivG+t/67wZ+
9uCGzIG97HPa6EyOXhzoT9cYyAR2lpn7OqXqtFZiFQCVYry9uQ20oLONcQ6J73rWYGMmISOoaBuC
FX0v+qrF/VjI5wCxAa/VRRdow0l7KwuY79lII+DeN2Aswuoi/NylrT6mP+rLauxw2Tol6cmuvGWf
SJxO6CwBRKwMCqypG7pq2S25rWTrDb6TDUh4HKKfSVgMgBrJIMmJTmSn0YsIHMnKu4MAage4suhF
KrdVjf2UdfgBbWf/+LBm7Ni5r7azC0D3jqQdXFvaQjrIh9HyyG2tnKglMjTKq+T7cSp7Bsoigclh
bXTdlyLtKDWQPYUCqZp9i97dpi8eZy9zb9s+XBsgNomgTvXwIATPuIvB0ewHoqkikmwq9LUcpV5Y
BKL1gsPoCW23absjBohiUfpuM4Q5pjilS3Xi0Sh49N2dDuSHZuVMgbZY+CMabAWwlbmV6eYw7Pzr
MAmLGKlFKViEDU8KWVklV/Ensi1YSFuBsLbBW3A/iJx2Jonk2TpWibYl5qWT9j0M7KO9GEK/ZcTl
nJ1NELlhMw6HbkrvKxNzOIdJRwGuvfT37+YD+c98e6WAUomM/G5HzXyR2viTuVBlKQJvPXP6h7fm
BpW0cLm5IXsfV/5LkNf6785uzLL408klkW2RZUhEi8YxisnpRGqEGqlhd4/fcN7EsLxRbgVboisT
EmwwZijDfHDfYhWqFtdcGCu0niidQDBrzNtQJEFP/Ov5CZVc2qmMhEdAo/APEkq5yb9EXBoiheLZ
d1hn/Mm2ocecyMz9G4XSGn/WJi3tPs8qasxDn/vHNlNM/+kNckVV9vWeHcSBDC9vtKKXJZ1m2Jmk
LWSnsEtmSOb9sIq7YpdizFBH4mrjPl/WhfmybIzp/zIAKS1JXyIDhRmQbsIvDUctY7FK33v1F5mc
DYTAIrc5WoeetoYL73CQgSHLve4xLE540j51DScm6vyWcN6+0S+p1eslc7W5ZKna/Dma3T7TBQ5h
UUXKpkMW+N9F9qt+2GGNFeOMDCJNmjMtwEtcGA7KJNsInRbSesgsllhzoDO6zgqUqrOcEWLisgxK
7QydyvSe17JKiyDRdben8KEb+UlPxrrrwQ244PFVM9meelCbtgJygz+Er+oECTdHq4f+m9krwZPP
jeQQbcBaB7VzmlUWv2/CeF5g+lT6NX1iS7QDRWHaBErNvkeum2i+c36zGxlw1XNpLLVcA44fBQCw
TczQlIc4uqNGkvs2+ggzKg9feEDQ60UPL2ufDgVO83vQMm8uRzb4+BDOg3gZxsO4a91vbETCjrE0
FeSSvQZX//qlv5zaQ/9ya8Xy/G5wsiQ0GmsZSRtwALbcUozvzMFLTr4Lm/U2pCsDAatO/zMJ10V4
rDWp9Z+a9sggtJuUBeQN0ezJDmy4QdeXUtB1v8RvreX7iRuDgZdgZ8RDdp/WTKEn0ZfyVOPYiF4b
pNYXCtRKiMfKLjmtc2byd/XhTzqoQ/W6TwPkvY/i1AYK0uR8Lre819HQdnsviN2QiJ947a04OPDv
QivIWfbpmArqFeD17KmzB3rthzJWptCQsx4xZW+0yEwtlIi1gtCo6PTpfB5e82bvqAw1nXu8KNdz
Ugl1h+BbPQf8P+0iABi/Ab40rGYAI+nmUyQqnqLj+7tsal9u2Uazf2S19YZtLH3OGfjHhLZEQv+N
UhVklXF6tjoDJFUqpOxfUXE4lkF2xZRYfzDdLkdJvGFHUWinv9oDteecnf8TTaNrk7tXuId8djcY
c1CdFU+Zp7uKoIOG7a4LynfMLlKXSBYy/+IanCF0diEt7VPICymbbUOqNWoINeWgIhc6vFkr+tYA
9nE7rKu8WgSTANzYGu7hCzdbimzp/5ZAM/ZsEC43vEU67+jXVP5JrMUahKArbMXlmVXjTWDLoFA7
jQqdckdFn6UoUYaUFW6cyzXdGF9FeMWwOlNXQt5xa5dEWBFmb6Me507UfNWYgnTJMEREl9oLp+9x
8MH2NIYc3WCOtx+74LMy0q54LSOkRdpR5Nufg1sB69U+BlKoJjj1DG6pBZ2Pqcjej7+GYoHrVHH4
w3yXnlS0cf06tMVnPOjEIJsRa68sSaKkecaAOFl0YZSPcKz+1QdbTjnxUFshZQqdRetUxDwvTrwi
h8hVCd/3NZ2g697/sngd5f9AtRySDvxo9CRPwPZvXWHv2+xRgC7VTME2t2NzRKyCiaIWdqcCFO3+
f6P72WRY8SltN0ZMmDdacntP/jjlbTCWqzkFcT+Y9+F3QQ60Gq//aIbz6ZI8RFXq0Gp98y5QvHNa
7MoM4YZ0DCY2HLblh5SSKWumKYdOvxIyn/9xg8HUMmrvBiZK/Q+KCMTL/VFFfbrJ4KaM7+MP9kBx
+G+mNYmQBO6ufsalQd6jHCG6LLkHIOYhaRBWGvLiNkMmNEPA8lL5+Owyb/d8G3u9VYfIdzKTx672
bHKjH8lphmvvGS2KE2jukHudOCS0uljlAdBW/t0fgBGG6/HMAo9FOIGOIjZQf1zA7708mnEdWi9X
aDo9EAk5/aOwVvB1LacuUjtgwOjMMzxKNn8+XaoRF/+SS90PEyF3sftlEfeqftOdw4pi5mPITykI
63+Bt8tYXPS/qBevmBkjVBdYlnWyw2qdZLchlFKYvj9XyhCtESPA5+daT8+2/MRDeGDONKwnvUzJ
kmMdIILsiYT9bjdtbb2X0d6nJiQMrJ7HtcaEwYn7OagDwi8h9Fu7RxpnFK4gVfFLzusSPleqpcql
Gp9lTN+P0g/lc3+yQaf6nJq00O3BEYNqf/So1X1OS/D0my+r7zt9NPqi/ymWN2FX60QZa6TSTX1w
r04ftp4UpFQJT1QHJfojzb6xRaIF6KDaeR7YhP+S9pLZ/wrSGRXKGm5qQKzopsiQ3zNgeGpaZqeQ
nE2+r550CkDGsc1ITmvEG26HLx2mdG8OKCJ6JOxPHmaIkkkBtaKOsfR+RVqFjvD05WBuclGhmmwy
mP+nK567PQMVbdxFY+CnrkYGwLBwofEfTe14Qn1QLNjZFxGh9avQib9wXayOTDmWOq8VGz4P2XxI
dN31uHdzQwPrhfYluMC7WgfIsCBCL1jETAUByc814dE6VqHVuAa94PCmKCU2cP/2jnScdphrq3Tb
EjTEVY1MIh1Ic6GLPd8437ne0RsZLm33Ia8DZ0kb0k9FM7pjro5G3TyLMVMjQK5ybDBhnQKvDhoN
KCWJ7KDd5zdQZO3d7WiMb5M3eCzriapULQpyaxOt/psvPuH0tyUX2H7/++678oe0kYZvCmzuFeZr
sNYF3P3im/HMD9UUZm1Z9w9zeKwvGL33FVjmz7tydXAe2sRLe1hoh5KOY3ctCPvIIMuXoP6LPtSw
EthBXryWf9S2ujuYs6QJYSQS0htEzA0clfH854s/jFakCT7/zWHnffxheQTlxwg+g5CDW2EPkfe6
0aX+yVoG5FzCel17hk2Kmg0CkF2gki1xW95SZ/7iCzRwH/vJMaFKCQluirY+1K0PtAW+aI6/XmqZ
BGmADkMEND/Z7H1IEmSv0J56VBATfNVBireBRVZCVHgtNrlP/EPQ4FHW1hE7OJiVxzoo+nj38bCE
zypmfFwmDBejNrhD7A+U5D4RUvL3+HjLLa7BZgFxYbGJ3hdLjRSooquzHp2s559fbRe1G+hel9uq
yEhedAA+nOrVP+32kfl3QAToJtfUNmfv0ykrecnZNctfZcSFKI4lAJqzH6xaMWuR6Sl0XE8OANvR
UUNwzUAc2N0tdhvAiv6/0wWcxJoXEcuKGO/hmEU75pVu1sYRCOmxu9p2JAJnewuRBBuPGTfNS3FH
BOgl5Z0NRYobNj7E7AnRTmwrB9Z9tP24KNfJ0hYoKoWDf1dv8+DwW9GXVkrGqlLXiYIMv16xPicd
lMQeEFGcGnK4XsW2wBDNZBCxDJgNCP/UsAh/LsAP4mMi45xjjTBLydYa1lF72nj4b1560pypWsjS
PyhYRHj7mIpV+DUf1ZXHcxQKYoq0rjBwCSVbRDbPgkb7C6lIsRcdmFddxg/ZpP6jiMcijkOfp74S
NMgahWFpGyE9HZBaUvcmuF5j4RbBBNGd2I9uAu1AZduiKbwY/8u9XRq/3NsVtdLnG6Ubmf581+0f
rc3sd/iStVG+C0C0ESmPImVM+OfQk8u+eqM3+8MtKnPvoROXM6FHXQb7UoR1PtntmA9WWhfD1xEm
AWyJQ8mf/4a9spVx0N5+I9uCUAs2Fd4z4L0/2tAt0IsfLCjLpn2uvnYB0NQUbRiqAGMOLhW7cVno
BH4VBrRIRJ0i+95IX+1mcb1+f3zygqeq5d4cQe3Vv0GAirTMHO3TnKaXUUW1+kXbKtilma6HhYnk
7zIDzfkihPgVMOQsh2+m4NXMaSweLNSjzoo57WDL/1K2Z0a6c217oB4Soy0Qo07YOLapOKHEym12
CShfwxYWpVHMSIXhQxrwx5innbU5CWkv5Rg8VFSuWNFBB1aZy7ZuNbmlBjTtCB8i+fDajjpi1wX2
FStC84kBqyWhjGXrcscooAKyo86Ru0jOEROOvGc3wAUureXfVnIRe0Gw7sVtW9iuuQEu5Lhu21pV
NjmqWeRA9ikR6z3FkgeN7xGcRDRk53rzraVi/TsJpGeIrOPHGl+W3dO5xfiExx6LgDUc7zsX1Hmu
CHiIhL7WDr2z+4qGgMZrwKeq5QqMHXP+sMAWL7ZY5QOei4A3vUIKiBRyj+fGLgHWndffhSgl4YaW
7ZPwOAtCTLQolNhN5yasjTQT6klolgopoVbEHG6muE83ccKWtcNJiUzI/MWeXBKDel3Gsuy/rE24
fWJCiS2qfoVl40nfOBa0IhJLue71dm8FOAU/vSmQArpUvsVQFvzWJnmyg3omCVT5wDz8DFpc+6Gq
N2copA4anDFpUVTGv1or2hMGPMiCbIiFps0fpgEPo+riHSS9l4SjRyIt4HN6Fndn/dEvdo4s5CLG
ukaDPJoSJFwMrohHVtpS4g4uEGq7FnTvd9aR5hm2H5ghsrFZJwAE70Zney34cffdFYvMmNmP/OOX
ocgJvKqVzJQn+e1vOBTwng/UU5HLHig0Xfk4nenyq0OlCt8vba15uVEwGEkP8FLiBv2PFLmuKZxH
e4Ca78op8q0EEHy8E9e7vZC236H6D2nipssCBUIcMsxMmKWtjYDwPt+DNdakFQe8na4bCF1ixcWH
gbBxKzckB4aGcN3DPRYN9iqtMeHJT0IMSxL2frR7hdSO7FCy+byb0cPwMThmR0jgtjxQUwAmSD4C
7meAuaHAWNnwmDVpUL0DR4t5jLVGzJBviV8tkMdWHXfu2xTLgabfYh45deyjcqnHesMmGdUXdKTK
SdUOmWGzzMYroDURCCsYPv8jwBSaHUDfjvXoNoJKYGILn6Pjq+jiZDClHCfkLNoUAi8jptE8tZm3
/pRRUfes7I7U4ucg5ozauXFPI/C8YWvZeDtHlkpGgkeL1LfwL2elnwxIt7CwQ5E/DyBP1Z4urKM+
kWf9NnwjrbpeiRSdpKYxqNAaWzTtKKKsRmjTwJeZKBnV6jHMvOG9u6JPfChXdpuDnVxHMHs+7uW2
GcS99NFtIlkuu109/obyGQKMU7C+IXjPGoMThwH5mwDp1758DhRYE4b9JqpdRhh1WfflFAb3OJ0P
dVV5iNPfEdy2Q6TXaMG+bODR/Cr5s6F/dLVVCLLOpz199yp6q0tjK60smw/7AZosOZsjWVQpzBSe
4EjoxtxP31HZaALNkepM+8RWIbm66rVEi7ZBxLS5XIzcJluRPAZNI/3D6EEt78ZfN3lr6c3N0YIh
OzYkYolKvED1V4F8xVQI03DGuqoAIquzZOPkP8EarwmuNYC38FjRWQDcjQ3LZnT8c2Ee1z3vAoMr
pDDxwp1QusDiDAZAuDqy3elnJtZWz+CGgQFsmRMdE2I7SkGG2iPTFt0q1AhDrDxxq0t7sKClkLZU
+71HeNTHTV6lM1u1mvdDuQkxs2N6HDiy32Qwj7DWQUQCGk41EvnBAzx4mg+OfOHWnp8S5WPlQzrg
cM/m5i2VpKJM5UY2A/J0hrcXwLWdEy5vh/E1FVQKGEHVgJEjG0YxK5D8UAtmncJiLTVaGQTvVzjq
sZQi3488nvaft7tTfgZtxelS2ErRAXlFrC4//UFuJRfPCSv6D5lnTsh765KxbKs1Tiebnae2S1fJ
Yv5UkvRoQBb9/lRWigJ0YI26vhQ0pLYepMr424mMJqdJ+A7eOJdoIg3JX0z3t5rHgYRDn1QWBPJC
fq8kdiQJW3ieN3l7Cm5/yvHXHHnfMfCEA1hdxw+1lgTA/hkzmOyAcXGyDfPhCjV6l5/eXqoMa9/6
1bOmQrmmzQjLj7iWbqROe4+pzSu8qZ7wKr6GWlvQmXhCP7INEtk8Qr71XgBLw7RkJUMdmmxI4v9Z
SIsKBCKzsz/uhSm6ib3q+vwSnkMzIHCOz9mWgGx/hb+UwxdOiF1DY85hyABznSqLPKDkWl9g5Qgg
GpQLTDtOw1D6JIwc32W0S9tb1JhRwtPeH/sDwXLMgLvMPRf64j0cmfvwCveBbbszftq1tF+vWgUK
NcOnSVB899YSYQtXXBXIvL0HdSCChTt9shyFsuVfxxrCUDQX2ept9EQB/OwQmCt+VoZJ/z94l3j1
Mrj8Vw/47e9mrSYaP9Y2ETB9AtXFL6xLL/2+hQcNnd1Hwn2oKCZJOGx/8epB/BN2t3b62fJGJz06
QD+fjLNO7Hmy3M/O9RmoNfTX5jovv8XLtKmBt+XNB3BYtkFdFG8rVN25j+Ro7ZxXM+XHO0YXg7L8
ZYw5CnbqWXQbn1EnGL3KITvbTwww6l/mN+hJy5trUfRFS0Z11GP3/xodXrVgKWV2pkQyRL8I76E9
DrPydNf/uiStmSU9kYkuKsfxUFRt9weyggRD4vEGUC7vCTFwEQjXzuTspScfkbyLxdZckqSu4PEZ
zdEfCgm7LUNBLsMgAsd/AOJCM3lXrUKT40mUwBVoBmdxwKTdOYYSoMFuNvaTXIe7DKDrU6WvaDOa
qTDqsyinZkQBaILsgkEGhbo2pblKHERt70nVG5FLOWXkRxy8/2D5jQs5QPr9eBIT+Nmr96l3xQGQ
+VYZZRhZvZfzXhZzZ4ETIHswtIGe7i4uTN0g566zbDuVHBwNX3Rhe7xm24m6bZbIo1K4B7CwgQlY
Thvp4IxRMJh2wLa3AnosJblFvb1lQDVktlZg1biII5plvuosYyTgGuA5td8VD2swedRVx01r1DH2
5d0wBHonhLBC5TcD113iL9LJALTF7MPqQXVxoXUWK/LrgTQsZOOgrzKlWgwLyXvIcnQxVq5pEqaG
8qwi55gVUcKqpcT6tLveJXBQb/JX2R2EJWJa0OSLvdIL8W5y31FoB9oybpnuNMCIi/Aip537ttsM
2OOD+HLklhFVlI1ciXhZW09F+LUN2NHBLAC1d3DnXJod2xFXAXPeh+Ya+RCgCQlBXmEk6RO279rK
16S8vLYeDVntZK75nONjyiWmeS30+1mO37OLkJUPjFrdnv+5yZJQ/qPsx1YSuKAqvrCesGUGGIAa
3CqeHwXT0QwHgjat66f0cxtRYiGqYuOT5/Hm7bDp/xtEaUEFnauayTb9ji5d1j3DbRQ6LXhICXjy
qeWiBAT+GWrlI8vKPwfPwK9ANKsSUNhI3K5PKJ339CalebsR5owNXDR/IZeHgphkb6bksancmEM4
VI6moeRW8tZDBj+0dTX+uVNSzzI9LDzJn3OxXUoIHCh4rnakXchdHEc4AbtevGgWn098g5A+0/R9
fV562ao726+9f4DHfixVK1e+zs/LCBS+o038N9rVBn8uYsjresaohAOumQo4SOrsf36MktZ7tihu
0Sv2Rrn4e723NNoNVNc3y2VFZId4toxPOO+bXcxy+n/nABd24ZY8P9Zpwg4MbT3D0HcBx/0zmH5t
TDl66fplmHxOSXqyoADVAx6iUVLR4BQR8Zs2suaRux+hX/+hkSk/dHaAMft0gBSqClsNM/0Aof9q
x5pnskZ4AGa4SAtG+tdrZwND2aFKnzQP1OVYnQloqD3KcZT/nUD6NHzUxU0+UWqrqHGNfAoU0Bn+
1isG9U5GOmSSn3fM9y+sNZV0jAq7+/tWhsR7pVFnueTmWVhfrBQxLNXvbVWlw+mqPwspVUBQdJI5
HKQhM+fmkb3udOHnLnGmSiYjwZHGlvtbSrJ8mhkyrAtt36OwCjdPnHxOJLQS8R+PkZJJgeiCaY6V
JQ+/kH0PebxgklP3Z/5UNe9hz1JhWGG/sprWn8YxamJ1vgTCBe46++cOVH+y+naMLaO3SM4FGbRT
bte/9Xsu+ig9tQ4X1omEintG+V6y0o2wy9Q9DgKkSybeFy+EGkX6RM0z9sZj3zhW1/VJgaLO2KMZ
FakrhzzRQ0TvIgJz+H/ZYwHu4dg7JTHHWlLkbIfvG513d9K9vZerq5p/s/djyY4fXIjbEaVfK2sV
P2NWql+CCr6Hymf246/vnA2ja8mMnIc9SzeS/4EInnXT4fsjHLdG6CMA/D03gA6N+bUsfYXGSgb3
Ej6jXXcdrdjXUJDoFqcDi5NhfDle4qntkDdBn2pKpuLMb1jtEfWeAHFQ5JvBeWyTBixEQpftP4z9
ZMytNukNycFSxBNxbGqTc6Xdtgm+MCRgaX8M5JqIOsXtW1Baeai4xDgPPBxUhIdk0GdkPTFcvDw4
2Aa8EvEW2HOhH2NgqVorikOswp9mkXt4aBJpgir602gZxNp17ziZBEU6fHxEseN/TLnj7PqHdjmL
Zf16y7/HFK+axMB9x7wLSYgXA10NPeaEtMfq7kJIz22681QYoAft+OMbkzj2hHwZqBLymaswCvYk
NkzvE3hydx1L0s8LMwWZKPPD939yk59aGvbh727VjwE8eoOd91XuisBOlc6pEeQxDrPPJwcHDYNk
PhNdLqr6I7vYVHSUc5TKlJAb5AHJz9BdPWZhAt7FlbaNGzuKu8s0GhwkrnGAvPwb9SrmItTeyhHZ
OTg8o0M3ADwsyhDdB+D7BSKTio/oTlTI1VtzCJTSrNAjcHCgsj2twPcAyOkvZo3gCZBSpaR04mME
zAAyRGg2Cq9QBB2crrWBvRgmeHM2IR4++FHa12nCnmpXuk1HmZyhYg9f9Tdaqfn2JQOXz36Rf65M
tWMmssBoiOWoDxYQunGxZNWYqXT9FJIaJ5CMiG+HEpss+vRrtpcxt0D25Iv6lSUq8Si5CpywddWV
zBGPv7vS7pPtH6c9yTJrIslp4tBm3pTG6qhYl6Cj5Jz96rT8q4w57X0ZnsqPIi89qETu3+x8fUIk
RVDiqqWHGuLIovsRcVnHWZkNDbKif3aCFxPE6pASWlGJxPCX/b4J9Hl8zIDR2yo7U1oPkmLn2pTd
cg7OaYln/hcDZnGUow2RBMEp9ge8NU7ra2DuKDPNr0P75w0BDtf8VUipnhiFOacZylvp+mzsgYNN
edfLqmgQwXRQz24NZI0IYt8xdZc8+FVHSZJqHPUFoBzaCZ6lV7PFsr5bcbIQxK+yeQ2B8hRvzYPS
/8eS7tMqt1OfGMLCGkX4NCmR34jaXL441NoDXSFtA9G20iKk4v6J56KCVyAh5yJM4lZxRYiZL0Pk
oJo6b/HcG6oBYuEKKDEdLS2e3xHnvoFyIxg8bQa+ZjpD2fpQMo0D45+DyKm5w6EFmMQo0ZB1HI/u
yP9CWG3LKez2+rCbkitWkb2HCqsMrN3DXJM+tiWSFdqyI/V/kSB1spb2IYnFJOZD7MzXEIbS3Axg
xT5/rGo0QA9AUz9DUohhzrp0IrjvJxFrDUPPaBoOKJAFBXgXiiO8m+TXFvmFv9jWIBeAta9woBo2
EWz2fdyOzrQjmvQRIqBDWkQR2fdDe4U77IRLjOoYu3p6jH2t7JC1Xf/BwZ8IzOQUEIejMIzot3z2
xxN4exJ7MkYv2tx6e70OUpU6UUwFyfhigNEccvDS+M1rrwV7Usp63noW28FNadxbv/n9xVM7rTTA
2L0+jlat/cbO+XIYo/35wRIxmvwMIsAbbnR9PQ7WcVfT8VEfcZJGonlc+s4QFbF+kJBi7mLk1Cu4
mEOvmBUsG7njQGsFxS0U1OYxJMEne24U8QinaZq8NlgRjhYkNwIY8iRfGZvhd6Ka8oYDIK84vWJr
EcmTbqPnCGbwJIJEqusi6JUX4XpMMtIHo/OIVBUCJpcW44BGxKi/ER9Mf3pD+Bll6D6AAsswYvXR
LoVzLets3oQAdcj5WKQH9A2QsQzOd2MaUcy7gGbdUq9QgXNcRzDAuxppBHJXsEJTz0a861RnmCVl
LFM1O5BwypUJQaC6X9xgg/tdMuZQBhrLPX1N9bmgHSKFXZMYOTn5FyP1OIZQ+RnzoUBBvpXXA0XY
Qr5+2tTyyGT5XJhHlgqI62fzPXvf5VoTplehxo2/UIiGVmF/DI87BOBAcj8+CiQ0NOssW54I0ReU
7Qi7ETSKxoDXC0sZjQuMQpt0lWnjYWycRkwYI2Z5KIwsjBnUmWfrLgskeQhTaohbSkrYU0L8zcN5
6sCCycOO5Y2kir/MZrF35dXtxXJp5H31nazbMLlszro61Vv/UiKfDvYhBxThiH0SEU6FbkuMdSiD
oQLpNIgcqGjlS7Ts44VfqgQchgP9Zvad/4yRbd6HLNInI7+LWOVX3NtoGzd/K2k1YioN1muyBMGP
L/QJt1MjFKceQh7SiAOzk00Ah+OFrrY7wOdECZAS8q6+MlEeghFTRPLPLexH5K/GTp48GaLMmCIr
VJ/V2gxbRg5uuv7J8tJuHeTvFhtYOBMOHUDHPymXh0QrP1CVv+Qlh0wKfX9YVQS6apirzMnzx/cI
BAiVIliXzzTDxToRBNHuTWJUJR0QZg6wa4dhzgaiswunV3n9MBY+hS4mKacMoco9pSkKlCoXzqVG
Y1sQ55pMnrJpChYVc3ySOZZjsdxulXMDCOxuS9ylQvvC36+MAXeDhu2c6YBLBgtaiafyNbLoeXa9
CHEI3G7dGlY+OuQCEa88kYHzqZKdTdGDCmaj8xh5Vi9Jrk4uQPTTYE+ilPXg2RrbOLA0UTMT9qO5
GI05JXHEwafCP/hSX59x/Dw51qlxN5dw4pT5adz/o+afAnc/7dB4AG/i8GBIBL/WnDKYcHXyDz28
dqY/3GZc1fppMVAQx8WMvaOtAJqeDRBKKNg12MHh72e9UHULsO1dfHMVP6GrKe9eZIlfQ6RIBDj1
hC5ITQWVFyUEvJKwh5nfddFkdmI2NZNWzg+HfM+VdnFeTguCp6J6AhlqvZ8g1P7TSlMv/5uaLn7w
TzYcDYJ6oPVoQL8gRJABYwwO3tlt4kqRy65eG55uQDtxU+12/b0xPVJOrY/MWRNgProd4TA69FFh
Uhv/GHmQFazD6TvE1BVrm9wTwCQMlq2s5FPcASgGmeYi7gAO1bPfY7TE4FbLAY2FadXuXZg5iyu+
ayXWxXxz1o9uEPWZtzVr6ZBkQUVLaTevLeampwyh1WyT1GsN3ZlcUbFS7seTkR3V01tuBrgWbEs8
CTFKAr+pMN0JUUlab+VMOVASILyQZuphB/p/gbm4ZGTsCoLGa2jR0HxZCPupaolWGTJqjKbwtkH4
O2et0P93uolLU5/2FEo8mD1m6te9SBn8gs0BCFcO4MLdlaRg9ztRN8bXxiIb3iB0fsiLBE3oWb2T
TS6Y45obeNdrXygywzxOJIBmy+384IiDINxdxrO4Gzlk2fIPpRNCYBT+Kd4ka6GAQgbyuQRjWUcP
OwYnMrba0fTSpSprt+OxAkmOhm0Zwl0ktO5djr7DNF3YD4ViUT8/oOSiNQURO/DklW/6PqkFx9i4
7wRjYf2ZwZePe6rJoXhutbQCjzZUvqxXujmsm+7So5R8bLp7eR7Zu/vRMvmu5hnqe4Ll6JRM3hmM
O1a2W/8JjvkyfmpRk4jJYJj8t9ROI67glOTsE+cPLphZVJTeAmtFTpnAyA8iRSSyUobgAYYdMGlV
CPDZ1k/Wp5JA1ffAK8H/18ZUwQHEn9PMvQCVRg6SODVUyfa7cI5hFYrLp4AdIVSIbpMX1itv1LlH
UY1Tn43JePjg/DUI3TRAm8ypvbf2R3nlj+FsC3L7IFJloqSOWeyHw2mD3qpn05Vyz8Wm35aLhD6r
50XM/9PjRSJLak9Tfr33MxaZ0XziSaPuZdI2acACbWgf5t357EhqRKz/iRjgxTl4E3Pxz+k1gbdO
8M5kIaxsPHTBYh/97k3WVfkf6FWBntZyLlL9E0NrGSNVOoe4nCl4uG9TdyY38ue2kXs/vWGYR557
nxDEmRi78UEMwtKLwt+xHEHlBnhTySZElAzHCytEKLSpM2HzIFPaXkkzl739FAyr4oDfVE3YlAMb
hrixPykhkyLiTaIur+3fitQ0g9GEH6eue+vP8RpidjAScVrQdCD5MtQBkY0KhVLOWxTl2DUtETPO
rVwkDlXrQqW+Q+Vv8YJX/BbL5goRkxdufmKRFA5628QzuiHLUUwC9dHY558N7lnfdrTRY9P5CfZO
CidB9QaAOpsVGBn3GzZH/IkvT9y7n3G9hWyF7w6yk708oFnbbQvbTvT1VWG8yHsHQBOK6AMRmr1V
ofLrj9VUr2s5ZJGeNRmbhLT3wdd/dtLg+TQwoSpzdgvPmfVHKhUIlRdsnZQtbM3WJPeswI33TpX7
RQjmTLJferUSSG4uXaJGn3zFAWdhadE77uLCfcoPFKdapdNVy4vCzcuqe3vaqb1cXoMSmLOIBUSz
ovIIUu5VJFdjLFBROaO8/I2zIvkLlt0lc5MWgHxrTd53hmwFbeEEVOZmyVHlNYBE0LWHT1x1OUB4
H4Bki/HXgzrlTI2Jspa3vCe84/CUuTTwmAuTHnhEe1ibeJPSQ/3jxGk6vVoD1el3f6zBL9IgYp9W
rgzV4BSqSfx+sptZhWFDzNDSpZztxw4TW9qehEZ8GVfRBLSwVgkHpTrvZyK14rkNRUiogl8udhZR
q75FAyuOvPeY9ycz9LMAuVpWtJ6tX5oXcU3/2DVtycp/fmd22lhTeND+Yb1E5hAliRUERC6OC1+7
b6VSDpGmDXyS0XQxkdVhwjSNotTOE8x4iB78n0Pee/q+7D61aXYgbE7WXgsNKqc1KvHsOYPRj2ru
IFmBy7N1duzCUs9Y6E2ThxmpLSLiTJw5Vxa+y4Jh/PFNWWBSwoSxmSX+w2KX5ORL2D3gzbv/g0qz
zXQuoRys38628uBHSBQmx+LuYFI1iuf9ARXSKQmhyxawSMcBkcxv1e91UdqjgBMpQCIFYFXMe75C
dPOnjMClivXqP7/i32rYdhOiPcZm4A69XnEeEDd7bzDbApZ4/coSLk0Fs/miFLQSWGSl1+xEZhOw
j7iWnMOolDIwu+jUfiCptX7B5pbU0wbTv0DYEbwN7LQdiYPnTVhEr14ID9dZthf/Hd/SgeGwVhkw
78Pt3V5xJ8ugR13/U60hLQzlQfCxOgjn3AHqu6P7Hz0ln/Qja9fTjggsBUgGgnlQUcsR7vJIGOlv
dWiMBB4dyf5RvU3EOPPo6G4QoBA1W/VihV8mO3/ldoM4KY2ws8kZ4luA/CnhXTZ6btN3+Oi0RU7B
GSN6mIlI3ryJpn/AvxiIrm/SuSC8vblS2K/VGF5Rz4OuMtLb+WnUwXjlyctQYfhDKzqVzmJqfoKU
EUuUQMz3Iswdkc2XH0nsdTVs9z3DeXfAJpsdezGc9Dh0VmKhfcj2CG0RmSLiNjMLw1hsky4cin++
BqkwSM2qZW3KWTpKeUhzKeUjeQqCT6LFnpj4y8a19o0dn8/iiXbn8xW1j3PQ1ZjbeO+MuARaF68L
8yS5ho38IcxWimQ3Glbf8KkRYP0eAfhixYd/AFERFwwvc7PqnxaISn7WihW8RdhtdZAc4RQcenOc
PBNE5+1iB/gEswdp+N8uVasUD4f/6mChRFqihTVcQMfk8rGXy7dauJCXFUXAkKgBCpRo17WKutv3
XEuxHxR+yw5PrsJ+c5TMNqTtyNPa+CbmfYyx06T3nMZ4fZyjipHUKm3Q+O7JVGBkCT9AixHmbcpw
bQb2TWllRUuKOpiZJAPj2XNrpzN/9MGjH6P4q/umdNLQf+zBxgaOef75s9vRxRxUBYFtrX4ZsXan
U0P8zsHWB7hE+D3E5qxsY7cE4QUOC9pvu2hOTHble30a1upaVsax0jLjDAyAugXSVvS+PfZS2te3
lK3cTSE7bjRk+JVT3zNgUPxa2uBz6UiD3GJZcCDehhL4z7/qUKXdXyfOWryk59wDD4BkfisefPIQ
BRxResDGBNLXmIAkQmLs9i42Li87v175kUXOCHe7n98sm+6xH+Uh0fUz3SK/EpSOuKObcDo1v1Zm
X9P8DN86wr+zi89x3fXlLtjyACyEYcjmPVYGMVSVih7aIVS9slocrTSFHiynsC22y6/BoCG+AQOQ
IzE9RiYVI6dNwaZ2qr8tAEmlpqR/SMLrqHWV77YL01KILikn16BV0/DZ2UgHjcbZNlm48LFuzL3s
FaF7qacqA7XIatZfAZAY2iuYp+rfK1ZE43spGKv6M7Gjb6sJ2RvWGH1GOXUzbGOOJ39GRorjvAEU
VGCsBfexz8K8Sr1o85ydMc+2DCdD+dPT1lSKZlCRNrcI3onuQVy6e7yWNrOzq5L+VtyN9v56nCqW
w1rAFwYeM0lQG3tvJqrg0SeO/+UMVR1CnartSYwQGI6cIf8pkRhnqJXxTriLanOnR7wOaIIF+g0+
D0Pjtyg2xqw9re5TlWrjVYnhEG3KOHKRXoEt2pe92a5c0wLlmGv9+lt6eBC+aOq/X2DXEex1TSdn
fKWdC2oGNb4s+6eZ3sXYjl+cdEq8Xufs+LJ4APPszXM4Jvk9NhIcSmVR5RC7+5YstYpC5vTzN2bd
yxblE9M+/8JPddva6tSus+ExDRXruqeAbom+oHEqDT0QTbCixMmpmONr/zMaYvm24p6NV0Pzq+1E
NUWLpKCV+qVRKJ5kSmQ5eEPbt9+fcfWoJ1qRLd7+eFXsuHadOS1JG9Hg9lL5KeBC8YB83OeiuWzI
8fEyNfvsgFtMKh/CZ1rNQH9MHvrzKBPn5+n7aCQJkfEaLNzw+V/KpdrQhrxFVUnqJ3ZKEUOQdUAU
9egaYPh/R8FNWH9feOUVteyUpgNXwnA5XhBsnlmBx1ag61ytoJmTYbNDGudLxbQsvoEHn5zEnpq7
JIUkN0X8jorUUGGogMmptbtW03NS7ztdeelhdCnJo9qdLArf1Dsm5735yPVmocnCicprEZSOwXue
l77aKP/k4I83oio+P5jb4rEtAO4kncmSis9MD9DgbIzi1v5MUqb9lvhE5fyiJoRRU7BaMkiTSjX/
BTPZsmhCSOPxXDspjpoKo8pRDvjBQJa7J0VwoVZ5m0B3ofA/xRGS2EEUJUapwLV7GAIK50EMSl8G
Zs79QWMi/L2ogI5g+Glhp3WawYyzH5RBil1unB6H70I2JS3Yet9MiizKgVaU9oLXxHUprHdlOERa
LMPpjqsLwKSzkwCO6yAu3d7hdB2DLDbq0MKAp65WgKwB/hiqk1wQYdCa4GBIEoJpEpIW71o7zSzX
QlIG0VzhB6QR83oRpM0q+doeupKVE2fUhUh26lnV/iK038LtB1DknddKfQOivokC2hO8O2znuKXu
aA9FrFXslt32OubdssNSy+fMexsfYOwuERcJ5xMhory3FkjM66pNKAJ/LqWaGv0cPhgx/NIAN4og
viQGFgXxjanxHhaL86w+8gtqjRlFVuYvTGOk0Jyfw+RYF1bjycrQBnaCL84ZSLHPfP3eJm2OtyG7
A5hr/axlZAH2fdKeSwwgQkeM/jV6WQRtwsAKAdT2inrd7UcchcL75SOwj0a4Snq1ahI2iR/nVF8F
ThcCGmSahJ8oN0fGAEqu3EKG0sSV70Pl/k2GTFwoEAEPhSXodq51hNQI2QJQv2T68+LPvfBOT4lF
jSUhlTtGtpJkJNl/hRSKM6EikeDdx1Jm0y33ln7BDW2J8ZDlL93G4uCGgNPh/AaRSJxTe+pzTMth
ikuMXYcwjY7UAfUsSAcw7r+rlszL6JYN099fmmRfToBDZNJlwyAEwgRjLEtbsdD3F1VyJkW4yUwk
x551dsKvjpRuCilt3njLSvR0YVAREQB/fK0jZPSjks3e2kL59Xw4Px9nt39xdtIT+NauDwhmBl4J
Q9/xUckj2hrAD1iBuD+f2wOi58jCnt07hqwyUeP3Mucvnx0iOH4vkeb2pn0evY7IDLOj+Zq5vf5O
FjCxvh4fLA/GbHSfLaXhxLJsNC0Yh0F8U4Kv5LIRnVTKBDjciikZSF24+rqUUEzTrXXN3spTimu6
I/zEuyn0/hIX+rvp1fDql8/HMSPlGq6vTklv6SiDSIns6ACktJLOYvgmdALjN+zQ5ELrK55sP9Lv
R4/RLnyj6u2SLlz2QV2Wu+0SHqIffNeoP3Avi4oc/RqSoE5qbpLrVoFIU3aKpoiw1csfxBbwNN21
lvpZUyuQkSsZq2Zi8jHJSFKwRxPsToFcIiFqZfQkvbKWSCuKTvZXZMd8/F+QRmxxeSS4crSdmVFr
ipw85nZEoHU2fK8F50qqwOMKoBHhBP5rNfNk8j4EGzz9y1BttDSm6bKds6VrFX3zzqmggqpkQbLm
eTYlGgwZ92vXEvaykgJjzcOBrFo1tZmmP1m5XzqcJxHZxT0DcNi7uUaoMC01QE3hlM+Lmow/LKRf
PxyoU4Y3UXFYc+3DctqH97OeqFY+n0ahLL2P18xvTxW9A9uwkNS1t/g00l/Fd/a9CG0x88R1h9sC
5GP0lu9SBfQJcflVGjjR5qjILfSV8svrpmYH64BWjc+4avMGzImjX3QEH5SHIFE5gAU+zH33lMJX
e3YhFJ/BUatx2IAHKBQOuRyWhgxeysagjaq2G2kYqJ7XQthF2vjUMjFV674mdxBWdmSkjreiF2Bc
cLm8Gu8LKwd9bLlUT3qf4AMF6zNlgkcwEi7U0lfBYgdZ5xXC1xzAFD2b1cZPHHLVEj4dUYFua7cn
Bt/mLERv5B+iCl1nq4k0TToDM7wg4u8X8xgv285ZwUaMj+7PFHC7QRkEd3ZciH4e0WxM4xoNMsYY
RawjdDlZ8BC0h1LnMNLeaFVD5/dP92+goKqJy5eqQfnwsKoLXyZVYfcduTN61eKFueoI/RivIOaS
qQfcDi7o53vaPM8qq0KmBMrs+wEr5Ja5PiXlGWt+wuPu99m+yWeNUEBnQaTYohP1NzRAMb8PjZw0
+NFNw8BHvSV8VgJFbh7J28F3SMcfYyGC5xWpXsvdm/CX76BazHetJBFvV9DV92b90wAxM0liOXWT
zQmmpMsQgUuRW4X3C33iV9IKkLZV6V1l/H0hx4EvOd7NeWEeP3tQ/aUokREAJ4Cc7Q0VQZjBHUPL
QGVr4flCIgo3Nob9v6CRiDv1VHWe9FG25azBjzrpOcNobf9odemEOjnahk491sD7D8+Gsjxo+2yp
fyrcRI6RU0NJ2fHK6SI4v1bADxDRn/YDU0oaQma6QCjTm23KAwcr+Uj7a3VaDW8IEBFRA+TKveIp
5WeH4glZEydQoZFn9vJxRs1MajrAakfKhvmn/P8PKJJXtcWc8pGIZ1NqX+BOXjhLQhfHC9HP73HJ
UEygUPMc3fMWbe+86YGlWoEJ5fXb0d1J3KLLz2JJHnZ33TzrAkD68ixIhpvC0Kl5A7zhxhi5U+Gs
IYB23XBJSi7GRP4fEm3uHEn3NmKxTbC3qKlXxVnzK5btCRBwCGXC7cElaJrHoBV9DKtaO2cQLvOs
hm5XMRPKBL19HJ8yhXgRTbX5RDXWheKDWezIp+l6zEX+pqAnKG44lZ/iv8WCmVjpFxTaSl1g6lTy
HBrS4O9r8gJ9zKmEGRdxZojMx5x52nvmhjdVzX5fGBJRnx9e+y7O+ACBo1LN/jxLyWZOO+FSt89k
cJnmP9WZ9qDSq2xgt2pUZRFf/TKx2QwKuoUq0WJH+9flXJCzxcVx/xRfGpmeGqDZ4jPbLaysHmkN
+P2UIx2GPv3SWd7oUDSvMMuNHhqeukyeVikGK+IPqS7t6CzOq7/lSYSy1SIffyk5Zej8rGQjK+1x
O6hqMua9OLMvOaojTlG6jUNKZrC/ID6jhdCz6TxKN8b4wp8mfrBqh4q5TTIKQirV40tqfUuo4k0r
WJhkHWkR8miS/z4XFrvsJMyq4yqeCaafGffY4dvwP4OzP87hDrsiC+NcE2YBPkm2GUeTszu1B9x9
RYgYbKKrmAMLDKsdlhxWe5XOXaNtWtLHKNm6U5DxlrV2Ngj7ma0C3nVJbUr8A/FzgRzyiPzv+zOX
/8GK0kYR8YYlK8LMxUprfLCErF4+JwZI3tNsqD/7p4OPvr7SarxvZYsv2l4nrefY+jFJJmU/kIB1
PttreVydWs7clGMxWNbsVaAxfbH3Z92w6wAF0hNiNEx1ThEMlKq0i/qgLhPtOLfL3PS5YqiCF9Au
GAjiy/bg20NEOJoSHWJRcmhMlW5X2+fSKmbAShIk4YSr6k7DKEKVwgnfxgqoVUYh2rUggBFQRLMq
vOrIFiGScoxjbuBzOjnCODDz0HEHh+aj7ES0LE4xSb5et4QSFO28+smq+AsYFoCjQXhy5krKSch/
M9VVjB52ZaKu1NtFiR1h2DxfmEc3/gXsMovlevoWs7fbibilOyRcK3dlCiQxhVxBDtQVzClEv4nL
3EmzLS6w/Wo8ShX7eXuU3V3DOVpEJDJB+iAiy8YJyCZh/eQzOv/bKud4tbfWFwDQlJYOZXoetgXY
5yF94Des4nWaeBpM2Acoc/NSLwzK847oOO/k/VPy7gDZy+IjpWvJ8R2HXEKQCh6pU2G89fbbGpwh
OeZUmYhUD9mh4dRnrpGZGlaJ8bfNZymSusvR7U0+w8+KrJ92vVzlZaWXElyNzrU2EPvlWjjarjBd
Q9+TL7/eBOybrK305dexZYO4CiuPmfxM+NnHTTNHfW/lsnEvEpgdjl0h2mntj8I3bLO55YLQNL4E
AfOAyhsOLTjwrjyni/RHGvSu5Ewu3vH7bTCAgZ5a/dohFCuGsULvkZEG1pVHIvPzr1XEScm0IZtx
JSuRaAae3bmhc7nNsrKXBWYKKOx86pJx3c94rojk4x3Kd/nMdKYI/nkQo2MXMtjNdU4HjkKP5nb2
JM+1yr5DbHKpQQLrleFimC2VT7dTCcODA4dqZSri5LksgCrnExp/JOQY/Vu72uQ/LwfXQj5pITb5
TAZkgDBkEfPIuSzHWRHsn6bRG4FcqeKGjlpXafeWsrK9dBrOt9htrJkFk7VHu91+CY7QUxCdxNMF
J7D5JPmA2qqD7Dg1UHDlWwFaN47dinEBUOlQKK/UHI1VRs4jTXE5EvuR+9M/kY7QlIOEKZ8DjN5b
E5aICHqjrUh8BQKYuBArRKn5b8jQRGh3fuAANdvZ0Sgsp6zRxpvSQhZkUKjdui1K7Pe7R/bMiNT9
ys/KjTI1LOW5EbF9noU+6ximpHvbGgVrRJPM049QdDEi9+/c5lUR4hozDoFRHbpJr/6U14SCYQpk
Sehi/YbWVHbSNSLmEMqKcKrXFVycM85YUD1AEwQnMPLQSWfStqbEZGOGU0w6sDzZAPe6LIZ2YqDb
iPVTn439M6wBzidHT2GroSz4C86SPZclUxait1E6MQYKPVaWTbjG+GjPba1P88vPvZ7RCHe/brX9
hW31igtMcWWvvA1ItpmqeZgqjMbOKmXe0EASllLgzd9X5i8iZPmb0NEAR1H/DW48ywqJjl6pbRdS
GLfDQ+ZtluBeEBaTChmD9KnDXl+sHoumVweuPKKNWPTANqqS1G67pgsXGsVLNS9vcUl4/L5oSPS2
CQj8P43Hl54ffCfsNlwj8yHJVzL5smLjbx9m27LAGd/GR5jmjW+Q85HkJG5kt4lHVSK8xZxzDNCN
Npp0wu7L73JLfOyw9+NYCwhVkZNrRKFiqNcgm7wgYvYZ85IR2gr0yFRDV9iVp9Xc2Ic7JhGF+TlM
kdvwVlqsAuuWO2o9tOEKNZsmNtLgEmVATV7T23DiRhja4Mqsbphbjr1xagH3LWpV+31R+Z13GgHo
aZ6Wv6aXg3PoWRrmV4y3Rh+Ww8PDwP3uLyaptNMo9UNSRZE/+E87IFo+IksOxCpqR/aaDSHYk8Cv
JRu4Gabm00f3K4g8a2jjccBcaIJbEEIfXIFDg8ZBMOrJfPV0gNkidMYWocIWeoq09WplZHisXrdE
kmv6SksoBUG8HM0P5tj2EG2JXjIEQfOefFOzk7zmq+n1bWleG1Bj3suKtVy8USzE26IaSDDl2iSx
/H2TPbYaRa6W6O/3AP4JPUvKAgREPyfJnpexPAbTeMYJ1eh2E6sIEYnKCeG6tgp+ibbll0dx+Fq3
p01r5mdkGkGgrOHmIiVoAJ3ecK9A3By9gCswsu1ywHs2J0wAJ3xM2xNtV6P/W5NUbqXEf03fyb+f
cH26UeVSY3IxX2smCzxw+Marmka+Vmj4vdTEs+eVfpKbLQ4zDUHt5DoqbL0l6VVNq+kz5rBjDyeg
EKhHnHkR7C+jA1KGpRNzj//mawzaPn6tGS6ibA4BLLludYDNIeIv3w8f8jLuq/35PMQacdIqzfgH
e042h3MYj4tg0I50EXzZz8OzcZL6mUZUjbvCXSG5++8o/WgZEHmhkYCak94G15oLfHelxLoe8tku
kWuQrWPSjWgj2u0WEULhCBVc+idA6nQsLCoIL9IpioyyNPa6GVSUlTNYqZdfcvxlRc8deGDYgbvO
L/jXC5mBNbt/xpsnUxRwBfKbWF4lceDsWueHHV+oFtJheC/9jYuE847e5kJ7eRNr+kM6GreHX/bR
/B65wHVsW4F7TJgO9nvs+Nifl+rXlGczfOXHE+k/bwNLyWAdDK3xMH/AaF9Uc6NqQgiHTG7Y0KQi
X9hcnSTh8zC2wx5ii0G53ntOg0c/Y4zNihC3THI4gE9JkE3IXNKAsRhMArqqXVhR00yj1CcZI24l
1C2rhdU6d8CHyYb71QRiCjishsYwvRucvsowqlbP0iTKDOlx3rSx5HI8o756MVNOV0gGUcevY2AK
Lzx5gnhumR7O6AY7tDg2lgB6PLRi5LVznreuS2XMKxXNX2r0sN6dkl5XjMvBcs7SADLzls5nQCxI
iV/V30dkHTv/3WDWoaN2khU16tfCY33tXzxU79PSvDucSP12GKJ9qtAJeC+hFDjBxdSZ0hl/IHDx
oBuYqfXsq85zKID7Tc2i2hi0xLdSql7uai+5L7mnFjfz1j1xjxEBecfcxHflef5uDaqs1OJQWMuM
ROmbNHbFPE0rhX8QdATpqQq6XB3IAeznIlUfCkmWh1BuULm/FpyiZ1VYLxZYqEhzU1vNabntXljf
DDTWXjX+pPtFwkvqVkL88zg63ESwp3loU1oU3isMwD7e3+K7RvA9gkuCGcLQLFMpZr72KG9FLkEA
jzGJ7SzcZeknDvvXXR4EgNAbo/QzSFL906ZDvMLYKRcC+PMtlU02VzsmC70llHwadxD0oe+Hz4/t
sEL09Fr58xOvbl7GDxpzjKdrYTqIGTwovccePL0y49TPwqs9S3m1xDbenASgOD8My9EAwqoAxo9u
dUQC3TnsObv98MkjpX8sQC3cCY7+NorVDU3bDTkvsN2jwAFzrHboB2fBtxOTQe9/XQrqnMkwoWCC
YdPkdX26SwImkzHqUChnuz61O8puBWrT6KElje5GDYv1Jxs4CBgTr+239p71W1E3c0MsOkSqrVa0
a8aTfH4irWLKLX+9F36DDLCwUwB7LZH7iotZX5OIk4Vt3yFWMFJ3c9V9D/eDulq0mds0uFKOdk/2
dPuVm8GVWvG0q91WtbtqRd7wAEa3GeZAqMFq5dS8euWXPIV8CSCrmpFA+Y9zrAg9KjYzZP5+HnYy
RoCyX+VxQdlPc/03olCU6VuCkGH6Dze0JZVZ1xEDCIljkX/XBGP0hPOsh5X7zjNWm1PvfBZSo2fv
iYpLMSQ/2omaS6Lb3jBdMGly0RVe1Gy++M7pLvhAw+CStjTlOq8Lqop0Bisi8JM+AgaGUGfSyORv
z809a5Z8DF35ff3GHO0pMk4t+f0qWbNmITSaGEJQAIWh2NDUTvGQKsYK2Vfj6Zu+Uf7yq5v0m18Y
R/XO5k4hV8YlXjlTHXZFXKDokw9Q6m/BuRHQwFA6bTAR/KPAJcXw7NU+sfDTDjgxD9S3V0IyYwse
emi2s22U+lqjy3ZgqSwXMuIDx+iukBTYvy+bB8bWw479kqOHa/4xPMIIVzkYJ+nglNqyGO6OolzF
k/zpGO5EjRNqaLFG0IuChp9L8fPWRQZ7FWD696anpalSnJo3pBurV9Gz7Aawfu7rT+SmBgDZStsv
dsXm1lGrsAeXpsXFsqiznGoQM6VmYwZ1FX9vnhl4jet6aaSu7WUEaTzUGxfmfdmhvV7C8Vr3krgO
LPPeGYa3T0I66YOtw12vRvlJolrIok9LXqIvpBFNzW2aM1irXoPD5NJjGRs1iGYMazrMqzin4Ywn
OXaMwqWBPizYDmkoMvcFjks5gDy4qdIJ5uKsOxyynVl3ifNCNc/y8LV9/n3kGjTKZKPcZUBqRZ0B
MscjNyY1juTboveh5frv0KswzC+6khEcCf0irPWKJZgkT4SysZ0fguT+JehzVW8voBQsJkE7AsYr
aukmsw01mOtPFudQq1rO9gwK5u2a8OCSBuwsBlNR3mWO1SGEbrizjhAeUux567bkY7Eywc6Sysuy
DgCDW9hPzHOsjjf2ewvoharVTndk09TXqzdhHCA6B9XHsxJntNpj6OUe3kKUCS+gV57gtMPsM7n/
+j1I37oK3QKEaSIx7baTpypADbGAZCjexdQvVseexByrkyl1uGrtzUnIf6k/FxdNm3cBEliaGrHq
sHzrv/tKWwwPQYiQ7s27Keh5ZRL6084V5U3rCl8lmaLMKEizYJ28RaZUOUSD87Rv14+WuABWNbmD
sXTyH5oWmqGyIJgoItJE4FK3ZpGATBgkYiCAHt1h/D7IHxi9lqTQHzpEQLP/54OQEB26jzsjD1hm
Zq98J/3xp6WusLGElStJvsw3K7fTDbJ6/iv0grbK0Cud7bzUVPoLWQ7xUyVcXa1HtLE4F2Tnwmh9
9DmH3d0NYnO6TEP+uq5paHb32aaYAq4q6mPyh2aA7qfE0GgDrTM/iG9uE+CVUMXk+TfWXiCQCokS
XeqN+/XQTfQOZhSAdJ4Cz9org/Ymhy3E4dFvFxp9BNIwMlyjbQ2hJpwRyLyyxThHbcJ7olhVqNNf
boz1OPCVHr6axH0gM1Z9ppq7p9hb4z4FNzpHedFhxY0xTV4Zr6K138sp19pKMyttUraPBnJKDROr
QAlpKPhfO+TvKVIqxaCvytPnwRdx40Rv9XOXKB3cozmLxdvei3iMbV+BG1bhB+OCXtOoeuok3f/a
U4yUnktQc5SKxHpeZreDKFEx9WI8kmkH48KYMqaP4tciBPfV+rIfUO6dpmYmXMM7lUUs7rj1KJCo
lFI3USHLsizCaKjRZ4mmdFu2uhN2iFsm0uNTeSjeM3YiwDWESqx8V6UmYhsRc8gFx5p3bQD2cV5a
IoDGXy9cGwwzwaCHJDB2s/lXxvmTM3uIiG3eBR4I5iD6QOb53ozWCrV0RWnhTSz73eV4dv7abigw
4S++quOe/scfr2hdILi7uGJ/jRUBmiO++akCf/m4r7Gv0dTzRoIAdUpCp9zouZSDB7UoOPc6ojdW
qeVThRLE/FIagdrt7MOZbhCcfEM5SpP4mSEPJkWgGE6tEXZk2TB41U31CH0P8UbqKV4DZVuZ694e
4RB3Yn+0blXuXx2hA6Cbj+BWvypvd4U2B+zWBIsYFsl+LjgrUzuic/4XBphDRNH+bcZgxsOCUVdD
iLNKELCvF1tKqgOtrolkUHfH0S5RiLjYYaLJfd1Naj8/QKshhIMd5ROFRLVptI4i9eMwhR2tgg+1
q3CEuKI5EquaHlw2KTPyrjtBloEUmk2Rn0GPB9/SUAYCQV5ofN/0sjriZ9xUmSLAjsXNZAFfInSt
CaZYeYey71EASpwfz3ihsvnyaB9GhDZAiQDYwH+Pn/6m5HMDqbCGhlGlEV6gQK67ci8JgoywJH7g
qclZ2Zw/8/bxi0DOs4MP5z4BvCwrwkBCtDdL2QbpsHgzqOyKiyaYQ9wnZdAKJ5CSSC5c4wxRONCt
PEe+U3MIwIBhLc/j84PpEokaFHWApJvpFDnO3xuCTbWUEYnUR6bXN1qQjOYD7BW+oDYroP9KOrbB
PdoVL0Az/lxk77tFHcr1tMCzKb5d4tlpIX0tT1xXSI3xmqaq7zmRj8zBkZzwfhd0IfV5HZSUUF6k
0iM/tzAJyobpxKXIxNv9QsO2pTj5TcifVBvZYdU1QDqe4En63sxH8djNx3+pF5XStYWWgUZxZBez
gV2gL/jKs4VT+L3N+nEJXzOCrm1YirRRde339P31n151iychKbxrV8aasyQ0o0TGtN72Xs/AJrmi
ugcMzr9uV8kBr3ROzb2IxAGtfJ/oc34gji3/QIyukWm1OBBIxj3SZn7dSVKrE7GKMH3ZgpxEDkYJ
y2c4KkIRKLHCf07FuU2zIfDEj8fC+PMieJ3AMOXF/NgSMLJ56su9TElWuoS9IBu5DooybJItWA8s
w/5VLveNkegMeOqxB+P14ckib/7m+xGd/N4svaQzCttff0pO9ajzwvdOtLpWyoYZKtQMkZb9Boo9
7H/G6fzHnnmsZlhGE4FZh7TDdFie4MwBT4DhzStkhwO72jonOzgv2EFG0lVFszUxLalHey8n2Ul5
ivLKduokoJfUCrnz5QlhwsbTqX4Dfz96uvbsc+QUko+7sWAAScOo6BWnUJcOAc8eG2mKB5WSnzyo
FwWsy7o0WTgF/biwR8HvLf9KE+S5lOURzWdKwaEM6oSMFQiocRrNtwVXUj4tcqlMigzYmeetBiKK
taFECblFm/yyd3yy77HCBzBet8g9rqnu6TE50mRszuw0aD6UJaqHdSraCbPYC52E88hUMeGDvyi+
21a5NqrZBmhhMPCbTKLp8xSIOK74JIIXnWvI1BqRIXwkT/VoSTLP4GUQgquYijomgveuGJagJLEH
bx01FKHuEmqh9Tmhx68hHt9nyd5d7G5wGXgsGS+zGYKxlgfrbyY51Tu/8XU/kl5fOIbEg+rKu6c3
1/a3l6QM14rncqCD9V/iUvxpC9ZFKAD2nfp/sDdoJUoMPm0woFGy1DMdddzclswCBn7z6nVKzo91
5+WJuvQrWhd6RpxzonbX3lr+iuJ0MB/R2/3Ftz2Y5aGnPKlAl7eUk2i+7DOhNo06JxqZPgM3SVFT
j0BcW2MTWjj+TdBH47ydQyY0eQbr1h9+G77MFEO93c5XVWwblckB87Y8NJT12+qcy8aIMARRXuZn
akipON1ar0EwCszEsnQADm+hI0Va93zUtQ2PM+JEKVPSaNMHRhxqof08ixX719rkjvFNJG59X6Im
kb6h6kPzq0krGeEpKjJGg77VTZFeKTweuPbAVxK5q583nMOFLULsiwl3B9++NgdTF20OhNwI4+ZJ
IFgwMj46SEVCQsGADK3jmbIx2pGVUNCk9G5e/N8Yy/cKzUqGuQ4gVFk58V52qL2O5WfjjuGxZI1W
tHjW34U6OWObHA8THnsMF5cgQjvn/GzP3MAjnaRhjDMVfPg6z6+PS2VYy0ZPrdILRKszwLTezyoz
nzI51FnJZ8mAl4nzwMPelZye3E9owdvvvDqC+58Eou84+qaykPrcAnnDwrldszs/+4jTi29+mVlz
2cy5I9Nbd5O+G1Ne41HAJNGVbXbxP1ZFV1oxJJrLbPSrh7pTUrNGF2PKz5Ruu0GrxGjEk2wkLviZ
xIgVRctZWtnXDKaEbCvdrTla5xdoygWNQF6aK30XUEeHdbhP6FAxhtjdII3RgycJzKgndCXUj4OY
OjPhujt1m/gCadPPcWXCgxwoiUxcSbgS7s0KjvWMLgZ3sQXjynXEE6eWjRvif/NomrG01ejN/VHI
+EFXvoJAe43bF+sqje7uRbwQMrwhiUHH3Sm7r5WwQJHdFdX6VaLFZDP6J4/ppm2zE792v4nC3s2z
i9QfKEPqCJR5bYkKr1z9uTKwo5RHPXFbMzSwxwM19U2vNDMho8gPK5i/JyY5/nFOYy8PzQkF/YFw
gDZlcnEJ/km0K2RMFjA1zGLiZfAdMZ5/UMCbE4u90cTbGjLWg5DixkPzbOHCO72WAi4P2oqKr2wd
V8+aESO1BPLxP2fFdqs4LZlbq2U2gKK/qYdghCP4hQn/lgMMKnBdkx/ply9dQHKjUbFbo/4FDsIa
OmllehCy6Ifx2Fkdx7QQ6WGhQpTKqE6vZJ25cNIJ8rNiWK4DdNUXEN9iwwAbLwIgYsiW4eZcrDYf
MSY1AuC/YfVbrgzc/qkHtTxJ/mGyzHRfRiscpXOywI+a8i07ag4xVyu6h6jsQudOwTYqD0W+EYcf
2FkVkNkR3WYSJ0U4EG1d2YIB1jY88V6udYziSIoIZuRj9JQhW0PRtZXdLF40MAbju7lKCCM4a59P
G5a1V7r/vHtzxQrXbAdOfDHVAj4oEmbkBk7ApjX1L0fuTwJIyRI4UR2A2VJYBX46YHljXFWhQy27
tAxlEaTlpHb0h73HAto7Fl/9g+VgQ+dqei4bJitHlUad56GsyJbmJ2t0vnPvo8yYrur/U5xD7/5F
FqJL4BkuJoc76A/+vgXermoWh/uiBeZxhMM3eNu8eJ03uh6ToOt4d+QwF6w4sitBnOa+EbWHe03z
W9aRRnAZzJENEimANw/TH1slCHFgLNKNMH/MQqYOS3iqcaEP0Sr8ZMq6vRltBYC+qqY9d25q3B3O
nby7pnwHfEk+094gpblRXXR5FKAU/tj0g/GKdc19WG4JVFokp9vWJvkv9a0IbGnSWYkGGkp0kmv6
QwIpIDoxv0Bf8uAlN0PSYRAr08sTSSW0gbCPk5TF2ZO/4wHpej5k/JPbjWNi8V34sNYzbmkKQnd9
hIdzpxPONnHENR44EzTBJ6x1LC0VNV60vW2EJsDTzVCol47QyozYMYW/T2M1o0rZwO9VH+JUNKsF
klKTZ/150W0WWr75NBVv31zYWGb3xafd7FrjNB12NES3dZQ6/JBzp5H/sp31Q+j7fQWFZiKtb1vi
9lp8REPOg3mNVDY8pe0nxQWMzFh6EOf/s9jATRCUpN8jP1o5nHc0VeOCWiNVLNWqrn3nUshsLSW2
s5zrrgECSMPxN8TUjJbeePcDsUSEHmTKIWXt+nhbcE+fG4R8aZoF9wts3bSYrVUNXMxuqzcma2Hn
08/QFXsD7w8+EwYCJ3giNdJ/cOznrkxdjJyflHnpqchyfeQqtKCughdycwwgWqN6M4J2ujd0lEZy
lRc3W7XO3ao00CCihydRsW8zzThvlvJl2srYw5PNAbvA+obAl7TjspY7sYl9k4X7cX3FvpGIEQoq
kY7F5R4+/HPSVHpwZLP1DYon+296oF+ZQCJkTJTkTdJjE/73mC5WGA7WU2+dqgnrOQ01AVze8jtP
/NH1btm+ixEuJZuA5LnaPMwQ24u+10vOA62Sa2tYDI/bzTHXj6RDStMCyczO5/f9+8vahAOpSSoR
6ahAHe+XS1TXDr1SMjoO4zZOXYJEd9x0nQ6pB3lmtmxUDGgpaBrJrNu04uRNnLk+Xi5CxaWiWnKp
A9QWR8C3+I/WTnlnw1YzFyTMYP5dqQdWYn5R+O2uWQ73/0WNoZs6J8BxZ7clmvZlR/dhpCvjnkQs
ebSlYdrg1HsOG0k8F2rk6vAuOxkLKc3pAznrHxdjI5r2AW/fBYGMjR+UO+60yhIKSLLFQyOeCNO8
VHW8zYRAAp52UGiWsjrdS9uUAn5UPS1UA0uiBXmDsbxBbG1B8B3LzQkTrofWtCn6TrW0bHGfvdc5
lxdYYEZtr6gBG5YdIGUzM//cA/BXXsICsgp+fG1Tlo2MSSzH7zLZnsb+X8vXdQxEEj9r1lnOh8Pc
y+0NvqZk4W07h0K38iApuR3sa8fE0L4c4SgyrrDqiKtVNmr9y52cQwLYNDCQLAjGTfUp/SnjoJX3
CeO3WFBQF7tcv5MK7ntbVkJ662Bc010yJFBQGI5t2RySYQ5DkBfnuRPIr2EJVg9JSIUUl1buWavA
KpQ484gtJOyN+Ps8B4XQV76ZJfKWK8KhHGCUjsN5hg0wzROiv8qaEDtBZHniapl1qZ5PrgxXQYZW
VA3+gtkyWI6j++nB79Ndqjygd05+3So1j4jozwX2Y9SHHcKcfhQ71lbXQgw1AVX2sxTZs3k1R3wm
VqsF4hQ/rEBml1Y5+DmSf50tjCiZOVWHp7qqkvIWlfUUjbME3f74Yg1wQgzCyPGhyz5hP4m/yHoC
CYOkygZYuLnWlQXyf72aKUZEbapJ/O1WvT8ncYL3gCVtS+CpIMsHYtoxVvhE1JkfIBNh+xGCGrtB
8TbnrXnlynrKwYoqNdM5mmiFxaCIcQXIPHgEIYD1rIIemz/urLMFYLPUIfTTgj9/gUvsMIcauXZ+
SzGF6rYv8DikRny+SU9VxU6Q/wotTj7gT05Kjy6TCxXiuJgQzt0oTCc14U/XXw2B1GlooBcSsCdw
OJdzjUd9TkkQdiK/LvNcYJDFGc7NmtfUz9QDHCjjpzQ3YfP2yDSZoi4NSNF3h7dJC5RnprTMnhoR
eVVEy1ylFoSa479jsOz6ltJvNXbM836IpKhlTwB7wH3i4C5t0pmL9S/KHAEvbq0+lE85tHuFLaT+
+wjthz7B7gFT1H2M61378Aes+df0mOc1m/LF5Hx+OQ47Kq+VBRcYZspezNr8xO6eQHnK14ECB/Vw
a5mKAFUQdcSz15sxtvK1ULT+rHpIVqfbxh0KFAvJmVKTGtNMnre7xU04FR93YioQ0rlp0BlIqlLa
+A/7P1h0nGVNV7h6Me71xvb8IF8mlr6QWlFS/yXL9ZiCFEU5pdpkq3B99ugHvbpzJvqi3weBcGS+
FAzlTCR6G/W1pstEtDQW18ecOSVXe2iWUd/thx6j/x9HgCqqyeXPwvD/oBtd+0bQto2fBiBR3itw
3Ju9LAK7+vHyX2TacZcCkvC9XZsfzXqwxt2XrcTYd+D+5Mwu7MfI0h6i9z9hXs1IPwVCPS+GLEkz
ssdiBpmKyHgiU8Ea9+tvzWy6hRBNHdqS+K0gUH5fLP2Cb40UUgIKxdW4y+yc5MG5x6lhurQd5ntI
YNmMEErd9HVQmAeh2V7WXp59tnN3jePxrm2R0gd6hfvNm9GguTOFdqkeZLylhrIBAU70eQ3IaAXc
28bvE3YJWG4FvEkfkHWedBq5x56m6J05YDZ8YeOJrvRZGEHBmdt4TMQoFqOIwHbadNArn6/Bbrtp
9BOyQnHnEt9e7Fis0S+oM03a9xPvR4SlIZwvjjtO12P6UITPkoAdk1QM8+JDjYrxQQKOMbglXG1M
yxVNjHLhkQCcVWfZcA7M+w7k9V6Eg17sSpWkEDKHvQyXCPTGBD5zmbbwVJkcks9u4uDvc8Tzh6dX
3D/mar1QekRoFw637g/00aZ3MLjRYE4pCFU/ieBuWT12Xq16CDcYtzY3FI2jazULAjVgJ205EaeA
I5aQcfsYkhC6zFYWiRFPLuk7yuZSezceW17s15hTYJgXtxv7me2/+qOIGjWuCPJovZ7u1a0BkEqR
p9jXa6Mp5vwzs+8c0D11mMjdAVcF0nadG30UAlKrRc5IBOFxbFnJcdwEMkvfX0HDSp0XZmIXkc9g
EdROJVYUG7FFo/BBSVzFhOsIji6i4birUR/vljc3DpVUWP39XnWQpiM+q2MoqZzxZXYo6cy9pUS3
GMCol3BFOxv8nvIh+WJrSCDuDrlURizGHOdkVS/A6ts7XKU9ApdMiiBu7V3xhxN/OUbD1VmzYD0k
b2hWKijVoNG9CjHHEysOwkfnhWltlo3AZUa92u0rD6CPukavgFPf6MGh9u/ChSko60S9mA5OV9cm
jPJnLgTV7f8FIpVyslWw3exISTXVoodOtayaCO9y7OlIp1qkAJymTjFXhCxOvS5D1kwYcz3Et65U
g/ZD6xjahE6L7qPLx1xQVlWOngroda/iBFBpeaM7tSj5Zw1WBlgmDB5h0bK5JSOyk7M+f7urQFUx
vuEn2dLpFBjseZJj798y7YFuefzdYH54bhwcx3kI5mBVGDXHZ6b9/KbBDD3lU33zA4tmSzxN+0a1
aGvJafNNaqBw9Fb26z5EgR6wfFDfrIectjIbe9rVvLlHeusEn+q7MxIRP2Mq0mz3xPS9ywWPWKFr
uXLkcO5zzy/11RIYR4R8TKvNUp7MOjcpoZEhqCX3gtt5TqBZUouvGiQu66/u7dA+kzReKloddn1z
p7QfvOTd7Pu8V54BQromLXEkLlHI/odH3noR3cAuGej7ngR17Nyk2U1VgucRrdRwRAkj9tBg6uPy
+6nO5JfNzfof/Rg1eP2nO0y8TqHhoeVDn3VvOQfxbJayC00vKArRkjb6Wmnjikl9fW4NYimvhqzX
LdsbJ0jFB7+figQB2DQtOrFpjW8BIOqgZtjCxH2nHX+nMILoyvZWGBCTPLTyU7OpvoK0oMF7rkq1
K3Hr2iH05fl2q6Fpv9YsgLjOqe7YrTX0Wla2ku3rDiIoFbCPo/J1peMzlORgUmhRF/5k78GQjfVK
sBxkVUh2gt2nun/goH517vqyz0PQRnhwW/lZjUum4NxIEQ6oQQJTC8ImfKHzrreZvG/v2HcGkEIJ
NX0il563fv+LeoCeRscL2m/sZ68AXDFhe6n1fD4ANYPNqm+MlIf9PIfQAgs18wbg+x7gXOp+f0yC
HrGIJX4hJi+ZiE57tZL6PWFXeOu6RXmI/9qDTU6YkkUjJTFcP5+imj2RDCzkM55M/Nx+P/B9fCUP
X9w+svDhh5So0GMOoBYrNW6lWSHd16UjDPPKrUpnoBsX+AiSuQ4ZR0fD50s5wByivm6UIBLaCAht
Q8ygK9/wav7YG13UMiQNdblFRprQRy2FgBFDcS4mGPaIgHT6okJLqqgjEgycz4D6/KDcHnQbCZXk
aq/AofxdIA6L98LFnDKnyZsawI1QINadpWeOBNGKaAoxqC5+iFDL2eEmNUJiEJ/Hj79N1tUE9fNE
M7FzU2a8LXHPiK6cRcySYBxYUUTVm7NWy6iH6gMRwXMfmk2Tw1sClAZlS/hx5gEn4ez1V75YAcIv
DBm2vVC8lp8NLmOfWDOIL8BlRlH7v+f3WI8Kb5SBE4vZ4fs68P+PJ+hiWj0z4SigI8NFMwpvkh+K
BObyCvMKcXzusnyzdTgp+8kXsIcJQnLyrTevsPllRsS4hBMVR9mCGniq7VCGXCA7TM6D2JnBJYNv
Fxq/LCA+DzdoC/SWfzatBMI2SsUKwI7bDeSk9RhHW/CLz6FHSdTnne8NwkPPVyOf2Y2cA8y85ycM
qDNJxfDayohCaCfcpEVnqPybaqDQlCv5El6/IN2BFMeNa2sH9TsLKsxsmlaKw2sDA9yFlSMGQQJY
2hVbd/NlKOJIBDDucC5xMyK6htYheb3N7+5OqcYk5jouoL/bfDZA+vvyAdA2ITJdIKxwenrzobdn
hPiBLx74aRGld8H6up4zg3icWUScIARodrHzu+gwu8g3402PsXqgoVz8Bh2qKjIIMSS74DcOTJed
44bw/eg82e3Xsh/M+eRiX04sA6hsE8Nij7wDuFjQ6D+8F67EVGSCHeULYlQApdQU4whmhiYKu7Mb
JX+sNywl9XpIQ0V06wZH2LF9E7dcfslaCQapqFCH7jiTDPAe9LHmaJyfPcvI5MnbaP3TKnz20rxU
43hi/jhnXwBIwR4YYNfMOIqhZvga822SDMUzajkPwCl0ytdL7QJoHb2YA/lF70176ARPlLoCASzM
ZUUJhBSYQ9s7GvnJamBEILrWBVCv45u8V9V4k8PIse5KYZx5OTC1NTGL0m1kzTgqd5WBGsz4ofAf
pd+B3GikhiLrli/ndNM/fElq90Jyp88XNgUDILIN6SpuXL6pZEHKaJRPz27kicUPFvgFI6c3sd3s
RnCW7n3iqJnJV+4486yevLOMomBdj7+15zP+SkIUGzaCeh5Z73zhns3YTPLhqmhgVbZWfnr983Kc
9iC3r83vSwYJwcNNHv3FAXCZvZxLnmmCi8myZdQxSJB6ZjXU9vYEzRH+hUDeupKCYcE4/vR4g4r9
okupv8vsF5EVwbRkVJpSmouESX8LiHyOjezF6HEfaSiE5EHjcDMdwPiZCh23AcOmlMOnMXouvCxa
3wCBHA7wJzBXS4zfuqXUYo9xMm69ZvpM+5AEM8iZChD44HbSS1LmE2NlcxPFowipWgs4ISTBTU2P
Sf2Wt0yuAABwn82VG2lZYaSVvySErvZr9VCL/Yk/E4paERQKuKOETd9eaBExi7zWG6IIRJZAhGRw
zofWIyhzXwQQGIIoTGEHw/AMYS5JDXBjV3CULmNuUBZ7p4Qniv/tNwXUsfrla1IgwlD7zAKDAcXP
nc4T/y9wOGT+OhEqiw81c2WYXdGpP6URQ+qH3hKHwg48xd8hhxwhpSLAfyeqjDyY6E2Gm75oSA0M
7m5gf6CikUqJUJNDvWXewk2lgF5PJC+BrVvY07l7VQixRbUnwULyt5rGop8EO0bVZtk3iupJ254n
Fe49yVEzYrvgs14mdq+5CqgFcbRSxjWbVFj69qTWkxJuN0gMGgpEet0YEFcudGT7BkxF6XEOhpAQ
DM9ryHyYXkkSI123m4O4JfU3bMJW1PPr3Erv0+nagNnzOvn6srkUXCRcEAo/6FmPP0uAc8ILAGXU
MFUM6xh/9C9zAX+DmkvC43VuiwlIDZUu+IXm6HU9Ps1mxJeiFEmBVPv/e2N0tR6y0U2hkIUuwe+w
mdhYQEPgHV9mDT6Goq/MtG+uMpLPkmJKdveFrYLmuwvb2gKXWx6HGacgqb8h534GD5iqfxkaI9An
QIKyX3/z9V+drRhrHeY76PK+MyUF42WSwoah6M+3yJFzUxWg8tm1NFu8XAc1ImbG6x1llFcLLG3Q
JCenPndOv8DjwExCeF3rsKJBbIIXLHg1bp+gNkryL/xx3D7v9B4n7myGJyU067eNwJHDTyA8ZP9S
+hHZamJFor0OAvSx5ZL0dAJl5TBeo4lk9CwsJSrzMPymD2ekJ2G4kK0fP716B4YvYAXX4rIyQDg7
R8yyIEQoWIPsOX+zYtiaukuVS/CpU9EZH3K6lTlZDdpsvkraxHlD2EctWcXHUWVoia8PQDM6v5CZ
KTmYAQzqBCXSCrwRzT1hSSCJsfifp+z+JppzcEvuqEz4ccraax9X5DeCbIS58AH6+hfXAqhlUGNu
bxrn29KtyuQ5nJK55K399dey30A1XN9QGITAIfjJ5GegY80rLKaGM3bz0/0F6PKGyD/LYTFJD3cA
49s9RKU5qDeuD59RHbjvthIPxileb4heaeSO+BhpJ20ZestYLendw8Xg20Cf7hXcSFvxwcqXikbd
cS+GI+lZ/kqDYp0rLAHRN3yQmhOtqyuASntM4Y7KOUtFbdAeoXw/al6QmGD1AmUEDEYTxQAVTqXK
WvuTxPGWwPwYBiTexPbPWE6StuakAS0M4ZQi8DCSs90nsahMHCfmbNytac7fGLFqFHmKRY2pcVJl
nA9x7Yf6523+BIt0+FMiGpXUfCtmf48elBHj0vBmWsYGfl3rxtjK0YsM1b37Fka3ZftyR/RDiIw0
GsQx0LqrXgfdYjisXLKyAGRU3ZVq13u57hTkOmaZ2Ouog/KznIqooRErEJvppWQvaVbvwlW9i2qI
VaBO3wJxOS9hxSUZ0c6rH2eMH5RJoFKRFRKjrdgmn6C015hXUX5NL/5FbXep/87LKA+Pf3f7AIg+
2NOc5+x3dWm8V/801jOcwjth1uF1tBo1j7jjBgKyfLuN1+ppV039Qd7EnTP1dZ5h+z0mAe+cJ1HI
rS4yTH94lsH5o0b9TwyZMCY0qvp4Cf6Ps0w40hqMHcXFrMQ5JeST9Hn+H5cg8CxuBwpo3do3YW/6
b4Z8DDcNBAs6EVFUqJ5UXvNgAUxeqVaC3AwCY2jw2mwKJFtrLHSnAGr/SskRIPUvPCJhOWpD6twM
gicBtIkD+u8h0s2PxZ4EJsSNYRDuqf4Qaqxfb1+ROsaCyI2ux1nYOW07JxXkJuj1v+YbDMLULGGz
V9+BqBYooFwuDaUeHDKdfcdNwMqTJepF+rUuSwqY0UBTglUmGnwHgQEcwgy6x+CyMfLZADpQPHi/
p1sMF1zDpVIO2PIfzpdhEGCSBsEblwOJZuytDlY74UU7hlscOetGjPIhkb01yUceHxv8bmLm4QAs
Vn4eDEolmJvBN+OTa7cSDbF7wLKqBIAgrp3w3vqySFImNsJFAfikwqT6yRQ/VuBS61lVOracppl1
yppO9FAg/P/v2ORNvoH6m9odxhGYAoU5/5htAptXK6VjcBJhlNdvATsKBonVzzrKOEwhZ6v16Mj+
KUK2dMwwWOPESF3AOzZP+B0niv3GYwFAGAy+dQi90FnHXoruGiTpKTvbq//iTLLGbn15u4xowC7k
CdqA+qLOFgXMSq0ZgO62Pzxrz89nWbbube3nXQQT/k1EXM/z6Sy83qlsw8/t5IF9xYYDH7BpjHRA
xLaHleo8GSDCbR3qaaKf7UE5sLSZNbI+oc4f7br03OmeCvgRoUTLsvq8mRuQ4Ygn8COhNr+ZS0oq
d1x4netRDespOMBWStGG9dBm263CLSKc/O+CWjDznSZnS+7+NCaIKLgcNe4E+GDCjXS1ymaAyHOt
IcBK+kQkHFAq9wj9n4Aw9mwxIvEmugo2QCG9XQQ6C8k9oI73zELCqVkhyxCLNk2j8DVYG5rwvxcZ
gJEz4y7ppX4z1lEeAmi826+Nw1w5a/02a5KUW5eeuEOp3gqMYEugzcw7HgwVzI9mAJH3NfiTscVN
uAFey0IL9iyr5J9bTuxrEkulHhFGrut0G4hKmoaap3jJwaZoDR3rzZ96kppNjwGiuLaVCKY3dyB0
ARfzpwyf2PYjpJeAiWrMQ53LABbJYiCXhRtubYyo5vKuPRAmmTiSUPYmP30Pv0XqHN+j2Nf8YyFK
ute4G2nCL30bv0bPXbU0f8Ba5xttHM1wpP42llTkPekD+YO0q+zJ6nxXiT5fisYcTpvD2qCTn8v+
dMioyY2P1tbkoL9PCCytlGQ17DNqxbdSlXzAP1aKpW4zE+36suH6nHp/V1RV7o+//isRtwT27Y6T
28Y0BGKa48JYiLdnDNRmOESmOdzMEAu3JUqKFGwES2CTdbq2a2upc8IDruAwqLGYANFEiRt71lhM
nJ0ShZYbCGKZ85WK3NYIfTpFuJ8oKTrzd3xdwd5cpuNX1hYRfkxLFshf8uds4Xo/fNSJGudas0o7
NX6z190aArDOYpQDQ04TGep8SsNA6/zlZ44cjL+riZpA9BewC8yWW0Mi+2qsMf39wAeXSnREsB+H
JyQg7es2lOqUkCL0fSR6b4GsPN91fYmXRjPLK5dUW3vL8eY3Yu29LiHlbUVJmvEfUIXTDV2DLOlY
c7p2pj6p2J4cGcK7NqmiERaYEkPbJZpK6/RaYXHQj72vxU8XlSXrSd4ragB6XbKMN8udFC+waFPc
XAS4OWJVX11cH3EemmqmbCu0YEWM4t/ZW6nn1m1Bisjrtk1RDrhTCU0LDNjohgNiWYfVGFHGCI5k
IuZXzIbIkBXaLwt1u1H1gpXBonHUGxBTjUOnXZnb02WYsitknhCjBb6oVuwKnaQFNaCMW1Ced5bY
irJQ/tva+U78QUdsFPYxSmku3+DK/KTF1nBEsENGYzc8T7OO0DlpiaYCMF8A938eGqnT/BRU8E3i
BASBMS2OR/GcpqtVeYak78dr9FIWq7HwvNYYEJv5BBvo3y1zZvpD+r+UWlTuW649Tn4lFEaclWLv
rjiVA+C7utlqTfABqwExlAZ8n1BUd9CnzPi5+MoGCtMZeMmWwH40LKtDC+91Q1kzWQ5UabECi2ov
mHURLF27t6pecKOUMYz/0Jh/bQz5jAveqivpw5sk1cK8xMjyor09W19rcbVx9xPm9h3o+KFmuz2H
UlEqgouAjsUuhHHMLMeST1dHzFGAC4eZcmeR4oRYyDEzl0INSm30SHwh+L1Wz/013TSdP0zoGflQ
4oC5IbOzlBMtflJoIf/F/b3OsEt37H5P003DZHNa79HaMgRhFUcf0yjh2QlFdj7ioOoYEu4qq+Hh
ozvlAVbqlgDf7rwN6lhP8VWuYDUDL599xfXqmABo7j47IBObLewTyYqh3ZJ9QCMGCaVji5lwqyf9
F+KBdPkZA1+9qQlGR8MhHIIW8j3Lg173GhwTtzyWDgPC+Z4Id7cWVScMY2x+oEZdjXh80TqA0Fxr
IYvOBwTNbY1O1siKHS7H8jWbDH6EPS5wEg6uAy/gcObYLVMH1lCKj1TPwrLl4QKzG2KgZ/cY8G+n
6ttByjXgD9HVwFbnR/O8NzUSRhtbmnteQbFcHp0dwPWY915Urfv//JNkZN3DSzOCSBH8aWP8aAWi
lUAiv5irLNiq+qppUE5ftFF9PxU3Uqr9EeWQBaVKWsBFq/iGRmW4y132cT8gjWCPWN36a6RrGxb2
tI6sLeFyV0pvggnUHCaK3re55d3xt6MeOTc9aTLsS3QbnnSasO63DdXpstxvpZaf/DOYdswAUUkg
yjYTcgMJzJGDocRYVSX56dw1Dtw9jNL21g2zoRRfXXQUgklSwbTC1bzxwmcVVSRL2kz/BCNJ7Xkd
53/7lbkj1pHkZfpPOL0PVxiPROimFE8Wxza3p7ZeY+e5zbMDvQAsX44fos44XjiiuoMmiEG6Hh7u
YAZYbfdqDm40Mv6ul4mBbXCNuUXPAwg2D6LbrBUVNRGY0N6YqMlNWUD7/uYSgqj1PwNVmb/9TpDk
D+Ydi6pgFeyAmx7lww0aUAEz8IYadKSWcCvrzS9kChOgI/ee4HEHC5T9jcssM8ueU3xAgbfUlwsI
wE+BwsCjRQ9Ha3BhZHORfFKgkVQ/8L61VYcFsnp8OpYC6HL4gpnwNLIMbm3T3MSON1TGWN7UyzA+
c27nP8LTY7qfOjhLTvmZ9uFDvgpKgWWgtEHsmrbMa3GBUPO7aGJ1XXCNO7UVKrAnBYONfexGrSQy
wTacQ6NrnLgCsm5L+teuei6KOSYgrQ4D2P3ALg9FZFBa16a0fs2MeKZSgzDH2QK/WjRU+IhOFWpO
Lk+z5GhhX0Li4M57PlmUuKHI/zFyKNDVRLus+bjRyd0K2g21PjFKQqDtXlDrnC9l/InO3xsm2eiR
LGtIbp2g7dGawUF+w56UAdxEZRqtmFkZfKWOePNlq9JI2SyPNlXRZNpjiLliInwUurFssobjKC4C
PaRXGkmLpviOMIYSraTMpkMVM44plXcJBQG5OyIaKMArG7XLVolt+jRtZ7kzi+9Mx1dW2jwComtK
kL7DQKXKvjI2H1iBQR0v/KjFT4efLrKDwEL6LPgYmcVh9Y8hbXOWsbLWpUOmiUtbzQShes94wEeN
KjY4xhqUhX5irrUrOfMpKEisXTvJyWUuzM3EOKfnoY2ImQoZCyvxcvaETkFnFufFxun7y7/Z9hAq
y4csKR/QnoI6JhsrxvLZI7Q4IXgi4ELIBL5vQPFG2P2+ICtrOc1I/tRQn7n/Fq+wvsUR+qzuRDdH
m3BnPW/W/V5RVj4FzC5P0IswzsB6/NDcAB8v4Au3PHZwAVNgBgNgT0R+pEPGhivYspdK7ib8pRp8
Jvy+BxuGCMR0z/DErJr5o/bOVd39tXS/XPfi+o/yh/JJvZ3cvzoVb2x2JYbvDyRFhjkzIjpQJayq
eGMpFVaxFAgJFcpSbQHgE/ff+hqcoXDV83POoOQaw8249IGDkAHIpnuGflbLlddGNET6MfH7uSoL
hTzpo0Nrswzx4RvVBipXGluE14cC3K2dJ+W1pB6f67UrUQ8lDnXZiJklh8hF/xkH6s+CyiKwOP0e
XgYamVyLYsQuwtupUCAF3Ftt3WjB45oYyTBoxzufj4l4lu+Fx/d95w2fcPBDYY8pSh/41jS/BUUS
1rSH6+2fke+dlIRhv3IArNXKfs86UnSHGIIr82PbqxPmZY0VCwzVod447byfy7w5/gXfYnoMR6pX
F84o/ZySZCz7ocbxOBglDheh2Dr/2cM9Uv/YnAqEBVfLrOQoZC8/fkbDFuDZq3NS/UIu6tEEaSm7
PKk9RypYPnObAUvRAmUcJ+3F9WdpmQJO+7noAiyBEIV0X5YaIRKN40aS9jf5OpTf4uFKopd6oMQh
kZiBHX42oC6TV1kA7DQvG5QPzhsz0Qxy1mxQu12j+ndcIEaeYYSpvSP7+mIceS+X9D7x3RkY6O+z
uT05E5YrOrWJvtspBfjvobwZoi0wF71l2UT0XQfPWXcxcCT60RUcm00dO/u4GAARuqaTa6ODdHJx
YUvqpBW/GKlva9vv0Xjgv+ShopD1mRzqx+rjMIjupKYKNVti5uTm4p+ifnMEvqCJTp+4KQ3heL2K
u+okKQmfkRi48lkFQNcCrmMUbprHNzijU9bv2oCNv9pLmfPJXdipsnZyS0n4iGqe1UKhUwlbaB7K
GGTLgJK4ws95ONe/qpySGb2iRNbkLr/3Wx2+s9SsRucdXNM8Bd51NlAsGvcu7BnrrHXsJG30YztU
ZvfZGXUMd2YxZ2xTQDEYQ3Q1m2m1Fo8RQnWz2xa7iCpvcVbfpGWVVxzU8zrtdOovtYyzoLgT0m+e
Uuzog5JWVGAAxl0FRp97pqc+W7HlTRt/1ml/Cidd5pWbNxz2JibMaV20HnIaIJKy6+rgLmzltwQH
iY/HnvOv5MwPN/y8eSWBe+dk3ZYEzewNM+roQ0bvcXmJkHLhXGIibf4sT0oFUkras3g382hx8AqG
jWacq6zp8x+aJFZEd+LIfMDluhB1aNCgXrMRe+BZevIcozAfzpf9lRfVTLSA3mLA00REE83kVUzn
MX5rQpmFLai8kWWh0QGvcPHuloGrNLewYoYa1AaQKqlxrXe3WkP3BueQUB3zXylMiuBsEfB9AKIV
KwlnDSHbwwCKjNP9OfCjWS+BDO6QRV57PfthdG0pVSrNIbpxhUzK+bT6tmLy6icSEiPgHQV6wjyW
vhBNYovx0KdAXkfxSDuaYj+YG+9NuzWo1EePI5LUw/kXXn/qxA0BjASammvIR8XWfl+MiVijXQvP
5+pxfA85tGx4jD8cTpMmNbUQzHBGqiNgtmoWa6zobJa9n72jHDIieowm8/5a3yTkgO3f9ocecwjZ
nYxVEqWQJZ804TuQMiHvElnS5DLkv3UH+INRohplcEkUPMviJysF8osvqo7TDkmw/2XRpa+qEVqu
sZqZXWek+FzcKmLtTVftr51Rrlo3jJpmFeBDBwCZbUcmx19QwTEtqgEtOQSVqzx887/FR5ecgrbP
OSewq7UFp85rHko7FD9q5WbvWjVTmsAYS78M7AQNAJkbcvZZmG9WgP0Qa8mwA+cOxCaHUCdCVsrA
z79qDLrPpRBHBwNIPC2rdt2BM8QyLlbaptbRuX+EaE6WtWqq54vJXNatLXdSdLfenei0uo5UDV1J
PCYRlnO4lftbiU1C6iIKj6wiVm0mA91eOl0A8BJGcT2wIZsPmsxvLhsAGdmrVyX24ImdjpSgNLsK
lIlmXSECQ5mk9ELtPYrk1r9slDFKEmQxVTGQw7ee0OjbnLVfHg2wiQDuKzibd2CP4WfL14wlFpwc
3bOfdyoOzjcPXOdXqhA0mwQBU7KwdDOrcVpBIcZtIDKhextJvhlIikGePw9HcIYR18/GTV3UMJfr
A9mkGEB1jcucd7M4+G+MazU61G+hSE3LpiBj4uIuaqtW3t4JUpQ+7bS/ZVij582UfS5DADPzmcx4
9iczfHYsvatzE18dVgrDbfHyjApYpWwA1m7P3q4OvRit3pM4NjNKjKdM1vIJxDnvv3JqHeA0kp+2
4/2974Nstnk4Uy5GA3i5KOlMnA76s/m2qg7lK4GfijU8Dkrfy2WYhGpfbsYOWMVrnaauQ8WSq72g
16bgFt015hZtGEtWi2+RXuf0FR+GeL3HWTP5MBA6hC7JfYcRgdnDy3ZB3mD0GFTh1n8cK9+rjVhW
4rR31rjftPYdfclzMgjAbRoqBJ8Ak3PX6AIscFWbGqe+1iB5ln0DnzvbihtvNOjyt/o6A7B8nlL+
yxMHU/KYvq6cVnrZIKX8RbH877MmMAPRwe+BKw1OLAiqYGLzXhtwyNQ41f+YR70/rJlhznmgQlT+
bTBZ/Vpzv7PloiM9i523Fj8rv2SxGulyWV1sNZCoEIWl2ckuEz8bj9nxRMIASD1nCN/13AMP1nMo
Ybtsn7r3scLEFucfo1ytAjVnhc0CLZxxdfmCqNAAbiCmQiMrFxwhSlRg9PUL/Bow8M9jXWxXK020
5NlKozdL+6tBklUEt7uVBdbdh78xAEQ/Og7XGDcj9fEEbaWJroraY1ejWrwx9msoivvHG1FeZ8wc
H0hm21X6tiUrjNkQv7jt4wTMA4PNbAP70+W/w52GzTE3vcO+XWAIm8TrJlgK9aVvNf53w7G5cLD1
ATZZ3D9J30+k0ee6WUwCiNkY9gQc1+TmF1QrnpzjsvVowoUvhVd8KsaZ/4Hs6CFRyEwqiSeiDszn
EtDm5fYs1qrScfFPYcJjBOmRvYfyyt3oaJV3cw2BzI+3MVfZetvKGZr1AcSHk5CE2zKeTklHDKAJ
IMQ+2XIlxLMRnVK9WtHH1vqfYKzB0MAKkY8N/bh/PLzhHrVBdkipMRd/ZD0FmVuMTcHczArHmgt4
y/8nhsLexkE4m5K01K1dKb9/ZKd3SP9LdzHdetZGSayc5mA4VIt+eB6wo20PpOyAgfgJi5DwBiZM
LxWeD/okdM+pi4HWsG0AMMZ5qTfKFqL/dLY1w9hLR/b6iEyLnC/0uikSiny22WoZ1j3ztMKkDQ0g
Z+kpmDNwhhFGit5MkFzMlE+QCDSKhVt5AJhE9FTBcvoLq2k6Z+RlkuequVfiGdt6XKQ6zcVeIgE2
I02XDYyoRYzUaZga66EfGuJyL6B5t3oB5p8eG0KcMDaJaT9MeMRV0Uu1jCBJEl3DCnhXkr1X6cGG
ovgZ7L0OPWR+AchL3sVQhbzZRzdLT/hRryoA0VlTAJ4dFt6Lm3fnyAwYxff4gMgwhl5ATgW0QTEt
gHalI8dfmc97Gq/HcNvhUZXPG9FAJVxjvg0fuEAkWFuvxVGN1U726P/Tcj357XK+pES91CN9UpM+
RvxojSROgjHlUDgf56miK6/xdmum9MrvagsaLr5AgagpTvCDYvrJ5+J7HwVAIvWKYBCia80y2VuI
n4z9h//iSef82uXlpbgoXgh4PQDVLXStUNetFTdGR0xrnIM3ORe18MH49j7+xHJMOgAbT6WJWDVa
BIxqPCT/s/uAYhWcZQwz+wcO9rf6Cxj9QnWCxls2lbWacxnHQ8Imop4ArENkZ4oFKfhFo30lqKIc
4h1AsxHkQ3zNUXd3vLNCA0bspJgHA19EH/ZOZHgWWAhFM5243qPRhRyPOk+4I7Mj9eNVSXjnC3OH
9CHLipiMHu8YP2AmYKLbfytsxjNleuO9rxHGGhBw9EjSQr3L+AjShIb2z0XLMMM+ro/6kCqh2v7y
IQdQbYPOX8dZ+nMo1NqFC1HWO3rINK/qjrbxJnjXcVx1yB0T5BZJYT2TAyRrIsW5fva/1a6N0QiK
t6EGfnBVi/JZNi5HdA/svyrdNr1WpHxI0Nvbh1gHCp/dvAfG15Q441ErYSZJO4gMoGnBoaGc0gCK
2JRGVkTSb6X3iiAaXomEpK4NZxY8azkXxQLao4Yr7NS3kH9s4HOPcu/Mt/hRSrdMroeREj26BROO
LkhkwQrvQ6Tj+7NxeWsbtLs0m5oywOFhgV4tvR5tAgzxeA6jrbimkdjDSN3TiIR08Z8ORyWtZanb
+cVqdYcylaWN4o/N8tCAq/tEFIxu8viC6yDq6+Km3TGZGM6jnLGi1kHLqd6qLRhTc/u4Gr0L3a2e
t1CQ1NcyaKBoVfsKkfRwy8dhPI1RTdsTIGB7bIHd/sRJayZ9+zUWyEssfZLRBhJn0lUvecMWyJd+
/D67DYoIVhm99Ax3ifx1xObv8U6Yt3kl4IRAqL5Pga9Av9OsJX9t0U0UnYGd0ouQExW92p3IphD8
BYlBK7yn8pKtIQr1Fsov07ob53MmN49O2V2kn+V/WxPhsX2/1opc1l+axL1Ccgl9QAzTgLiRegvL
BmZzcjdqdY8H/+wacz4E/Wbyq9FbOyF1VYDXwjZaLR9l1g6KZrDCeYQSmUHl25pDMWO3+GeJO3wU
ln/+Cw1Tn0iLf8gPzrtGR99Qq4s2EwY7BQgadPDHgN9MVQzvX5jJ0T9dney9XUAa3MWqoVDFqASh
ADDU1ZsKzEIxiGFXAQPXaq1yhtzA+tpNLDi/oiH3T6EoMsCIRHRn/BTHq6nX03IsxhLPphKexXJZ
o69U7Unk0OEUt5/JdT8undOU49cg9I9XGePsmDqPJP60sl7r1GtgmFwJrNp4Ev1+7rcSUOmn7ZXL
jLTpfeKm2clCn9iz3Yox8O69vJLktlyXh6ioJGleRxXM4FUEkuiQ71RsZwyniROr+1FU9NWllG5l
4O2oJfSWuf/oulUJOBUMCYOdNRmPKkUNLOYzkVBss3rCmIrJzMmsS1iA53x4oQ1dn5Cw3IBOac7s
JzAmNkQXeKW/9D0OuvB+vMKBPrC9eJJsB6Ud8VzjmiB2DcsVB/ICx5481j1nOUgWhFmci78EFlcC
Ins7r4Y4yHLSGrHh353Nf1BrDYraWjyhDaoXaSwst3URehfAL1APpgRBOAU78xQDG2c5W45279vz
L3zEQNBYSDiJW+sQSJ3HMp15bZ2odorWIOAtVYIJr8iHT1uQHgXdw3ThLIGKNs3ZliKwFeuOSepo
EQhzZHvM+lGyvxo6h+6qovOhp6VKSCOlEmHHr0lN1vvxEwHAKz9PYsG+7vCeaOcFCVx1z8ZN2dVP
iafr9kfLwhPHpEYw/bZjMUJaEW6Bz8wo3902PVUmeafsqQbB4ixGkBx9B3NiVX3LMG4aO5JG7UdP
/xF96THyZA3bUXHRT27DOz5mKaS3OFrTg7GSxbyxuc04viDzs3AqYXBP0hZEypP7TNpmP5aCt+3p
cgCIzni4s3RXEMjR7Ui+TB2W7Dmq50sHDS9zngkbLx/qxoXWFxXv2+7fCO7eNJZKLDCFHaIk10O3
27nha7yoLoKIHTUr7+5mkEF2M6HWblnfWfQNeXblidpBlwCDMfGfYWupSPSQ+me/B7df5eYAtDMZ
cghJhsDoIpFJ18zh+YJs4tGXlWTe9+Hm2cFvakUVSk/dCAgv1JaUtu2gG2lPrHN2o2ErbWzER4Mc
Ddi8I8/9Scg1OeQRrsPAlCi9a67L7Y8VvjRgHTy8rgo3/YoEtaZURLF38TAejTExBejTjTOy8lDA
BCblQtMlgaGMU4at9Yo+WGAquCQNaIQyZwDPTPAnG9VhkfQ45QxNXa2T0JrS5vi8WBTBKvr12Inm
0biwHpCd3ccJDJlikuXzlo3ukJggOwB61S5X9sTt4NqvyxyBDIDCdFagiXKVHmvgbsxMGjZBO/n8
PddkkKwD/ucHsDFFxEloi5n5FZ+kM8F+gKpFsBNVM5W/5OqMeAIVhcBTYLcnb6Ox8td5Jbf7F+tX
cIX/GXo2bxlQbDj157Rj3bdn+ZmWCGQIjLz0Scx/2insdduWnXYTe40vgZX9BaMDghCM+At17OPe
n/ScCfsEDuavVLqmXxgH27ZYtJnAaWwt68jhalyKqSjWuuhEst2SKx7yWvAeSodSM/LWqEyUTFuP
UO3I8aySC62G6BYehaiPvpUfBDyt5QriCkIQm/q0nzni8sIFIsU/0E6b6tqvY9Qtznm4ExybV3yy
HEAwhoG+ZN3sefFgEAFQd2EwQuShXCYh2JfVrgbdQi1I93avX02lzNBIMfA/8AFvV1blDF92Y19d
ZSgHdKadNYEom5JoTHDBL5jvLWWQNvmYk6L1TLVEVdrxUWZQm4rQbKhlqpaPTFpSM2pskiDZXaBK
q7J2VLUtlLehHIP12sQjdr2AfzDSzeRhekSP/hPfJkdHcnfADD1QWjxbJ2S4xvMS0OhjCkTqOA31
DeYSxYiuIOka9YMlpZAxpnBzqv46h+WMU9jgEqeMMOdGaWba3do8GnyiXUVQ5Gp84K2Er2XR2ug4
+yHxNEkjgEF2/D6BOOEna3/fM5fSVD1O52L2iBKP3AeOAZupAkwrnA3VkS896XijM9p7HVasL8HO
JFcRrckIlhO6RymL1oumd6VDzmADzzsyS9fo7QHeFF8VIRj6Q5+gJB9GTPY5N90Oyd/yl2aUNX9r
3vZhtZXrtNwnuNt87T+ezlbNt4sM46Wl3JOyN+eiafY/+3PXSwkBUR3yCngfbKP+2pa4jWfXTcuz
owZBaZxkzW3mu4fLWreJ07blqzicNcbf/1KLKm0d7N6tv9+4Z+YVrot6TcF/m90QulFCgq5igySI
vuSdfyjNCyDkmTSdhmmvtJoNcXzfaHBO/woHNveqb7P0LwHOgnAkKsSXBCLce21OCUx8TaLEpn24
2MG2nUP+ry7EBe9KmC9VrfaicKT+KIvaNNuEC8rN2WY9AM4tuYXuDndj817K0Ej2SHHTURMUXzFA
SiL89tNSOXOuJwqyhO5BBv1qh2U8Zcwbpb5hqJqO0U40yTdsAr/r54d0mm+IwkysgDX/AxMzU7H3
BxkEbnUDajmUf1Ccd4oq6h7vfW0KNbZ5o0WzwMra4mQGj4lSnYtD7BmOa/1p1GlnFEGi+wkE1vrq
32bUMQVADOwCs+ppPFCaiBjRWykv0S/LS4DrQN3WbBRxmgGH4sOcaxlg4/90fO+PuqCPmXNhSNjn
dJFSmLNRNwvro+lNYzVLIQnGwKQfszKuHq1ULbmyyGFku7idSL5RWvPjyMV28KyiGVkTd1SzcpHr
E0WNsKgbr6gzGvDZ/G+9P6WdX66Mks4b9W9Z2XFW96bJOSoup4UV9cj2hAo0l1t7OfZybDmis0fG
XyVrwam37tlBH6wMoI5Yn2XlXaZaeqICKbFRqMDji/LX1/hzpdjRvXaDUqkAKsxynKMdbQvv3QEd
d6Ftun1G244vy0i2mgmCUji/8U64pWA93fGNvZK3+lFh8ghZn+urnPI+fBH5euXHIU3toe78cZ+p
m1MxLli6BJj2y4Tc/As0fWqSoF+i31B/dBYt1i+C7ULtBrMAIVOZx5d9WEg4+c4CSMCZ2AdURCPr
yi+HJjlBb7Jy1CgsVf40L/H/w1SHNTTdvMZoMdA607xVvkjmmqSQF9Yadz5CYz8S7b9+5yVO+P02
CiOZe54t+YkZ5xhqJ2mMRGIceMU2sdU71sd/ocvDW38KXa+k8TFbxMX2/RcmWOdV6geANcTiAMoz
Jl7tmXoJYlzRxLeaS+9qKmgtHnTel6HtiRoTMj5isz3ckjhPKntVOlXsAB65RdaRUnlhimyuGeLp
5F7JBkz083Xqk8COnbd0pEv+pxIXunmvrjnCLyzkTT2fxWXHfAYMHAsflRPzlYTeY7YegQESv1r3
cgLqxczlMMvIDX5IbZagPYWNKsytohf0UyHsiuvSAA7RoVC8+KZg86Si7mP12e8Sw47aNMa6OwhE
tntgntxpMRHvWEPHUusrxw3mIYYSCmsSWgJoM0gJRCPQaYqZe1izj6zy8HYiQ6spUX8acsuRw0v8
n6pFp6Gan+HgM8i//dhtc4hogaUrVvvc+II4Sz6Jo9Y042uBYHW3e29N5q/KImoT6Vsiepu35iDM
pzUt1pn7/wAf3MupqqPV0ypn1ww0VpzjGKe33DEJmukvGkCiPbxoFRfgVWyo6hvMUq4BI/iiHBJZ
vG1Bcwnc0+EUqTLoYssuEGOtIxN1H9yLdJnEoK7d3MlZNUzx1U0E3ohiStWyUEC1heMGPxE6iCA9
D/24W2ihMnloOeZZwXDNxhS8MKvnd1i0t7iGhWcX6EbW3bXs1sMrOuEVtwWbcVN3mQrDbmnV2ZUh
Ia5Y5J5eCJCkggydbEckNyeMp9KXFtA+1dMoufPz/+ZdVXpsakKaY6z5U3PGSoQ3jmukH5p6r/WQ
XCHld4btvpBlfG7Zbnd8lhNaMngphpVBZNjxojT3bOrVh0zpC1NIE5IvHtkIqCLIoEZNcBQTfymf
Bp1qDbD5VY4swm6rPDaVnz5bANItzzyKSzGuPyDf9PKDdxJARp7VKi07nNY+3aSVIqasjloC9CnQ
1AZsydYM8vAtMNmEvvluSU2AuecJ7UpiZTBZdZ68zhpJCq47c1aMhXmB3l8bcfeRgV3AAxzdEIxX
gsGCbAKoaYDnkXxH6KNyXj+u7IZEIX+VPSaQH/Qvd2YWW8uDIuZGgfHDFC8DlUi76Qe0wuYJ587E
QakA0P3LJHixkXxS6p9NXBd+ozo+pKV2bWJNp89ylT1GN7nNRrChGZBcIGBr6Cy/1PmiWAKfm4rc
Z/iTQL0kaI5hvin8If4tgCg89jZ5whkAXgoqR9seMnR76YYiFV9iFVZolG7MstIG1DcpkOci4SYF
hSNSl/9amsvk3aQigbSYinNqBqSnzkzWdrl71/Np2F+JIwIFHrBFs8v38jgLr+fUlzKusPBdSNSJ
LxOB5+UAcgpPOhHUIzTqhWrkqHV5JNHG9Lj7GBKzL6Owd5PTlopbkJD/AX2QyljyuIzvjz9ul9Hz
YMNHU9KILdzbQD2KHht02pZyYnZeOxTvHlp0WoCYYSJOtYKoUch2e5AUIPek0jUhKEn+OzUnX5UJ
KONF/Bs3gCHH2aZm9sms3NA7285t+/mEGlZ63TiurVQGmDqgW6msV59mGAwSWkHY6185jaoHV0hf
c1//7PkY7r0wnFFDWEJyQkKjnOLXfswrCtNPcx3jaoU9JONmEWo0RI1pUWIlOg4OFCNLeXNNTPLf
mM3TycsTtWBQabSDOaIKr/ZJQqeUM/lkh3RDG+9CQpRcIqLsJdP5M2e8l0OukJJT5xrkMtnfYv67
whOrbammXDNgBCHiHia260T7MYmik1TaObYP91+/hWGbtD5ZGgkU2uEH2PrdgSTKHJ1rHE5fveXf
0x9azUedG7GTAwR8/m8PwpV4DYw7hCAOuFEnME664xWl2NnRuQ6waIrcZaNY58048+O3BkU62N4y
eyuECjjVTgMqxObuGWL9G9QVmLNyrXYioqcA9KA4L2yc5CuKnfPElRr68DO/4z46Tq6hWK6bu3Jl
W4qmFCWdxzF+sUVRbELaQVKeOdhC4UdTPzHIjeTjfkth+6lYBI3jsXitHrCOIPU4nOR8bNWAHyi9
F2GC2+f8I084+V7RCHF54NjfGXXO1S2aqEysYTE4zEEi+B/LH1BUmn80L/effufOUMKhLFghiVe3
/qfy7u6RIXkGeakyV4T4BtZySxT9UPcAAPRPRUwoGrJbeN0vpTibShmM58o8zdJEKOMBTm1UXD3S
p4q5enE5QGbWpmwDnOXzbayJpq/4I1yamk6rE18ObwskENP5HGDWW268zEHpedrH8lZnbrAGJuSX
nzNx1EHTWI9StJSkBTV/+4CfRIyvA3LrXORoutUxkargv0xSC2liMZEfkZYauYgpK6mIGcfPz00n
nzn+jg3kEKb30Dz6mkC9jxBAa1IQX311Vde2AqxRkuDyilEhUt6S1XDi01YVqaIp1ir55ATS+a4S
cwm2Rf5vG1Ad5uSNH3xV1RtvXQ/3o6bYOLN0CrMEU4ox9qigFgbuJIgQC7UY+yNivSIr36DuxScx
FuDhqGQcF5GRv9WMkBhCXB7euOCDIGXNzNMaD2go3q3U9d+YBBsV31GN4IXOHh4Ph5ashK4RxpmY
k2K4KPRC2F4RLAvgdyZxMuZ9LkJhFmo5fNZfAbYVcC1CzDLI9jyvjFVOFvHDmFHLnnUvuLy9ODII
8TaG7G7UgmuuqW553/oHc4H/87ylyvFgu1GILLY5BtWKANaMVQQbmAtYa+hdySujTzwQxTrf0ola
ZVLU+uz3kde9GD9QMX0chFFNyMzmdGqyZ7JFATtg3DrTwEzJ0FSKVQ1amJUyDNcN1qFl9cZDVM37
KUcHnwHOImtRqVZFh59EVduEG6Yiaema4sp7Up1OmnNGxtye/bABOH5Cb7xO3L9ggiC9jt2Pf16U
/wvKSO6pQJ+mgsxR9IHu3+1rFyNytBvh9uoqpR2JFLiGcKp1gL9W/vxaomUEdFK1/Tlpu+g594fk
S/YZfhH6sUGD0g/jungGBzWeYSQ/buig1jJnzUeSJtXaruN97GyP4LX1H+wXEPaQGEUBiLJd00xl
waWzZpA4in+dXlxo7kySECYKuNrpUSlgSouLSwm4fDEbe8FQed/bD5Ctxt/kXRu6GAmq5LTSgD55
L05TBMSXK3ADpfmN9yBD8ytxQI0gPGp+Usg9iF5rKtJuV9pLn/OmDe9wPfJEodmeUugPFq2qT28g
PYGXpySocMipOG7CW3MimGXqf+7o+ZZ2p4zs8bc2WX0cibynBJ0ZVt/StGwg33z0QsK0Y4Z33YDN
clsJGs1Q791GF4kFwZgCDdXCHcxvRW08TXk16f6StKjBkBtsf1HQRTCDi3Ty1ZqNB/1SZwQbWGB/
vcIn7RU6JP+5uMvMni439QY+lcG0RSKKmk1UjLQ3Q/dA3E+CFluHff/YI0He8ROALcMWM9ravl5n
mg/aTsMSLFS/Of+aDK6Cupt5+ZhQYp2rMMz/eOEGgrROlKjQfeeUljcTrp4IBbkycLWKXa9xqap3
NZ1UrCQBagitNDu1Re+BCYAKQMgnmc1hCoOYpk2LKQwSVYp8QQwjTxtSTLxwsaNh7g32GzVHL3z8
gfI50iRS1h+vIMyJaV8RLBgN+S3LaFogg601+JVfHScd2Rp6magLdpyHoAEIR9MhRHMivaJArarI
LqhF+2oeqkRe0XANfwXSvfJYm8d2QD2/tb84elep0TDgwYUn/vOSM3DPhPGoPPJbxOcijVUSO6cd
UiqDhZHjTueuJ2XM2i6tcwRYo2F0QpAHQeYIEa4vEpLmh5vRRb8hg9SkOqjmGEmdyZOtN1XG3MJP
MCV1UuN3QbsYoumoov04ho+FxY/sIlj7Uho34DC/xuIf9MNcQ0L9D4f/Ots4OLI2WVMChMymQkxu
VfgQz9f5G9GUvbqDaMLGuENfei3N6a7yd0I2o5OBt2Uz2eL6p0Su9Gxjps33KHkITZ2qfsDvRLBx
hNMr6MvIzBv6SJGFKkSmsRE4AOZWnK5+XcchCFt0FFxlUT6cl1eGRIxZX2CcanL+GQn96pO5xAqI
RKw93+NKwdwhA+85sgVOeFcUPxxzG1jxEJPcPZ9T28W1MDHrNC/BCv3mjmiQyhKBOjvcBol5/DCw
Hyw79jLHYl8qOCiAAqbITlecCTWvctBS3dABZB5sqKuTJ5AITE0b9gT8lHdPjWYyx6MqJvuE9Wuv
6vAgwlK3pqY3CigbWP/N0t5skD2a9PygUpx7vkAuh08oCwG0YtACNhWL9jayNSIKQ55K8hGqZxMY
UZTrEGCGWBj9VqWq8p921MWTTO6afeKHPmjTHm63x2JcrpzML6q0ZDhl5QrFuI2O1YfKwJ5NEG0d
umLxIQGNZ7mRxAJls78zZm0zpzb+WWj72mMbt0F3j/3K0+HyxVAECiPKqNx5v4/OGjM8PSxWFGPv
5lMNTDKD+PfgMMuv2dmPgQspQ4Bh4Ac5xGUHVn/MzpN7hv5C93uFE48YJFWWORqMaEZwAIkC0SUQ
jr65iqKD6VMfMfpGT60Z2kCaWOAjDnRmCM84KcowNeKcFL2ygH6VV1VXW9SfhZfvcKol3g1K3ghv
L3pHrnms0ojcd6QJynHQhtrggLp/U+Vo8gZ2saODakpgDD4JwnwTKOxesc/kvmsXTlK9v8R0N0fx
SQ4kaAb6F75l/xN7Rb6MCoPenwBVJYCgZS7ZgDEJbA2yGUTvxx+/UunKLE6mfF27YRx4S1yvgNqa
JC8Pdg8ylJ9CZTzLXbUE1g5wZZNZn0XJdZHZPmEnjFlpJIJoTLtMF72WfGxyZ8p6l1TokfQ6THG5
dU1FAx4i6FDv84HIdFfaoDHf6U5HruGWjljm4/2pe07ZTijfKZhfU5J1a2hPQRQEgV20XjsAQiGD
26ySqkQ4VhPK2nK7rPu1Ai9QHoMfy3F/oi64v5wcO3SEUsX75gNju24Wa1OHcqGOxVTLfuBX27W/
MDFLZO6trFJQx9LD2xjDi361a+Vpqxlryo/TNVgICDIHu05wEOtY9ROQ34w5lbBQQ22DkvQTfI/c
9qkr60pnADx268/Up5ga4UZs0rLtvkMzGpqWobvo+GvVRTDDLZaHQBjRBGfi38kU/NK7wAbBwWBp
gLTXl286OTM3wxpG0p8ssv9HZ+kgFLEDW5JdJDQNumgOh/cLo97pvoL1+zQOzMbfiiI+rC2w6tqD
8pp5W6vh/nM5ZNVTABvI//1u8IbEAu2jB+zluXplD990z9wzzSuBOau6zTTUi2s6LcNlTlGtowAz
8ztMUvVKRk2TG8QiWHT+5wMOUDpD0V4dlr8BdpzfydxXo18V66LAosizPdPsCqLHls8c6Tm57+E9
gcxyDFjTLknnY+8QsvdWno1hah4DFEhSuvQGHcx6Wypo0nnTVwK0XGigf0E+qpqq8ClfUKa6qMDv
gMElRTRjh8rvWSSJTiyhYZB8OqRcMwWwpYkGcfVb7q9ZTmw3BTXJX8BHyIlDkdUYT8UndisWv9Cf
Vw7k1+E0PPyft7Or3tPQXcou2Fj3GVe1ttOxiydvU1fsfteXUJTiPamaOx3WhoK7aTpyM/9D9VlH
7UjEuoe32old3aKmAKm1UyumXQaZ7Sgs6w9msmi05m02mgDsYASidZ2gYXYEo62htx9/+ZqyYSg+
6Ct7t+0cZqsA9HSE+KvWpdN92R4NJfO0w0Y/azC4zCrCrjTYBdkjiWnDfapyBKJMzocdtWNVBW59
MCKUMeruufzFjmii5tUcTpGODrdVKO9xhtIZyrGPDB6+s8dJjeFhVJSNmvRRaeqElwEmXJ3F6ZQI
7aZSZrzB0kNnScthTsCT7lZ53QO5s54FtXCB4e4rXrjRWMvAkZtTwkQhXenXV3vOi+bXgGzDho4v
0o/RBYShVDgHnvgvt1oWMBOIRRXk1ofCCoZ+JVAYqPSP7vzfocHwGYuBs8o4qJTHpown/VQDcmTL
KKZljCk5MmXlknwA/bUAoIzh+6FQpA6vE/gud0wWYR66nPbaTsRtjYUOuPLAhnXT2SyVHI22t8Au
upaP9Mwn9q2jxEhr7AQsP1/wP3RIrWW9vn7F5r4afRiQtFWoRx9ZwL4OzWyzVwWwPtINpR4lIZg3
RC0JUf5UnUwo5tTfVDsuQqvc6NAZVKZ8Ipz60x/jW6vlg76/70TaTHGgjTvy/lc9vQiUG7UjWgmF
wyXvUlA+id6Fbt9eKGxaVhqk8UkJvPa/mFbsRHffB4U8Lu2LmHhmmyqbOVDamduON1KQTJmCp4Ku
7VYbfmotV+doHE+w511aOK9qfi47kCPdCZ2wob0tmfCFeg7jRXH3nMB517KmEaXCqf4DeqAKJhm5
Kp2FDusvelNtawKWkpu7twnX6EVwNveFzDQu2+zhDigMCDUdpYdYW3b/0Rfs8Z28Ut4M6vnKYB+K
AcegHqfMsXK7sB4F2045Z2gAmsqCOC1rMdDGfFYjb+3BSbUI1uglpnwPzAfe6B0PpkOMi1UxAkUD
CHhFMZ4/u2lS+rl0fAnSFhzfuMQN9kw9jF44WaEB/OgW2XLKBdooP0W9eIKxo1AdcnBe4O1b4uTI
ZYpCDRD6vYdmVbvUD4UdUqn9AmXG/lOZvBdAqoGxYFBFhYrD+GKGkJZTNC+HZkh8yvMM5WnDb+V0
4P5BuG27s9odVevns15JLDTqwFSlVybu/r9o0rPlcLIe6A+ghMbTwezhO2/xSYc8rherNN9vqaOS
sfPTfhywi9Ef1YJr3qcVyv9ccqwECtzad3hhNtDSzwu4y9O3UGJn/VXE1sYs33kSd9moii/NtyaT
ev+Jc1JCQS0Ka8TIy6IfeF+Se93ThZJ/tJOYGpJcXZPtj4eyhqb2x0k+zBKa62KkYjVyjkgmmk77
OrT+zRsTnsWq2K5Xdjc3RJ+sHUL5HWC95/BfT5geUuWWLx6jxBpNuMw5rLZYcClWz8a7dXTK1+Bi
Gec2MZIXIRqKhL474DQsXleW1uXEHbQHCCjSO1ve4LUVnCY5C6AOFPNsq5VoxA+RMYFUihmjPg3D
Ax9guAuRFcHUy1RqUPai5/a0MRFJRzjSS5CFVl0hJ1HYhuTFWfsl1H8mCXrfDmEu7Yiz6p9lq0NG
L77t35dQDcmSWdjHtbCGswweM+mb9aNg23KQg9V+mN91W8k9JfLAqCt5nN8WGjgPHrCw0cnS8oHR
mmp5d7WPiu8j2mnQj1+6AKwMtb3lDD1QL1DbVgC3Im4o0zQeUmMtHEf+NsYDQ6TIsP+3sZHTryqC
Suq92NrxhDuuzFSP3zucsFvOLP5K2UD7ZEoE1kbhZbikwt3KrmyE4hlo2CZYfx2FpPNf2kfmulzc
hePkKfYLhIOSm6F1OU0OKVFwaCqxSuYGkojGrXPa70M+DeJ9VTdZd1Ylt+R6deKUFUzpChAuLXNy
QWV05P/doWGcROD8lAGrXcoMYrU22HKE4e+hOW/H6BgRP6mBIp9UCVIYxUTRPG3+tdiJVI6e3d9C
t0LFXZNfxCyImpfJS4XfvC2yPSvR5Uzu+sWhKaKFgfeKLAjbFtvvA+KrLYuPZwVxtd3yS4wLA5Cs
H5M1GQg+Uto2kIXlvwwQvowh7VCNiXFr73UfhMTSVF/Yplix96s5kdX7CoWQY+WSNtgjLP+1nu0e
Sf8ca5PVgkZETWECyzo/Jav3QHL+EaHGoaEQjoZgmNGW//lllF8WkA4TzNWZyxSRL/0dLTj6H6pn
P+2/DYyCSUit+NtFxa2YbxM2ChwIJsT1c0BLAZfbvdF+bgYjs5z/0/U7J5UCpIilN52N5mgT27dk
GQaZcgeT6jE99VGB8fHNLkzcuvbj2z64BcTUyW3cHJVSNiGr6C/CwD8ol/hExqqlDZjShFTFYFNb
EePZZhSPhwI+oMCq2JlDthvwrJvpOq2Gr4Whjt7wEAmFVZFXnDKVZlj89z0iPqqAMu5pFDkUEs33
Qz2zQrILVuKjM7ZbISKP7nrqO3HrvXhe7PkH1lO8UBbBTaGtVzJ4p8O27Y267oaUcdRQrWOfmhS9
63bxwu9buSqMq5P/Q4xp7L8TUGd8Y7ryFGrRWVyg6xwYF6hLG+Ke+V6gG5+FDyWclQkFyV5t2r60
9Q8av0CJ/hVS/sCtQWpAs/6B9s7hrf37kAnjj6PBrNg5cCwRrjX6tUH7gWuIyzttsPAdhNbCkNkZ
XtU2YpucrcGWjCSqgggu6qZI/KyUD0g5kKc3KwlDACeX+3BgfYYTEhT3+KsK5nQFEercWlNVEz88
ZB5rzZ2anEDH9sxdHldOW0FoqXtG4dO4tFZ7TKcgh/hCBs1yXROw5o3Rw3c/Tqscbwx+qBhP+qcG
IQTLCTH3o2e1NvEs2Mw9pxpk1cOVeo5KzXVGuz8BdLP0Ph0S1Ed6lJkYjgkvoN7L+2i1KatS6FHw
rVQCiTuC9otTQtE0R18xJxr+ftKbuzJBBwlMqhSwSDN38UO8vMmCjM/Um6urKdaNhz/+VD2hLkCJ
ACEs+0cpvk/lJe0H4F15uZmb7cPV6sveD1Re4zun+2Lhpg3tLgsoaZCjLvy2sbW/YCm/w3JDiEKK
TByARjymzlE1B8ygF1HAw0T/Ae6I015GeEhIVGxQ/Fj93bElm2wV28iHVzV1MLHCJBEJdbGZxg2S
bCVoigVex5Xee9kCFILhbyOVbY4LnXUtMXuLdgote+jfoGz+806xJPD0ENp2hr38rc+L/P6zGDWR
bAgQ/omh9jGABythxYoojB2YlMnp8x6S25DGMet2HGN7kvTCv8oeM6hviGbpivhNla2uEhOgiODw
ThtXHVGs10HRfwTc51/AK7MwKh3dDxRWuKrY4RzT7ADumbZS7xy+XxphTmETDA4+FisDi0Ub/0wY
Izeo0hi2CIXUMslyvlP6qnMeG5JhQ7O4LSwKEKjk+IFEg6k328/6z/q+PjH/MQBBha2GERg/wScn
z0gxUyCqV3el2zvJhfjpBBGHrV+KnahtZ0RNn1g90Ar5ngFumgSOvOIjku++NbgC0bPScORmmtn0
uMqGwbPgGHXzDpecIY2ULw69M38TRpcrAUEDHIsPgiYVZGfTu8s3Oz+zka5ple7Iji4VGrS+98dl
nHEH2mgSU69DGO4KPxfEwUNMjJuCRh/8M/qcLw4TUTVj8etOGDZSsVkZDGjKmYMWs+ZgElHPskxt
VUg5QUnw8f/2f1qjZ85mGy+c1aFXGBtFWgmd441b+0ahEgx5G7X+4zutzxZOfhlACJHJYscx18bM
JROpQ65nZ1k4UfVlmf9loM1gr3qu1typd88vfL+1hWcYy6rdW21Vx65ZHWYqQstG8JvHX8wb982E
MYTGFEAu8BAhZgo7m6nFiDEKBenrsS/zwm+gqlyyOHV+9J7yGWwJLihtkjx4xFxcXdSYD4nh229B
HgbQ2EoO/0HehrPcxfhSY+WkXZCbbC0g+bBQdy6OK632+My2Swc+lzst89P9rRYXG30kZJKzlQKC
s9rMbetUQTQxdo1msf9r/GckGxn4a2WP27vpXQc44yH2A+3Mviztx7To1b23mgWhCVDma3SEaBVr
mrMYp1CtPJVunMOKvyNX/K1Qxmk1Qx0EGpnVWZ4GtdshjWBWZJXjRGMqvymyXgpViC8F+MjtFUTT
47VcqL+VIVGYa67zaFSbNmAkBWf9T/EDENJggeqmVBERVYX9s7q6bbc4bAmUN6X6PrEs8cIcyXET
tvigqwvsdS/MvmhaBAf3npTyxpvfwbfIxFSDKO/30N7EdmzoQakPlPC/aaTEOPJSrFk1oVkOigIV
ICIBcsBhwngOfGq80c54wpWGZZDgZcQn8/cgcY3KhpMk5NxFVanpjmhVoXRhRxvAvDKhGjXK89Jd
3b4YjO9+HhJOs6EIcqgpkNt8tEc4hZCQ4LT+IAhNkGIUP4SMdWUnYBYf30RZiVP9r8JpzPjq2UzH
YEbHrky12giw/LH48ifL77HNyWVWsjOwoS4y7h3dRTwlOGcatojryCHTw9/69fLxTZE+1kw+Mzk4
TIkUn+YPmTthivthTaztBkg1X35ypt1KumbDf/T1XbfsJCF8LVbWDyRkhj/q31CzCdmAW/m7E+bR
Ivxmxm/SEmLwy66BQem2K8woB/TkL2GhlA34e8IlYreLEJ9Yv4tLawUBZq/5a1Y90+oHrNLKkVXj
sa1muENW/lddSt2JsW2JCxifY0DFRrvUeXB6Vvu94OTAi7GYtsE1wLabxxzrnifALv+09N+YNLOL
q0Z/X77dwHrHKNnFFDVtrgDezKQmrh51XjzYDm/G3c1lA5P51U9UK8yRtlpN0CitB4RWRmqozfVL
LRln2NW3+ni6Y/wiPRO5AqCdOE0RBCFYXuYyp/1YRu9Xs06T63flBay6L3z43qH9fwr/Kzl16j/2
jWNufznAKARWS9WCd0iIpRchJbDes+e72tOCB/DJXSvxe44DZMZPWpnmJAO6V8AT0l+8Kd/MDY/6
JymeS3Jwd6f9ks5qNKcXoZiZEY7Rl8C9IHTXXaVmh4L/7cWGbpVGnzSrwe35yH0HYD330LAbQ7H/
x/fdHmSVr0oAquCVDiBS/+56tSoo7WgteATgBxmd/Jet1X68yu9jZUDhJOeeCNfn8oy1RVby2toP
kU7kGLdMNfNhq8AGNZZ1sS8JjFJB3DQuKs57ld6QWQeHCAKx/GGe7U7dHSXqV+jnYJsdRQRP/9pE
8c2mYX90Sd6/sLE9bnsQ8/rfLK1QFGOqZU8lrOj0632csa54XripFhXDMp+1iuhm3fP1VuOmKhCu
1ZVx8Jjy/0ZHykFg4zw1tt+XFj51iMUJ5lrZScv8kAqEThcKm0VaP1sKmYrb8q1RH52bt/NQdxuq
fx2pAysvxf0P4fckOBqYkMCGbEtb/Qqr0PGvCrXlRyu2IQjn9ZvoZGmJ+nXHlrMtf/nj8bc+LOiM
TzNknKnXm+sTRaedpsRhN3WyuUX22YMiaU70CfA93XTVE/6S9JLso975klax+PDNZ2Uv6hIsUrBb
nV5g/TY159l1reftbXoRGD0XZYjjCjTcZCLG2nX2PLclv+/DSdFOGWK2mkgpXIg8hbBGRMoVk2NC
P4xtPx3clmumb+9HeFZzjALArVgNXA3PyhcrP2ua0YEnbRbTn0JpjkEk5DBk5ZJ+e50ibKZxadye
Byt0jENeuMq79TKE+q/uXApd931tPqyByWtVSoC0f2u/BwRm1n560u79kTCApVR71Z5FP5tbai0O
1Bg3DaFHByi5McoFHHBGpVrgxGj1bORJtP9qyTL4twvpojSv40PJST+MP/ojjP34LZT6KO/3NN99
/yTP5mRuPdWg+Xt8Ilfjbv/b41nu0JiBdnrVZy0u4Ykt5NPI3Kei5g43gaReS//BmZduTfZ8vzuq
2l0YZEv2jnbmLVKrdXHAs1mxMcigLtDIHAy48gbh5bxg6dLrzsATDzxxYUS19Ka96O2CPTOrtDQz
32LJ6NQDUCgp7l2IlSv71TfERPnSyDwOEtgzL3Y2vxk/Dlo8CZ9xeQwqGYipvHkDc9OvdGDXwlYT
/mCuoNAe2A+DI9oT0el9nTXR7ncRM7yLJKqAEZojZlk5mb/4ypfTiL8ken1iOGpK982MvN7td7Yf
Cn4NJX6yIALstBqGSd5QAn2b68ZtZwtBOgV+Jp1wwSBKBwSSMOC3fawjNA2Z8DzmXweWHGvYvfqM
dvfmhgaCZxak595g/cHCZT63KfjmPQCnE9RKSsNPr1S9ymCnhHMwEucFMb3VWUO3m8OfK7ykM1cK
/g1yEsAD6jp7luwSyHcvLcycSdrCCevBl7hcMdaMQy+YhEUSdl2eKoBhdapCsxFTt1O99lQ2D0jP
JaU95TwUiS8Xt0hN4ZLMaeBw/FxZYwvf7Ol2BW7+cfVjUvnlZy/8jgEkooy8PLy/75fD30NGg6eF
ZMY8yP5kxb61W09ktghOV2TtbBZpLRta9JftKncOpM7k5vr+Wc+Ny74+DR+/YsG5WZNBuBmIShrk
ELgwoDAQ+anCKh4bKv19ngotoTxSxMIjyPdzYsXk7COjO+Z8DdE8VBQ3/jekXyoGrdD1SWJ0/XyQ
PHLeye1dJG3t9iHMFlXYxAl4SsoUxznCBnniYHTenhZFkbwNzCISdfGQ0krmjscGogsaEEr0KUsv
0+FAoQr1+pDKIRfg7ccMKHnq9k5N/Jiw1whOypSp+l5b8rxtlAT3vaeA3Yz67y+SuwaW0lOPloG7
OX/URQ7L6O2q07bBzHWZ/Sd5s2TejbQRxnMunQVvMAtDFGR2QOyMLkXbfcqo47fuQjnVmJSNTwBj
P9G9NsoR3ZLzfggz/1E9+IEHqsxy/6S03sFPU4aK54WSSzhZEoh0c3nNQQv60h33hJufe9on6SUA
WOJO9499O2S5ojYFnLcHJWD5eZUqu54E0pX8TWCibnYgsOdgZZLcXMHCfIt/BopWeNiAwbZNzTkq
r73WGd+ike3PzC9j59VONlklwkQawsxxd6jeo3gKF8Pc1/bnWS9dhtKKCU6ihGoVMtTFSeAqPfQD
AR3ZviDLmpLZB1xZAJgEpjLYhZukp+pCIGQAzke4HD3ip+G4lgtZtFLmiCyhrjzaKv+OEMvzQpgR
KRtFieDRKbkLR/gSONbjUVJbUP5pbulUjBuQ78yGm7ytMFbiB/nFyGUHsonEyvsBXrIGMnzAjGkY
I8QgL0rYs9kVViWN9f/l11h158I0isT8pk+mB3ureg6L+qr6yyKoLDKJVNz32+a0yLG3mFjbdS96
zMJIEqouqpPIQVmyZNI06N5tkhaU9ncTcw8CdCGVmWH3dA4ZCuJMezK3E5C5yqfhDnsU025fJgP5
Vna/DYRisislQ5ejhOeg4rQ7oRgNhdSG+ohhcfJRHVSAob22QrM4rJ67Oort63HZBPKYGoSkyeqj
VO2HLP/bVxbwCPWA7hg3DlFGZgsgmLVLrL7eZngvFBZv67Fp8PCc5p19reybzQno6exipLWY728w
5skJ/0DRCwkwOYzG1mmfEP1ZgdvnQKlmEcAykNPZqPY5mU4sddaMPYdOiCcMb90hl4mABgITaX78
GJuus5K0qZqYRoA6C6fe7U9tKjp3mDv+vM+z/+Vg+/X+irFdgn2TuTjcnKOYcl95Fo5ZAq9XRbQ/
hiUEy4+vyaB3qj/S81BlncAPn5aSWSKEvmoMODFHxnhPBVnuOIZtElGZgNCzARYIoC0M5z8oqDmI
McU9rC5sggyJYfTwv56LNRDwRv/1MGrTj1qggOn/JHZHyeJqP1AQ+6riINaiqnvAak9lZ2KnYikU
x8XwduEYlf+l+E6mYD8q7zJ0Vcd10iTr9BCHV5pzVz6OF9UFcdccDqCDfP+5q2LRQlL8iKrAK/jt
PWS9pcQcqHny02E+iYK65b/Cso0oIdzutNfM+ulswQtMah9IEhkDIa5A2OsL2iukjq6Z78pgmNrb
EpuaPVzjBLF+ohfCbiKfLQQVoYzFnoSeJpnfsF06BfeCoEJ11yET1hGDG0q/X0eAqYfUyHSodgv1
FtrPg0L8QpYl233JwBRQkrrzq3jdp07B4dLfIyCJLHp/BMkNPKxvPsTUWU40pZgQQg2iBaJF4F6k
W2JUdUBQ6McihhBTjHSzGmtsIFo6zpY80NNp0i3BeMLK+5eN7lUlIuuUJd40XDikH9maD1KHa5oo
bFGfxvd0BNaV2bpX9vAu+1wvlaiy330qOo1M193WJEHijCsGJeF5gz8L5HjZUet4g8Hef0ttqeF2
0Zz1etCN7VPPZFjSMTImdBZptZFzTKRDrRWaYckseBk8LqZoJkUl8oMxSNuf1FxeuDY/Hi6IJRZP
WzV5+4+apq+CPaqX0DkfSYHBx6UbyYWMk+TennH0coBG79g8LG1hmG+zT2l7gTlGht/yc3pewWwa
GpcObTec/fQOnPyrLZIr/EzUWUHkjBnJ0eXvfKUC2MQ3HzzcUypbPCuQAlL+5SPbPJk7+TPVbGiy
/J2y+RtIO/HYdTh3x+S2d38+BLdKF9lwqPsIoV/Tw1A0c6tqYofgQlnSwKLXCUWXIw6gjg5WkiyX
qdNKj36GEXIqvtd7uB5kXKWNQYCkDRliIQ/TbaJEaXZbO54dvObXLqgldnlYDveXW+re2AWD+GjS
4NGAI2sRmnCxu+4M2fHyxAbopfXzk05dh2YPGi7/g+afm9CtlCpfn8mVFvNTWWlYFAh5t2HVEbEy
voLlkGSs/gxeMlxAHOBO3c0hBm9/MxQbebd2QGThE9hh5PQaotwV7LvstNPMAYyiloWaHWBWod2R
5UNQCnVVOiqd9pYIF2h6sy0fTKkvS47bf+Zfw9lwgAfNvIchnMRH2yISV8Y3CWrFj+0c/K3yxKBc
oHJFmTHU91Ifv53ruSvHh/YM8AJeAAl04j6+nZfjRHM7/oVS1aBF+QWTmOs3L31Q0L/24fjQI84e
zKLuWMi7wA9yjz3GeRaA5IHfR17PJwcyqRuuYPT4rHsPlRamZjIMgQjyb/BrG3n9yXGL2iWq8HMY
0o8IEPNTXpU6o6+b5wKFTOSkXCipGvasD1xyopFHy5YMkXEyc6cebMdWDemGS4CEPubdhB+V+thw
pzsuG0D18Aq4pvoXrgmDa/OOasqWIoY52JHYiQw0xRAD2aD4Ffu9vCxsN6emmrOK7o9+Xy7S+gZq
WF0ob/X7iaOB3s50q5KY5dLtv+p3LJPB5c7XaWGkGelluLqdTxwoGa57hXQbfCIS3BP0jYItwXo3
2DqKOkvwhFp0GfIoF7GMUfWqj5xpfYhCRO+DB9u6VNwszjg7CI4AuJAzZxtekPswQJwH5u9yWbPt
Vq6HGiX1YDe8ApBf+T0nTS9DJYvsDd6nBSZtc0SvePYG6wlSoVLMnqxI6YAs64IKhmbic4Xv3vq8
Aum3i+0TcUggSduGbX4XOB+ZbHEmUNb1r8HGUNuxFMltXD+YoqjPgfVQMxN3hFt8rf7SztjiTVPW
NxqUSBux6jKyDloR4BleyHKxJH8T6fsoka7cLD47p+QuxB9k0KwhXEwh9/HlmCkjTYugJmrrFyy8
e5/d00ACBs1JznJXL7L3nupRnh+WRNGqW4j9nEinn/f9WjeO+iX06ujw5uMe8i0Q3txfv6DJHeB7
3WtpYYHclac/pfurkc7EXggTUfcE8P6D5CczwRXxGh+3cSgaXYY7GaJxqwhS/6I0t6n0B0b0R4xi
HZmyNSlURvx8I8KVhKRP3pwKvkVAKXVeA3uup9gCFkdxJwDO+HCUeyxTqtlCO1gZDlkNe+cvXIdJ
atmZN43TDkSfQneHkyNAkAZ307B3gq7HzpyhO5UivfjEX6UynPN/+6Go+BL99DDKm5zKqtZVQdG1
jdWbWHiTkaa0ypWNwsOiOyciDjhJbI2jUkfs2Tfbo4hzr0uBwq1tae0yi4itaqV0bf8tAzxS4csm
Pd6hMOIv+D+F7cPDOiAXEAdyyoKtSx+1ndFj0I+S6IxsNCieM0Zbtl9VQZkfo3NNSPhXciQHE2Ow
DAHP79QABSh8i49CRu1jZQNWXU+gJxAbnM+1J0ZHwRSmj2W5t1kF5JJ7Fx40cxaAVajYW1Zsugqg
yRNBgk0kR9e6rOb/WRryM+5TD7tvFGmqA3Uj5R3mi/ym/4A1+VDp85khy4D9Ix813WSHQVBl3mYC
SClaa77z2/ow9FuY/PmL2AjGfKvh4lcFAYfleYa6qORK5QTgUhIDhYX1rrR9DOovNuPZ+oY3qBuL
8JVml/UtoL0CYGffdnDnoQt0Dqt9HKg838VAA7v7QkSP5tdcgf6FegtLaByTKcILvrGaz2woYUCo
GQZcVvzVfyIUrndbAEAps4wgszJGvHM78grgs0yA/4LzjdllcvKl5UNB2Tpj1BI9wzf2iiHLk/ly
Az32fO5G2eg9XP0+Xg7EK4qDzbMLVL+wS94KhVhEg3vbjuCHY5gJf4jXBveSRQJYGNGZiwruYmOb
vXs/mOqyvvvKtV+g58vrWSY4GQowZH/8F+x9mVdzQWB6EHyj8WNwoDpXrMsbO2885N0tqy5g0y4d
6eJWkfq5CI8aIZmAFMo95ti+2k55NNH+dfIsiF/MO8+LFUbNbUl3nQEdalG6Hfs2lWMityJH0yxS
xy6xZC+e+z17uT6BEs3po5+X5T2sdedMUv0xTDgtDS6K+Oh5K3VOZhgIxCmAT6JUn1Via8oUDsre
HnRR2fdpnbtbViciM0wpelvnHTGA70xdXCL2ejikuXF+dFDPCE7KuUCK4UPZkOHPxsIeoGZupl6v
rxYX3Dxv23ymeYcCjS6AsFLd7l1HbEvLYuf1/NmxmZ2VQzTBhrnM8YQ86Rko8VBiXNt2g4jeDFQn
VTF1FVvWHaIkqfvxOot80EKkoM+yAm1kRzbMQ8G7PNJxrqpUjgrmxYefHbE79ft+4m5Xir/vqWGO
9HHNsR/i7BqH+g80S2vgi1gQHFR0BgeBsDymZunJnsZZ9cH1BE6JMYjtYVkMh2fWJ6wmw5fM4dt+
dxSdS22afhFNGRzR7kZuoJ9DOxBdat9YKAB+X5KndTV0Mx1zuC3udi2lpghzS10Ud6GLV5hR1qYt
W0jmjRIZ266GTDAiPCvV+nchQ+AL89+Rm5yp53YGjn6/7h5onbu11oyRLVnceL0jTjYgM2iX95fE
5lTJIuhsRO+Ar3gXtOl4fQCEDC9/cWUWWBUQLOl4mKhbax6Ub4GFBMfykvPEolKettzC0fcn+b1J
kWdcZjxoaF6QoGCVpNUvoXRCLpz6EL0a8kci7quyiwbvC9X1D9aG8RnqrXoGZEbHw1RUdZ+rYSn/
SaVFZTHI73GvHDXikGaMYn/+aG+QVIjGtaIACWe/zCoQhLenonyq6VDt7t2P4e5eZFHbG99X5SWT
H7wtQVRPEGPBccRk+qyFyisspJ3JiVQ48oajzQrG7h2TlMG257BJhkcRdlL5Eq/lGfZieGSkUUdV
aLwPfV9gCRuE5/eZ2dcWp4kulTLigR99zsAtdee5Xe8NwXKp+vDZZIf/DfS7Q8/NexKeAlypBJYQ
jMQuq+/YQAcS4ezEXcyJrQhfHFLNyUfI7fjjQWBJ7qWInOtzns9huwjDbqGEnqCqnQTUz1SEWAxJ
9efZv1GnlE4r5RcgFDf1az3bIWrNx+RrtCiJhniJRXjBM5SxQcdDbhWCAnvV1NRiV9mNxdxVmx66
pxUzIM+9dMriZWik56Ar0yb7gOb80/yL3fSf078kGRJ7XioqMuJqmfNtv9mVXOXzRmRZrWI0rZlG
1ai1+Ux+CHa8fecjzxmIn6YRJIUKTr6DqhZb8USSsE8KRJtPs2r5X1eJvKfV5iZwHGNzZ/AR4HH8
FK1gEkKZQnlLnGBrdaZzv0/tSUzVu7+fheLn/W5RfJYbUWQ3YNlH868ijDetep8RxbJyXuCd7zPq
VKSngQPdjQyd6Tx+Ak7zoao6+lQrNAGHvd0KxZ88VcNX7YCGsSikexT1L6Js1v2druCibMCPfA11
bzR/lQSUwQW52HZY/z0a9n+e1S2B+azshX147d3nLOoTgjEqdmqd8+5IdPxAaiooKX2Vj9Cg7RQ9
STPs7ke770hxyl2h0ksvebMd1XxcO6PRGvxV7mKLy3kBrB7aAatnVS6eIYYpsggmUEU+VF/1+qBp
/IhLyfwLErLEg+PfPuCnjLsfBcpC+LDHtioyCcTbNH/Qtk2sBOk2sprFXWrD+2F9clOGZMoyqS4I
YKBcXZILtorhgyBsTrutWLykrmwR2GaEMjNyOJqIHFeo4adG8iVNSJReseWhWpeHCurItACXV3lm
T+LVTeEDrjdScViKoWIo1V9aOJzQ0i5ffPfYTkzFhUjEIUeQgPegYMrLQZd2KHBxRxcC9uVCFYUR
QMIKYV9pmsjEEQT71VT5XAFUftY+35/ss0EE+ocVJdT+aw2yDmG5uASGNkCnb1Xmw5qrcJyTkYa6
Ot3ZHSWsxcZ35NcF7Hk6UO/hYQe+DRL9njCEX4HYpz9U8J8yHy6M3WpTBXI5701u8uIsUsQeQZuC
o7A7QdPR0BSeKoBHhz6G3Z8UN8HJATe2l4wGXbonJIDJvQyHBB6wijwxpcigvy2uskY70RCXcFRL
nyl3jQb4k2RYZM9qPfrSwo5Onjq3SPhvfFQCr/8zxlGOCGnlsyunY1t+yP8I5busgQN44GG3HCPM
4LoXKHfZhYh6dHn8iLczH8CmurJ3dUPIBpxdJOSptzQ2JaPf2nCAu2KeV6wULZZ+Vb953F1rAaRc
MJ/3FVUyBW1RoOuP5LozK7PgE7/hKzZHEM4IE68aU4VkQgLg4w120tzX9OQr4mGbsX5oPxdGrSV4
07pmVBbrdUKYOjUT33vMQIQ0Q8pjkOFAO1j+Y2pfIw/JICapMVhcyisCZJam5+me1qTgIvPXD00I
+xbIO7r/QLJL2Fpd6D2IlDzI5z4sMfOeZA2DqlZFH47O864nB8Zh2FjpdT2hyv7tSiuVHelVdw2n
aH2xg0aDVonqsexlZTDU7X4Ew2mlgBEBWGBZrjmilIHKoOCZwyPQJOlUcPDrU2fyB3DiRMr/y7LP
ZZX/m3EZ/q8sL0NPJU3nuY0TtLY2mw6ceSdfvNK5java4XOX296Mtk8Mm6xSaxQ9Bg1mi3quHcHr
6nmT1G3NGFKHUsRt9Tv0bwflouj8C/vOd3FNYRcSh7rIyVO9ZAMovhRx4Y0Cc52vQj3JCIzjfrEu
tTIoVnTUsII5cKpWMYOzaUFnl6QOr0YdZE2pwuEZrgmP23I6TCcmQIZMrCB3S8DcSa/ucgK789tb
tO3HnVPD6gHP2Vg5sbotvPPMbeqWEk6IaDkjhIwbJWvqRLkeZ2pXmRF0bO4Pq9aTDYLuevEGM6Mt
a9WelLXLwfq/ZjNAbpU+JecNo7M82nyH48/4322+xB3e8fRWSNKYdsJNrahfys0mGN43qteIVKYx
E5OtUFKmswO27BZ7C18Mm2aSewXpXyf/OFLd0nCKyX/u+FFpeB6OrdbIxgdvIpG3+NBwU039aAQz
pBiO4VWs7kr2X9Dzvu099uL6HQcIMVLJey5YsCK+wT2cTCG/ZtxCYG79OcXM2MUlUsdlSBozE2HI
0W+WeoQX6ckVwXp5Ft7kjX3+7ux3o2U79ulemI0/Dk0C8ojg+g9IiZtkj7AGYonAOTZMtCwbazSw
PnpoTfioN4I1TVE4PJe7XdAKPG8Jae2yVLsIq8oXVhQkTIcVpdxSXfLRKFBb78YWveFKxc/RufGi
yGgFGmY0HCnELTBmJ7H96E4lOXB+1hbdGR3R6IArrlQNvSvWdqI6qL++w68sLDVja6EkBXhfovmj
TslmOMwRHZLUmXk3z8P8SDQS+JTs1ziW1nlr8w8FihX/TKCjpkSi1ygZuuWF9jOtgN782MWrGVTj
HnCBB3SfOFn9yzTQ1MoteeRsbUO/JivU6WLWh3HLIIGrHvMQI1tkzkZNkhrhT9qe93zISo5Eo8JH
8bGzol/YVbelgiIenXogAAALbLirYQukujUjEdVe5cDtFzn0o/MyrBo5b1ahHdI7OtgXg+c+I9d7
H9yw8iLtB+PQp4hHSTqYdNn8De3zveLeDdc0aWcEetGfoj34YST9g2MDjqhSZcsK1mRprNfJP25y
9XgXTQj769YjMFQpOSgs7wzWfXSfkRHE2n01VcK6QxkJ5TxaNK9o1uwoFZovJ49Tt6bGZXbM/3uM
fy+eMt2dB9GAeECm2TXt6i4PJb5vBXVusTXxoNlI+WjiSlf9jTTE60gtMm+Splg3u0yF6Ugl7WDh
8pOcGlkyquI6rEYqZrtln26/TQn3DVmNKTrqoiMaAaTxbCCvWdo0KJU/1BYypjgzn3KTOzPpbIMD
ieLnrLUnxzau8eiZbZWeV7ZKSGruRSTiBsel0s7JsNmMQQK/wLgwTZOvxBAiULzaQbm+jQ+ovCHy
o2ZxoHEGfvyO4/aO/0ucmPx9mfO4eOGKVJxB+lqM1UnYOmD5l0NNs58TsMduVf3stuklN4YEm9ST
vwTAvSMP4z3zcvr9aQCv+A+zhDH1q/hZS9WZnnugA4b2+K3mPmNiPS/3QpkMHZiRxXRZINobgRZd
oGoBQiQjzgi5gEW69v02dbMtHgZWcdJIatpkUz0Ppdx+Z3qBi99RucJ6WB26hWEoP6irt3EJsGmM
hcG1Ynql+q3HOPXiMtyW7Ni3FLtTQfcB4kP6xWakSSIv5FUatKm1NDG3obX7lQM7FxNtH8eZ7Q+6
RFtox7XwCs4qiOsjXcEmeB2rYB6A9bBARLUttZO39yxt1fNeGvz1ZRuZL/gN67fSoqLf3o2L8y2o
MVRYwGqPfDR4DQ7JJ7qBsQ42G6qB/QG9TJCdq5utLc7jj/qRJzx8LXAt3sxefPNwzA0dEWeJ8O2O
WngrJvVBrWydtvI0sr2F3Pt2I3gKCrOfUP+XecT47zif9mLVIuXtVNj8B41FwVLSse6rWAk5Orhu
pJSwWQXAxrHkb6KADM6lmC1pPYnXQ3ac7kareY3ET5SBgE3MwPD0oNvJdxmLz9i70wg0it1aZRcU
/2wYY1RGAZ1KgRnnpbJzxARTN8Lu7YGs18YKhHQUtCO7TdopYftKefoIQyPa/ukNgzpGqp4Ys0HP
NIrNj0XybrCjWQa+DMLsF0+klI917SY9hAYfIBy3nShxmNfP4VKGRTtXPNQ3VsHi2+6KOox9mbfG
J92vWLLYd9eBuYjfNEdasvcYSjR2f2LxupJxMwT7Vp9CzOJrxdKfGTmTxKVaNTh+J3GxivSP3jA3
WnJ5mHerv2OczuDQV0snXURxccftxlcWy2VsxfrrROKRONjt8yCbFX4nRHGUdRmXS6tOXXN3oqkt
c0Tpx1qVr+nc5Q+fq8+WY1pbvQSqcOmfTJS89cfZYT4YWN62yfLMUC2NPkrmm+H124vdJG81O7cK
4Xko4lTtoVpLu8bln3KyWXrle0QMIKrPTHrd5kuxf1IyGqcdhW//U0Or35/cPs6HiulWfGN+IP6E
nATJljjespAOwQtq4AxWsdgyLDkdzdyD9U3mMyVVER3CN+JdQ/wVsy8Ogg5yqXpWKvvvRc2av8AO
aamagg7szebudLEuRnU60cF3kReObydPOmOQRUHtc6MFJ3Tq4ysdb6YA11XzEm0exNqSCA8Ni90d
iES1KOnTrZzhdX4RaVpNLDZNGeQuziv2CvArQi6TN5mTLSHnmstRjO0nOs+UM3H7GKMG92TG+94O
V/7f1aK/+6UQqs1+1l9PHidbAf4op0A/fRsUJ+BLvBUy/UCq5Sflg/9kYqftQFmRrwZMLMImCGBe
b2zQrRzYJYX7PVWKaman7AQomYCY2a8c++Sy4qwfgfMJmNW7TYQhqJq8mEPqy7MzwSCdTYCEW/+v
eH+SKO1XSsPLmRDBMri0l7q10RYZOMZzTDNPVETUq+MvHeGn49zHc0xIjfI3kQu7ElSrD9n0MLpF
TdUMbXOyXh3v57QwDIyL8dIbgr1l1hNcls9bOvUTcXavk1MmhtQzSXUs2el/cF/JgP4IvOB9/oSf
Z3SHcDL3D+18hXs3UF9RAnKj8gckngfogEWO1J4J3JFDdDL9+Au1wymPWPbjGzxAylaUxObhDXKP
y5G3zDBkqTWz3ayspg5botpNR+uwf8prJJ3eyBB8Ll/SqLmZgHSbNvx1XuBpvBbM3tdb344s9Ldv
aL+BB6jauDXUGqGZG548/8Fa5zYsPTWNO+QSIZEPw2A4QJsePFEV72kmP0kV9qkVkMtxltb00vXE
pzpTVwewTkayd7YIzQy53tUpDX9ZXYUIO5k7qVWGKvyY4SmbVDE3StgqaCnzoANlqL3Mwi5yR6tR
z0my4PgQOKeFD++Dq5iM94PKvzkqU5JZLGf/PWHvxQ85F3iBTxWRlTxRrinHCLdhZEQMkQQ4xO0P
nnJVrTrl+OnoLqDVLLVAn9evnTto4b7ntQa3s5Ps3TI6T3PG8AWpsCneW6GkwDujI+yeSf/C5MFD
3T16uS6u31TOnFbaFQS2UjFERSAGMA3gwftyZoAi+66ablHejSRlSlAz8zVjNlqN9Rt0Re+9qe5D
+0L1mulmLlILAe88qqgjcGmGT1E95KlzaIy7wT+VsFljeZ5U4D08DEB8MJcrwJowgHiQcQ7xIE1j
hNBKyd9s9EF729c9BCXBkzBNmn/3Co+CP7FcWRfCXBBDFanflLSVXQQhkDavaGaQSd25gm0fP/RU
GScayYu+6tE0uyYMoaYSECUzufMCJLs5r3gC0rBD9xafSYOVg5Wi0TXdPHKnXCiPsVyuY+OpCAKX
QPCnd7n/Us+4u7xwkMshJyS7tJfD3sFNEEEmoNicXeYVl+xlKZHUP3zgeEM4iKMWRtbCU32ENvrt
ualeTHZ9K71PhEviJA1Hn2BlNl150kRztQOKLLOHGigoeNUzh/axSsyqAeeXuHiue22XSWun4ZGk
zUz79TaTEY//rAzQfejHdSZBJwBpOXGMTELoDG0usyq2rEzgs9rGOs8gP+TFVhbEvcEvNTI0Zwke
8OUiuX3iG2gLDpcEdDtDZRXv+gtqPluuxMz32rNMKZfknr8n85FvUDSqnhCnuGNH3Uo6XVJ4hzwc
o7OUpqZFl8n/zuGodqw08PawhRdRPTfh7wargps+N1cIMcM8rdXEQBmbg7CZmQPZ0duw8t35Rgm/
6BxMxhXbKLiCMq+T5O6tEauDMH0960w1kHEjCfzuRrJ0tOVdHZkEN+ju9zQ00/CNHU0vOrCMx/cg
y8GUCBB3l67Mm7A18onZZbI/n93hq5MbtmRX3+CTMqArPPIdufsPUtqXU/caTjoqPe72nEx8HMCI
rMkcP9U2CKOiydBGAmw9As54hHCdbafaLml/BEHHC+hLsi683vtNVxT6tdicRWckwH5JFj72+Pim
Xex/ENN7JF46OF2CsOY2P1bP639D6XWRy7INssQ+IANzWxi5gK4biA84Kojmz+qakmCTm2MSetMu
/I7sDzb40+9R8OFDnpt38CpibplSIVOpnbhgsK7U3zlSY4PQesw/iKfu1F0+DjUDCDMesDbMYnb5
sb8QbZ3ZQp67NSX+DR/6upI2MK3DPm/dbSxi84rfHItrSUiXBijOZqD4BO+2BcmbQFORWQqrz3Rk
gFTGeyDTNRK250dlOQctXAqEGtDMHDymVDDOONl2iaJcNH1wktbFqWV3yhezSD4jSbXktBzjGepx
y7vSDU5Jdt10CEcgTr169LlI50iepBw+6uuulFxAagmqNHAgTmOrv1VELzuJY2IhPXriymOVG+MP
Ugai9wwimWhFkDeaHLdSYfmfsj8fhhD4ymEfqZ1jVNzadC61lvFtEAKnlkZEloTKOcjc33LKerG1
4IxjO26HnCyvSe/PmhHpWB716NZy9SGQfg5MdKDsAhHUrLIkvl9gupWqoP21nZyzXE9+rgCY2oi1
14PBB7TcoocJ4eqAK0Q/CrqC7IGhlhrLuh89qG9SHuvmRO6VNvvhqbLItMRZgEFi3lcNODdKK7fh
UeJWpmocGvb0OJv/JTds/aoxEm8GW0AoejniF40MGMUD3iqTpRtC/vx9o6w9ewJ/KvhjjyrjLwnY
gwuUUSQRUmTNGpSzJVo4clIMpbjeM2Q/ESWbtpl5IM1yPVKNqoNszh3kkNAG6edkMydBXBsII3Nd
J6Og41B7Fz5Oqa9kmqhpITUIcUACr+OisbLQA35iZPJQdMste+qLQLHyONjEufPs4qQ5u60iTIST
sViUtyznM+z9zC0dr4d1zL3Fekq87JC7dlYlotkQhf+9wEjtMk2XQGcOtDQ3GOpqOMaHzWS3JldK
kMYisqmbRZ1jz+Z/We6H606oOxgNof62I+b9d1A56a2EE7OoXZhLFJuK9bjLn4cy9z4CK1PwHFyI
xP0G/EaSiALtoVbSB1vG9Onp4+E++s61qf+bx1SYgcf4maBIHYTGLfmWtN4ZFKHa3txGDGzpv5EO
kySsFcXfYj66DTSyONe7x3P4Nn7cHxQim7belno/hSLWhvam8WQxmF3gpF4JT23WYp5Qjs6AgGVr
/WPINGciU2+vj41fGeT+PbkUK6Os08E8rO3kSnXrButnw16NNN99YmWpGmMrSoYfKJipDnGyuUyh
dk906SDmib3W9soVLsfIWh26pjQ4oDqeX2doLzjKz7ByVm4aJiXCVyhUakDPVxxUk9+qHxlKnNYJ
fGja2yROizqYz1Cx7KxkqFbreHSjr5kpF7ah7lq6amTH1WvsaryvsONCqsHeIbPcxtZEMRkHw0/W
6QxTLNTWsIN8/6486Uor1J6jhRNpSJS9h7MjaRlHN51IKhC5uY5Msl80igyyitfnArV4jCO8yO23
hT6ZqV2YUeD7fH7ZeT2W6lXeMO0jwNB2891R/BO4Ov/d1SCKTEfPhtVPJAYNCwsxXEBh37lvBpPu
pLrg/VzHwGnZFoq2HvByKyXYpBuOP4NHSJqmVO8RdKJtGO1r3lH1H3yKkXcaaLhx0JsC227XA/HB
fsGgOBudG5870f2iYLC+sSRbEIPFaNmlLVDpm2n78ATz1ePs10HC6K8OV4lsfgMBWTUsjC3lseyv
HT6mZKMn+N8ogOfOQ5Fxuo/jfA3/fV6ndWiXAS8pQB3JO2GMfU/wl5SZT2Ymsxfm6x9oqUeoWtAA
KGwFYDrxxxqASCAynwjd5hAx+LU4xqGS0AIwfGy07+iN/UQjP/mmiHxPMFbn97bWz8Io9+NWzaQc
FVUIqbvaHdrhS/qlvR1acbLOBIXG3ilgbZDdQrY7K/3lJHMuhpz0DJo/gRmcjAtsnlALGVEcSDgL
3ie0puvt8BQtnPfJ3mZUuiji4JwSyU9LVqXnvbnojG+QcAmQfoaCMDXilxWLuFVblhZPMhlUuRrL
wkbfJud14kGR4pafn5vRifFCBaKl81ha6DgdrFdrrfAmZhO2NGOGlsFdts55H5Kaf4ULPMLd9uHo
GDhW8oPXM8vHvK1JGzNhtGxxlQ4vqKdQQubkn/53cf+tXa+KnPS8Bd5mMftKq4c+8sNJKEXREhu8
AmR1LaOXvHFLTGFj0Y7WGlt4ZiJ2vADqnaf7pslftq5ZhpjhSD6AMVwQaGy2lLiSktN+Xsx6+eaZ
fBhHSdVlf3S8IKMp3bQ6aKjTtiqjEyh/Tz0ArZP1+zuLPVawBC0xaKhRnhT/4Gb4ob2QGUari5Hm
Hk8l6qQxltoVx0/BM1DaNByfjOyv0WCV5xzJY60aBgUn/y9q1yLjwbhLBErMMlN8jeoIB7n5oYXZ
8+qL/7gqo7LU0Rl72hawDOU4sRIlLLCVHWL2sSK9p/lfzmP8w4178w7wzQNX79FkTBdlXV5WKe/u
sCqwTDSt9h/K6PLTn+rhYYjzncXkQRNMDOr4qsDQA0adxgIDH2M+7QT1TqFzxkq5ugqB7XILZJBf
qmTO7Qerk9eFsCbHCowVX/4Z/ARZHmJjF4DMKYPSLJvPrFEpHPMzGK4WtdTTTkRhOO1YEXlOLHmd
DDoKfk7aLRJiy//pwkpWLZHO7aTrgWOzth89huopVI0o9FqoGnu5Hv+o3bm4gakZCC4LgeaAHZW6
npZcWw3ewaL8InhyaQvo7ERk04EHKQRToO3BzaDYveBCxDlwpXDqerhZjRJ3brH3UhQNz8qyWIak
69PLTW33b8hnshsjEfIeJ1Y8VVWoarTSypJMFGk+EKcRkM25UFS85UBW230Wo3c6KjtYJRl2f3zj
ha5tNdVjHLWxAnUAd5lxzHJEFrkRZjRybsqFPlLaZDryW7Acqhzn0lLtCG2lMye3pMqz9OkdoIc1
R3DUWJ+R6G627uy3rQJOt1UMn9GVIKz0ZmGPdeXIlnZyGegsZgMQq27BpA/sqVQtvI8eC3hNMO2m
4Xmdy2UT0WMH3tZPz6cEUCCqs+UC591deRBkr7M0STyJM2JLNWHR71Z2JQcAZuaT5MRciZ+OGWhj
nNZXeapQ/2u8qh/A7Sjb0sc4T5BT5IYHS2FxCe9yMO+Lm9AZfEGLpgz8SxX9b3xylXVlEZbPSBiv
mnsd3DSWJ7lCYBG9v4LEmsGRx+m6BIYc/pRXQAA8a46luy4MW/dYFgzyllfmreg/IqQVayBpuOKh
TJulQEkznRQDGXVA3XULq/2BrSpPfBbVOZi6v3Y1VE52ltv5k404N7VMhGH+FnQC5om/mMId+Ms1
6Ih2BqmS5eDq2i/mSaCsht1LuiuCkHlqd5z3vMnWn8d/LfzK/Tph6hjjknXi7i0QwuA0giKRZQHE
aStJuXU+kRFiuGjYRlkVk+vaJDBjNkab/5DICt/omekqeXHJFfjKHsXZdT3s0HEoSMX7N34kvIim
6mhQTuqxw8Sk+kh6XXeODinAhKRF8yoyg9+IldtId8gL3xC3K6LXp2W233hxCFZ06aCW+4qzb3wx
tMLya8X6VHSPs7Pxh7EDktaO/5urZsCQgiIw2EJM5IgjghQMSB7DRjDpJDkLWX8hrT4+oUpt3Zo2
RjmNmzO1VVfGu8CZha/Nb2n980FYmVbSDG7l+iEOx7foEAa112OP7cjMEUEogjrobsYsDW+Da4QI
bEHNDnbNvQ2ETs14FbbLGuwZrJei4jOI0Pa48XX30PCPYtt+1M6T4sil8Dx4ok8NgN4Jxf+FFc9f
2AkRkRM91pz+/weL5woHUQvNApnzX3vD1BfxSk3mmTLeSu/J09V42//mPlUIylmFs4CFvWI6QYzf
CrFf9eIHL70iiacCdHAaqb+koNfxSP4YQ1cJ6A0ee5txr3L0glBw64nlKH9tkb/osIIsxpaXqL3s
NGgzQV6Oe0ZnyMvtqorn679HNaEi6KXNFFymTRRbMcW/TtxEbOsObd/voJvHJS18sJz4+mugeGWo
14fIcxZmFRd7qofFd1D/ns0yAZ7WF2Ix5+0Qby+iNiFl198E3OT9EZ+ue/AXAoHjZmmlQpD1JytZ
tpmBV94EewSzj2M+N1Cd7bmItCUIHzWAatH2vKfy3NPEpsCZ70oqyB+YdR6WoS5ZkHDtPST5yttl
1Dkz/r12uQ04ucCnaDYfY4pZeeIc35c3nXY1xwxPhQSsuW8p38yd9a9jTa3O/t+7kHCAmYCxfbhN
Eu/l6v3TCWZd3aVJx0PYdosp9+dVBlMoo5dJRyK6dTIVASWR0savR59yaYu9bXht65C5DcRoCICm
uIAFI9BXr3a644RpLR9S5dszVay7FfXYz+nBlIv/OsobImC7IW5m2VHgVzUxemj+Tkik+qWy0OC4
qtFEVTwwpOdy/FT1CeL04cbhWDPuXfm6YFb4Pn+QhoGR/OxbDkBYVMmP1vzfUPCuqR1D/3t0DIGm
6/vCbr2g1rr8zijlR92gXHdWSwrtDUhRTtC7RDcIoSyTCC2EdpUqQ4nG8w6jr5p4QphZ2C7wpIje
yCjCT3jg43m45R5XuNzM2TTwCN9ahA7AIzl9P7tvFBIFGLBAriD6xY6TYMrcxCLb7Q0saVg/wZE7
9Qn0dHR4b/Bq8sS5/z8r6CzRNMqSBwf81bi0XvWCqZkFRkfcZoXh6CCAWY8wX/nr4N5tv/cJ0Msm
xvxc5BF2Pt/4deMSLXvfdYWSP1lRbBMMyx1k9h7zXvBI+1lqSAJcWY16DKwxd/9hBTBBj/h1zAD+
Avcw+oMe51HcSdvDCCSjsd2ruXNWN0+aQ+doXzwFCg5Q+5B4kNYLwi11VNeAV/ES9hl7VmX1ms13
svsQNnXJvcwQGaepUQ8dgsUDBLM+y+475y7l2cZZ7V1Kmxce36+3k74Db0ug/OYAiMryIBsHPOmU
zfBrU5bcWXcGzcAlzXIfrDQAgQoZEy2wWPcEA7Kms+LsCPfAf5o0Lh1WRjRDLHuwbhW53VDD7zUP
iQcWZcI+yPX6ta8PGKAFMjJ5nDG3y7Ns9JshsF9JMopqp2IdGkDCFotQvYAl7ut4n2APk5OYzexE
T5Qv6WSy04EH3GtKTuW0RFBLkzBMGVnLg5MKxlsvJaFP96M+Lfxz2Oqgg1NKHT736IgTCrGTW6Hi
9YAMynA7yS70j51KIz+Qg4Dwvs4m9lpfe315FApFKrIYgeRb1UDnI9HnL56p8+A9rmJg47qS3IfG
VT7RIa+qEACfFX6BoHHExHsINtoAi6QmfAwM/uZLxB2u1esbE4HCQL/d2hLxNYtyQ4A8QeH/sfS/
73g2osJEmJGD28u+qOGXx6/9XTZwwcho+Sayijad5+pdYWjBweb9WGEAJiFB2GVy+7zDuUmM6pRX
OBF5lvOvGsH4SlxbykRS6Tum76WorYOAQz0Wv6FOcrTuuI5NkGQIQ4d0r56YdMku+MgIRYt0YTXj
yje1AKBByKuWm1YVMWX/HnK5Wa8S6/TAeiQdK4kTnxySdG7POGH92jja1dlfjZOW8R0yy95xjocC
ZSoYmbeMGJMOHfIVvQ2DBAfsfmegrJIBAwCuVzgp2viCz8e6fvzbIvEFK6E6rgsiUOuSZpGRNi4G
NSWLQjw3fva0N1COlEeiJ/pgkGB6yOfzM/M0o1LNuq3/WYW0A9Htn+HeIsRAfYFyIqXWaWeTOi50
P/6xjIctz4VtE+4SyAXx/bmSu9lhslTrKNyv167nQJL56I4ahde5fvg2xCuw/fmX/NXaHaCaWl8c
kvLqJ93ViRZhqq9igfK8s7VqEsjHL1Aq/ac/5mNw50vfxoj9EV7xUbfcL+DhiyDTxbsaNFt0c5aD
oRVACL+tFX8o691ZQj5lo9RGAiu+ukovEjBSDkq6+ZTe8ao6EozFrxwnPJV8vhxuG9dJcIy4dakd
9TdH+WqGjEVfoDIFh1egqfJTGJ1DrXnKLNt/38edmdgUZP+ShbB9nkwuBHlQKC0f4GIfAEujKRSH
RQs3s30DEgzsENidu7gsuCmkUrJzIhEiHbsbtvusXQ+BKtvo/5wXIDRFoRij9M5TgmqpA6l8jTNY
/QJjI2N/q+L59T9FSru7nrUqM8AlgN3p7crzt2mrcL9NwcecUL9cArIlB+7HWMkJdv1i893THujr
EDU860P6TE+VsmyhbyjalGnKE8YUjcTiUXxElKTEzNYckfdugWhqLFfgvDCKNln2Q9FNvrFCZoUl
fsKVl2Swa5HOmm41QeThuRaxrTtUa2YFYWo4AKWxGnz9qWkDYueJrKwBaKzGahfRpgAEKHi7211K
GXsaKVN80LEb7nJ2uo1eTCTygbSipJSgtJnvVoZ4y6+oqnw2z/cYq2A3DkOLOzNoi5XSh3ObxIfs
CWKqV88TkVgtjZ5nqVFFKkQtTH+2f0mtX0N4CEDoD98zgyjSmHFaCV9cnvN49YadQxT3nSMuCIHX
mhSwas3sJYBuhcre8VPCibsyc/dPnuH0cufKRyoFoEqFqF1eWRVoOdeXC+u6DcZ/8gW7W/pKsBmw
Xju0/q+ED5fh+jYe0teW4H37swxlGKxhVL04Ez6RfUxpOdXG9TphL15jnDwMA8M05zVElBIjDksN
Mo4z1ppzG5ASsVeUPycQa6lWxgDg6fGuQhetARrt5esRbrqSoqp+7qMmfz4xsLopASdg87SeX2Lg
tAFgws/ORkwC/czsI+r9SO7psMcQl1M0aOuyeTQi4v9yH2T45EMrNrl5mfsLH06jM7ivxeyuTTyx
2mK9qudHcST6uliTgj4kOmYUiVBMe1j2zRlUYK1pRbN+WD3HMDDAQMgPZjqok5dAilML++kk8oXo
JAvOcFuytOZlMdP4PH297l5obwLeNqbCCmUAfpBezTcP5INUhIh3WmmJqyjSlxgVKNYEgKJ4CiGp
9NAY4DPzFPUZvStZuSsFYmB+bquH7IL2oKTou0tBX7KKlNraRy87SjicDPhSV7Y3yTyN5Xo1mg4d
ldH1VZHmNFon+rv6Q5HZGTMIbD7y/GPPljWpI7tWDYQoxa6o46OtAVlH1ZdL3D3Yllfz7mh5TjxV
i+nMOnsn5V1eEee7yWyKEOPgbabfB2kuD/M5xytwoxMskFY01ggi19f5lElwFWPK0ycyExGs2zkA
VmcvFSzGXMmEf9+iRQ+HwT77GuB6L/sryS+23apvxYJbN+45zm+ihEvi/OF7X/HRkT3lwFFNRJXr
U8BftnHQwMqFU151mo2eB24OYOhZQ8bOEIZQ6S7A5YxAOSF9nZMotWazA527zdE1ap06311025ao
2DmB09iMaMD7UD7VsPGxeyxeZsp8oOtPWwjI6gazwJg5uh1S2esTWB6AZ2SY+CnoZ628oB87CNRG
7+Fbv+oHgCQpcrg3daabE6RhQDa6AJXHvALzgYs60DYZMl67DYrLKa3reJGPYEGmq6WaxzEVHoJL
/GjGURYQPbU0rmzvXMSNTNU3RbE5F7IOFlycmoZmkzhoXkjVpXFCqj8Vi0uA42aNpALMqrCsRTxA
QZOrMEYkO8fYGe+HkKZRFtrfQG1PG9btVdcDhYQDOK6LaQ8NzNpnbFbKUgwTIzipiqu0/D7JEnZs
/KTIxFGtFO7areWmHnihMSCYlsAF8ubxsoCSLVfjkVdY+WuHoowWeBM2ptPkOWOkWA7KNwhWhzuT
A6zJv+ebvU0Nyxh16OuPt6YyTMwzYQtSjeUGOP4Uzk4nJeAPsRYENOyC8wjvvafAKhBuCclZzOpf
2j0vbTFwTEcnzdaJaeOTCZKPNcS3UL8l61gmnoN6pIuSdHxOIhk2L6r1PGoUFfnm8EBLjNc+pHgD
BbekCa34on4DuYvt2IVLvI8SOqey8Ngounu1P5etuesBcb1jO/haZi2he70LoblVUyrUPlovDc9T
hSJb1GVLff1fVXI05++Qt2S7FiG+p6lfGIKT9dtpK6Q3D2eiNfmHN9m7sxSMT1x/qjcPvXBUhe39
7fRA6/EqsVn923W8JsgI0BcDJQ9h88a8++liiZV1xVcZXjIKVKZ/HmAnn9Soxt1JG5uzn+a2LmPq
we5KrEhc4dDTHYwDdMlRb9rbmrnO3JmMMK7rgczhEBLTLmX3ytdSdbiL3ViyfCViyb9BSgdRvUm1
KFXKBo2nyILP8m9KLVWfOgdTTM2dWDSptPdeeV3ot0BW2v8ZuevO6mLnP12HAKH8RKkcHZ+4cKAS
e60pzXQHiLUkZRPKekGTdHEzJ9XzZMYtHBmxTY90vp74ZXBhvOoYrZG8BhxI8vz/yIwDlM/XLdj/
A2Q/fWy3EGpUkxsiqXLmcCTuFWlo8JVeWFmZUkyRknn+d8+x/iiEYg/BtNGoIxafb6q9ZJ3CtkPs
w1dMUJHhM5Lrj+31DBy0xdCGh2GQrm29qqfvnmJRjUnf3TFx2Bs61enpSA1iJpl3MVV+Mk7SmjEg
DZmF3JyFnP6HcmomRfkGOUDTFJzMWuJCvk7MUdsRAKv0tURWwyGnMJFdsNF3n1TiQJm8dAuZvQ8u
h4C3+GnCnuHUZxPGs1FLyAQVqRz5urccs0xfwQNSYC650w+TeESbruuibcgo5KpwedewgL/B1/5P
aXL0mvrGMynwCa/8NCMEgWzJNVwYcebU4lWhQBcCOHDqE4L2r1gkGR7KGpn7v/uLjuKpdgm7gdPs
pNBckP9FCtomSVMjb3/R5mnLvKfgpW5XDo2QDrGkkJJOJuygbg6+uwA0cJowQ1ycZ7jmSwVMcDZA
jpHdt/U0nYVRDEKBq/j2uqMMu8CoKkAxdRJyqPNp+gWNBvnbICeypDYz1yp0iQo933z+6nBVLE53
PJbtK6z8J9EFLhmi/YaPGw1NLKf+kCRGgS2PI74Xm7sowDmH5Urexylg3rulxKLTiqeIuSuVptTd
1AYim9NWOgyTzfsODVMTKyrxQVdQmCxnuVH0aqbqxZ5nvDVn9Ot4TOR6wqL8j254VfPFshtP+ulp
VODcB+qBYdIgc3DB890Lt/aPoHnY42fs+nt7cSqIcf6kIm4S8HoLf5vW85atlmUpas5Y2gKTgoPI
U1QYG1D2uxIwPjwQZdCco9aEThYC7W2E7Gu3fj0ES8KPuub5YgbGWqopkDKA2DOL9ScY1LCTDdQz
9wXi6D/YPVEzdgDysVExtLuIVzNZ962no9ciaQejcgPxXhaKQblbg70yoH3BEkKcUxcF/cE/Fhd7
bFN9d7aL5UbP2V+FrrYbG/2U2Yf61rYp/9W3CjtDrcgZDDwBgNjQBRZx/aWxDsgTCWvWXITc+CCY
enR5HWLMp7GNZjchd8CLIFSK6ob2h+F7vwJ9Xj5ZCl1jFNEyhKsOVace4y44uSiTQ5Fg89/58iYO
hnaFI/44afGH9A+kD0/RoqArB8AKgORBHD8Rx2/OQCePH0YmSfhxuqlIaKVMJWy+5X6yYKNxQt0J
pA0eDpLJRfTv4hfqgMra6HlW9gjIvzNeevH9N2ZfWMQIbpY228aOQZmF7T56XyOLmYL0cHdLZfoZ
Tfalxim30hxn+HqHjHV4K+PqQTq7Ui4WaYk6w5vYnJmXJR0wSTHAV8VKTfndtaILfLjdO2/EoyqO
D6qdX5CXNDdfLiddGZzMxqZYxM7gnz9mN5dMV+cP/DNiPr266zu9XhrsYOsorpav5CxWWV+2UzeG
2NFMdougvtkG9h5edqy6p2ap1FCrOLoRH0VGlc8wJdW5pPZEQuVP7RS1S3XPal+9e0kfQ/i0Zmo4
CZiVXSE8EqTqJ/NjTvuKd6GQSo9is+GbPIeVIZ3TUxTZffI3BnPDSBozGxUYAj2ifJa+FDxbn2Es
301tkHW+i/FQbIdcNQ4C/BRCVjQzuGLR6ddi+RyNvdksWfkAyNOx6rRTGquNWcf/OzoMK9A1bpPE
q2YSQan1pMMDFKLGXuhmOKkRbU9FnuZa6usNlzeHYb5AY3K38djOS9bgIkbVMIzM+xmvE0InmnsY
EghAIF5/3/bq/GopTuZhjIi7VkkW4PcDBE8MhSdyU5YaJo88rI6G5jMzswMJcqVLN53t+qDzzDWF
eatXUga/LCS54Am5dvc6J4ntAKob8n8QypP9czuO9ltqutUaibLIFEqQHphqk5F7xta1bl8rMTtd
bzkGXGG/HLeUImaAq5vDViLB+yLuZpGeJk0QhW9oysUa8x4iIAyV8EgwgbbjAOb2a6gaJMo6ObNC
4mQbz7vf4uoOAJD/80ORlpAYqgliNLQeR+qfAwI6sUfhDou+ub3PgQEYVSDi2JjE+yV9MGqBKi/H
4quC+aMemurHvv/oA8UGSq+92Jypw8nXaC8l4oq7fyICLpuGmVCat0PC1eYsTsQUnlTRvuCj44CM
ceTOnAwCrciXIMJpxnv6poEXPvONEbXibZPtBfNFEbV2dEBc0mjrjpu6H9CGTs1fpZQ74eB6SEMI
G2a8EcmlyUhiVD6l54VPl6fDwGahlZeyYs4TjXOUDOX/CmAnn+2Ymuipdpff+AO6tGl/fSRU5PfX
Q5FKjIdjIM3MvQFjRybjfl4/p70Q3qeSvmkWkDu46kU8lqmxsVFglIkUxmkwZfjpDL7y8/KudOp4
NVs96R/0CsJ0/eH1N9795+aAY40ErxbYN1aXI2lrRBWkKwCSdo8hfosiZuIBqshqQVxcOGqAbj9D
8VSsP1ykO6HDocGXvIZA280cYT8KBZhLyybpFd+2Na2Y0oST2w14KbcpoMBR+XBY3zrlv9cBtQNR
9GUW/rOAdfPRy5xUVX2dzWH5TuTuxHPqBvsXDmdekilA5rTBnyIr4WST2M+m1zdKDheU2u8mALB8
mCOzugYv9WsuKrTC7GuD+jTN7e0GzQx+2u6tm6FkS1ggXfAAiTpYQCJeDTg97qFV1ko20Ed5rjd+
KRMmLryReA2Dbhnq79LPA/fRvt1wQFulTbt389W/rma0gX+jX0fU5k6Oqqd5mOzMeNV342zcnjhi
2b6SdvywSv17gwkljZORbMnnjbCZzuxp8q6RpApcXnV2+grDnUiq3kwOfPMi4VTRq36Suq/K/hGT
FusSc1N1/e3Q4sSihgcoMrC2AKq5LJc79sfzCCnqEbh6SITi2ecNbn1PRfdHF0fLrgG4CCfutRGP
KRTEYypZj8PD+Lbb+fxC20vRTSoLWFOUJ4xU2Kty1RxeIz5suhS9zCIzLjYN2hTbaCR7iprHvhpM
7hGrW+wvl2KHFlWa+/ywXxSoaWv9MXW3jclSGniR736DzBjS+wQXt8Fv0/u6NQYI51sREBYpNDOE
DhtuOiJSRTr5TqgnfTqwDfJPQPVZRTIb6Dqjw5Enyi3u9cnVXWMD2QU+ElW+grYLQqsi2LNbVgKg
ATjOynUgPCKWSLExktJBvJNzuyklvzMHSR3rAfO+JL/4qLaRR9zd1KagSCFJx12cmym84BTgLB9g
vvXlMKbmxD2JFO62bRsOMreAapuw+4CAhYXL0bSR5accpvuppOUwpmbDddfo3NqFbD+Vjggk9ZgX
KxPKvCPtM1M/pnccKJFH7m3SXXSrXD71SNzxh1BvTxHDgfC0xgVSYe/gmpQuW+E+i1ZDeVdrC7fl
adleRf6OUEWXgPX07QZZtLUoI5fssKgf2vIn+2AkeZ/yhl8Y/lWEtDDjG+UwEO5d/eQXroU1V/NG
ROl3H30KUUXs/mjNN3l9zWKNq3ftZm/BcNis9dPqAhQ2TzkyV9ASCRZR/wlkat7BZwyzixNMXsug
ruqxeeSF5TkLEG8/zPvftT7u821txH0aa2T+KzGcgm90nY972zPEH3STHWfBJjlhKJ1XhYJjKsXs
wAQi6mM+qCIR4fenecXD3/neWZGpfX2MlTB6ksrnDU9vFp4nS4s9oTB8lL3RftLltrL9/iMkN6ap
rcqE+tAz4iRi2bga1Tcmf+vTeON8MHG2tZcsGs+EoF0JwhT8/gmF8c3+5CkZYYodqilClAxByivr
E+6s8SabVkPw0xfB7YbVS1aYRqRm5QRW1/q1R4xAQxrJzBE1fUhC19r8pIomIEMW3gG5YfvIWc7F
3Dr8RGZlF8GXDQ7cjLyf1Rh9s//GgR8SHifjH5KiK2b2o+OsEyvMpnwzP2LRsY0w36/gIlULejb3
dNaFne8M9NX2OdFF1nDAH3vcbEMaD31mq8s1TugAhryfffsntdm+A4YIc3cFWhEhB+WYefgQuzlo
bQohNOo4K+ni0uMHW+zoQGGPu935E/bwZ6wdYNqfHXUTj87MQRmRm0YqX9GUy7ECJI5PCUfs8XC/
cWjzIVvp0gycuxl1qQtFkSUyJLmZdvhd8MCl4/gx9UsHdfB3u0uI7ciMyL2hlaJl2WvRMhYlOshW
BGJqnb4MhLZG3B52CfG8G875IynkkJZt56ZzbmNfkHiTMUKavITCXI9HpNwPxdwgRwCxqfI5yvs6
hCcZ/SERlBNBo3+fkLmZXgHvnW6ntBZZSzx9M3hPXgKVatf4YhGGPJEj6I/nIkE0f4l/eC41MSE4
xEB5gfHlQXqesa13I2C8Rlxhm7/Ey7dQyZgW2ZyIXl3odfawfcarmfarvyTy+hgM29SSE9OVYGv7
RVv4UwD2xfR1/Bo3QFSvYxvkRgp+x2jDCxRUaAcup5MTOzG0bn946hJjvQkowqutxgfIrvaHOa6j
gER4ybO3VN27yc8PlWi0IowdoaYskICxlEt4zXnw6fWEgn63U/4LhgHo/r5U263FafvEshpe3+tJ
fSZ2kg4eTDMKYZpJ5/123UINYH//CvrdX1Py/TVKWvcGwaw/rSZ+gzfu+c5v6eZR3BfBpcincTFe
uhs9bvqgy2AfFLupZRre/mvkPJpnL1fCNdQGPRzz4XC+DDFgjZf+CWfwNnflPqVoJX60E1WNTfsP
kYfpyp+foWycfet2/hM636savQfDarBbE6g0EDgmKt1+LEFSC2HqMmigFOGB9ZRDfX8vqQ5LX86j
/dptEdrmjj8fuL1WBkfqS4y9x6QVtWFzwDPnLbaPa3fe8rpsnxMBjoaxzJVXbRp0zFq3/ySvOVeg
n1/SKyhXADSsntkt2tp3x2cmQwfP6A39i6RgElSiZAT9IUaPNqevzB3uB1+KHk/Oem/w4q/inqDC
4Ink/X6/CfL3Nziv6FRIbeQkgvs2TB12rmMnK4l6exIBlJhpQvUnF98V0SjZoUI2WwObysvOl0za
oEFz6BocAh4+eQtutOsOKti0tixVZMg6DfG2OyQmO141svdlWCpCJZsqtpNOjXWSQ59UUXOflFpA
JLWJfSwGK36nCaYDI49hUcuOXWgI1rUFHEQ3fdAr2HKYvL0NPnCf+yxIe4rPTsvfZ7HPgNJwx2c/
KPL0KAj9v8HZZup2T3xnlI9xcAFjcV+cJApc/7Ks8QbJoGeDCsHeq8GBVypZffEZ8BKw1+hj2tYv
QW/QvgXFMexP2ML0u7lbeLu7Y4jEFvrvjfjNjJM4MNl4foVM6M4pDgFDn1sQ1Da9baZjXp/XHr7t
2jWPBht2CTj/4DI9bckj2WiU4DYOnI3cEOCkh5I06fKD3a+dsfa6yzn8K4M/VofCAr03tn1LEhI8
cXY9w24Jf7pNuWWErmvVwviJdsTQ8cRK7y3bmbbCxwR9cfI8TeO8HzhYI1vUyLfUelFE2NlTI7DR
JSUnPwIXE5ZXeCyc/1u7wiV7Yth+uVOHe6YqRapKQIzadsqtRa0rGR2wpRsuXI/nVLL3OD8yi0Tg
PjAB5+tChUQIm2wDE+It7Hjj6FbMuo4C2ZCtLBMkigRyLfLWA2dS9tKshMSizUGd8RS4KeSUsv8z
i8kLuMbpz43+lCdlLhztoxEVRXICFktCtyB4xhKPSI/9JA5sqMi6w1XKjCG3ONIavDYEMJVxyT5w
2WCf5LrfKmVhA48uweY8Ga91axH82pizOXqssBYglDLpmtGAQ/7IH5EP9VJ/F7ES/FWZ/jm9WWB2
re79p8DCzVjaHO7brkmh9DwhXnN1rELWQ2IVL0FObnFvOMCMZxWKnO9UZmKVVbV367iP2YmMyFLg
yVmIX73cb/dJ/fRaGjlVq4pWX7obVGYHceJaYUOMclD0ewZrKzW3Dqce7x5T6NfY72BjJrRyUMn7
U1+RzmYoinw/r6dz+lcpxgLYpMmMkKggP5coOlrCfd+87kzxO9LkSBymyMHOJ5EAmB4YiuSiW3mT
JouRWkK5Hu3LNI4hJ5AvnawO+WUPZ+8ac0tGUGtnL0txU+QSMIDN/Yh4RUsUZekxmCOyjherNvOy
IYdFWB8IB3CV1vArZjTWIUE2afDZfb5Kai+kfs8NYrS4uRPeTGujiCWGIXr5Y3hOeOPyv4VC7BUM
vvoxVIeWysEymzFity5hwUNJRuLB2tKVNwlLvsaeqalIzj0gUdRvEno5rsk7BD8dUFeiqqZc9deW
5y51oQVhRek9KEnqIaDFWJfi1YiqJtsDR1iJFrLXxOE30WlApnLxGQaciMWmTPgU9PP7SQL0xdJ5
DgF9+zOQx4jc4w1c4snkVA0LntIqmXDKdZZrpHFcF0KKm23UUR7OiDwgjGjEPjpUtOwOAetUzoXn
gG2WhzgjHczZM5aEqLCnZ68V4bY8bGi94Kj9Ek4zIF1s6LKrkgBCe64QHToqOYIjP94DdmGu6Njr
aQMYUrw/wWE/0uM0Z/Ly5vi1cjtw1vW4SyViIiNLijCOEQdQgfgRbP0oTs6LUhbIJ51mnG2Jk4/Q
1oUuRDghxUyakzUq/eK7554HQPPP0CRbBZWKiUHJzND1UrMmLHMKkqXcp0PinvUnTSTRS/jTIVmc
RgmQFMOENCz8qm3OqFta3ROkUZymkyGpy39IsODPCIDStvYi3oS2LEeyMIaGEDqIFLQGaiKWRM1J
zQzsMXhDhBa5TxcHeDrWOVL3XposGWNyH3chsaD1UR/nGoZPA+/9u2s/cfYIZzmQMRcB4W6E+q11
h5SsfZ7LsMPMh9q2uYvaCKFfx+Y1q/ACS2yCaYYNaNJLYZ7vamTvYgjEuHMpptZ656APzMBub3xW
J0GaW7gQdygD3XmiINzpyYyRPhdm9Y0p2dqXHas935P4T0BK1n8XRF8TKMzwbY8/TRUH/U17424M
c1VfyYfIEk6/YOvqlM0r1JkQyzluV8005fJayXgQRsftCcU2+LINFT2sGGPXfFWGIN9jbbyCBZ+/
Aafy+EckVdwNC0oLmcvXQIjgi8cdvX1LST5G18A+TSl7j2e5tdkgz+iDV0BNlVrwjSp6udlE/FHY
HrjIt6G+Kmu6XWb+26bO2rGmmtMGLQ8ik4O+YliEMRywh04veICUgU04YNY5HlNdJQTvBr8NL1+S
YLW9Gif2MACxIjkmoYvFuOXvDIaersvrm7E2CSbF5Ahi1qWAagkbMq62uyHq1ZSlEqpi/ssJjBvx
GDdY9ZbbsSyepsyrVKL9up90/UaWxN+ix+1A102kSk47NijIi9gW9LC0zrDQ947LEh1bLpBZ0bUh
p9umpvRkOAYx8zMDq10ALk+9c/OaUQ/4jblgFcTHUW7+ox3CJxQ1Sgw9hdlxSawckKr0My3geL1E
6bNIpO7F5ODAV0cQ4YgB3Ax/yQaGi/LA/oQ5EMbrOIX6zk/11wgVk/pVwNVOJ4vrC9Ysf2P8WRn1
Dmb0+Iv0HVlZXwM482D502CnUFbGc2WmJimxYKgNMZQgqb8UIW1UODLfXyV5piCvyk4WHPrPZapn
uSixJbr+dSRhKSHttpTLWABAGzN+yutUozv/LIy+8gCz4dWqmZ5vKr/B9oUGKWxe/TAx3RXrDR8z
yNDGvmG9ZNF/JYsC8b5dsNydbJxB5Aj7d8SVLha/Y/SfdzHhMPKdLamJO8/4+fk58EfgHJvV9wgN
5gWOIaEcpe09V3jSg8GIrUjvhAxJe6Fk/u+z6DscuISxy4Ruiz/aGRca/mM4l6BP2Sb4bTTjqQCb
1KWKtXCdAdn7VzLChv/wqZqnzGRNGdcq/kL0P5c3VnoYSvgxLgUmDwr6umML9zEnQUeWNCio3uU/
4kTDHAAnAHIDCP8A85O1/WMlx5eKk9NV7syp/MqyE9lyyoUd35fKmB/05KYbFnPKpZVv6MtJ9CNs
eHmpiioLkMZ/ahE3fS8wo5LKBBpy/FayZFfBbte31g33III8b2HMoFUWmFg5lygQpn9SHGFr+MUM
+JeLFXwpFgUS6hCkieQazHvnvbQTT1G6BKpfUr3DvYR0MDJ8Sg9z2bJ6lkvUFPw1Zv1U/2jO1fl1
vBAoz4oAdqAbJCXSM/9HLq5KISzBBzeFcDw6Od7pYlLHNdShwfVsYCg/rPnYdR46/hdWHhk7cSjM
oz84CnrltVpHBkIErRfDkf2OK5AlRg0RO633KQJQCrpVZxqDsSFv/8JY/m23k0fyxCrJwTSh4Jy1
Q9iKcm8rC5jlLOcMzDakz5Cdkjifp3S7tuil53Dh0MAFF6FuX4SSPJu8Sglil1WMfhTL4qSRZu1A
YRKhH0Ws9wcnOUIP/pbDBuozwi4D7lKNbgFEzpFjdsjGB09MuIbmGrO0n3B0jVKYNV87uhjL1tk5
00nkVT8N75+uLCMPlvp7e5m4EOeBbkkPNmb9pkQC2A7EZlWXG2bavZ9hs0IEtglkDI3RcFpPJXF3
C/pEUH/z+zwxu+WhLwak0EDKuahWWNY8xCrAEWc/woRD0bzTnhP8/1o0sF+ktGUP6yJ3dfILFuaW
k9BLOBzkdpbFitIVXxLddwXPLU2LuMeb9k+9LE5u5/qinGJxquiKlWZeaxBqC/kBB5XgtwoxCEYd
9MXAk4V/xt9UtE4MXHLqI/wEj/wBmon42928M//ZD0k0sqrQ8uvG87bnNDp5rWhT9DtOk6DuE7pL
cjxj5RzP+TS2XE0SsiSAMHskO1rui6Hrw7hbrV41GzQyBeS5qMVUmks14289s9sotfRzQdbuXowW
cNe6KH2y+n/u4AkRwIjRNTUi3lNsvhZyOXjUQiYLfsCjaKI2Iw7AzieaxiEIgUPtd4PNLhPGhgCY
41GSUg4lQNoBblRfzaWa0C24k86rRXDzv/wL44dpWSiJELJRriR/Gp7jhbi/NxUzjaq0NaGt1DJx
68VOed2VnuiMJRqNO6MFGKM/zz7xP4O/gemAgeY7vGixk9q75Y8JF7SfS1ZxFpMQQq4gkd7Fvi5K
xwupeMvSYumbrecVzIKRQZltJJB+TXNHIF5rE0ftpI/qCXTlQlOPufj8bQUleHJaMtOb2j87XiWg
ICwBldUAqmmMv3rHjPJgjKZwdsYr3Eh/Phx1nQdb3HSXrZpltaIzZljdf1d1Htb8+VvM08ZKlgXv
VYTbSwJrWLExS0VY8qR/unn4uDrgBTnBECPDH8PhazgClSqckLCP8CdmSkouiJdQGtQcXpPVvcJS
aVWIJCuYMZ87vPOLCvxJy3jePStRoUhtEqvPQXiMjdv2JIeP0q9WTtkrc6+c2l4GL5cXgUHvfgPA
Q3/Cd4RvwCpGlmllHs4HTmyiairU/ZM0rtRmgIe2L1cOcjrusyd6EJpv37M+uQhggnc73GXNDkXf
qZLWV541Ua9nWxqVMOCvTLV0XqRlGwMG0LFEpDzf7bL+cFJocOqZv7PKm70pfEbfXohs9Bdlya23
rG710sHzCrJ1a1ITJvzoDMxWckSUEqhA45ahRQZRnjwNHwCTV8ZjNXp3oPu4Ho4ZdwJVhc8nJ3E/
7xKakDezaMwyY2rzKghjfG7+xqUhT7ScjCCr1TFO4sH5wXAC8kNxfUeZ1z8srUY5NzAXpR5NFIHX
a9kjGmCTwJqD91+i/2BgJ3zTNm94LBVY9rT2y2fo7FbpYooFYUil7wO3Q/AB6RbFF95qm33NB0rr
tKyH04aMSm8cwNWl0E6VgvdKm36+pIAUU1zrDhhWX5rOnIyht0+ktcINVa0X9/peJx9M/CG+l1Bm
cP9CzImbP2jyLo0ezAvWYeB9MGBDFBPGHypttND6cZBT7NMNcB4e5cqTey4Bfo6uMS/Pm+AgjKz1
MZpLmeV8XWdvKBjYHcPvGdY90cOCGNWiGxiHUH/PWZ9ISICoPTkxqjS1kReyL2C9R2ayMV7aA5Vi
KtQDHQRF9dvKUokKvds3pKWZLKnDD3+BCfDHTc6JyXXcdS6n9zWAiSQQAZ6EcEHSDMgVmFM/exXi
Mqcc9YO94YmbLSAvMda0JwJ5JluDcqHiOA+11FKbDb1QnleJUx8a2qD/fOkpttMfXLo11J7aVPez
jkuoQHU73UKitaEC95l6pdSqKBvhGu3I/RUzfIZR0/PW2RNOtZwV7jxyF0eBcr+lUIFX79C9jQkG
nhZ7+U6QbebQ84baSPEKAUDOyK7KZadeQ3eZEGcUowivrGQsAyPtCVDJlnqwDLoNnkpo5bezzUQ8
LLtGH9QuSaGNwkcoWlmhag7l2o+x9R3/f2LKvJeiggCQZ25jkqzXiorndGyq8jHE5hq9kD/JmN7M
PgTcNTyPHAEor1vecHhw/uxYPGwkvQpA22QdM+j9oSMh2MR02GblOJXShT7Hxz7zPvxYP/g6AiOn
KpJAoqJtGsWpWvHe8WfXeHUabKm1Qe6z5Ls8ncW3qxFAvOMOCSLc1L6IeXger7M65PGEjfUR54xq
9gWhQKpA1KklqDAyCLwgJ5Jz1O2/iUROeJ1Wt+yZ+voOIGbjhGA7qmAKRfNWNDUY65uifvorbLVy
6UaeEaCoFPrWkgUntT5w7Mq3xregDlelo3it5JvZVEvEnjbWqCenOLzfdhUU8FI7w1g6uCTezSC3
M8xUeKNAXMNIuEpxfyOyvMJuCON9B+MGZJV34iBh3HEltMt9wNnvTzSGLuZAA4xb45Qx3MvcWnG6
+gZzBaE6E2K4cexMyOQY7HvJ7PZmUgrSlkUB1BQStR8Y7LkrANvPUA17ybxV+zIXczyBtZ9kFarv
R8dG7xzWMm2iRz//QiG9s+m9HBORHTGRLDagEFyL1aq31ajtCWuKkoaQLGh1wVkUmm6fgYvXyAvt
9tWHYmvDtOBvrt4ZJGyrAm77Gz4HDA0lhqL4gesLcF3X8ddfVK63oX/Pzy6sv5+zIgVXJkNu4Kxa
c0I9zkFu3NNG3fhyTBmJwJ/hZXyXVZ6HyZFnB2DZhynzz4DJthieMG52Q1fQV2OpEnjqhwn70ve9
3G5FRTQ9JnjEEBW7Pd/A4Z1cmJ8YfkQ+cZ0EQfNd4ATUWpaXWz5VlfgeI7oIOn1SwosSIw+xjOBv
Y7vt4crIbvqHJYaL9OkoukcJtj7IfgdT/sFQJWSIs+woLHokwx0/pCTSMQ2dfdc3kAKSEk7VuhgD
tw7FVgMswD+N8KpWrn09boyUc/qAJlUJCiy5a8CZLVgSRVWqdyXMwvrcMRSUu26vKDYM3uGLafyj
3tvBHLJ2n1oRH9OkRhFyYpdNK1RVM1pZZ3dWIE6i2hUX6qY2TYAp30fZT6XMc8z+MfPIWOo6Xl43
Yg6rkQ2v+Z0j+hs0JdG9XRODpXUUO8XVVJ8eXjRFXK4FQj9y4gcvgDV+AgXpnNseiBR7UcHOF/TG
4hSs027kj9s2ujiwQQ6ppW5rN/fHPGJc/AU7Jzl3aCkik1/wF3R43UZiDq5ODQ+ZVL3jy6WHhbgM
cJNbd6NEFYB1bX/PTvziGz8+Cc0APRBWPGh59o24WQPb+ucSRR5HwDN2wQTkIywSxMLITTHMxzdg
kojcYRwR46BGY2C+lbU+ZimfbbtLimXLikfm7eD51xdCFEd1L5f+3l3X9hXaosLSLFjWuGvZSMJl
3jl1+rnh43r3gjzekL+ZpNXOgawX1/bm7NXczTr016tU+r8hjoQIMpkmWZwlqNYzmsDqcoVl9sUT
ZIWOkXXP4NXx+pS2KxWfDV86ZvF/TwftLpPWs4OUzZ2RWrDkqw9JM6xYmgC47LWvxFZkMu85CSgv
wQeDfGgCGbXJDQZZ8AGvNg7uF13WAiAp9vjVhYDVufQFmwfXh/xbbscUpdyY2e1QOYCheRtbrZ8d
xL8Lbw3FJaAUkOX4LeKq/c1Ra6AqWD7e6tIisGd6AfOzt5hZXsVAmBPafVX5cplzlIK6LSjinBXG
eV/eyT6nsag5ne+PcNyQCz4vl1IKFl2dYifmK4LVETHs3wdhmXDCw/QQmrBh6mqlrw2tIeotYgfT
vHHuPjWX7pa9yU4jPRbcEqzrcot/v4iDYifLokjdqzDav4nklqn3kvzKsjrZvW10e7Fot9pPV7Uw
SDOmQD92baCzhlhNla36Zx+uHRA4MRsXl8HxQLfgs24aKfU00ewa4TWHZoWwPFLsdKezKd1aqBNt
5S/ehOCHORQk66Cur4WvPoRl0+m96cVKqYH7xFKtoST44B9YTBsCZL+xw5Swlr/61jitPU1MeG75
viT41etgU8q2ZFqkplRUXcjvCy0xztV8cUvbM5yRaiXo87k67svIxsJCb0nbuL3ox2Iv3Dv3Kh/U
vKgs+K3RtjBvWkKFZ+uu+ZhiEeDydg6RmygECSxZmzRtB4WTv07XlIzUhEZ+ZdKcCNaHVzlTiDG2
/UvWwSoZDJOpa7V8ZrnBAE451qwsKM+ANOhkvRg579i7Pwq2pJGn7t51mLDJKhGQ1V11/EMc2AaB
c+D7yDYWStRNSUkplIAh7RzqyRnzgut2cuZaAxQC4QLK5eeKC634agSYgaIHeb/HKrWVrwXOpgGU
EnTvjjSLLgt6lQhtEQ+KqCb8duG5TSmruWNIrR6kbRrOC8vy+pE5Ly8GLAxHSiwyxCaPMq0D8w2O
ZXVAXrbbKosX30GWQ0ownfsjuOI92pmW7lFvnTfca7e6zC0rghJQhenEpfj6z33lqF28kzitXh3v
lHkSEyDEF3N4Qb/j+SfbLuEH6IoFpoHmF249QB3hS25CQjWJ+Gg2pfkB3KfqEFktQ7t0ND1aTk8s
00Ns/8ZPYJ8jKLm1MmULzjS11ZLtRCR1e5jaJvcEr/HcBhxD9t+0SEYXmcoGIrqM2kCx5q/trikR
/PfZdsCanQADWPy3b3yyhSrtfGwmEPoEHGoLTJ9QIV7zo3UFBD022GPWDTarI4uhYcSoSqGQDAgy
CL4l52z5fJt1jptuXxW2TE5BPBMLgf9UwM/VB9i5ZWtgRK8XK80BcXQkGRq0EKSrgeFJsI1btE0r
F6yDXODLEc/L+px1FDyvhTIWwQWEzFYQV3dDf9fy80DCP6bXPUDCn65PDGsM7uPIb/UVbTOdy4FR
ySnLkCKvEb6HZ8Z11bcHfTYml3vjZUtLM6hf/1fprRN4HCujsPHWLyM7of30WKO12ai0L1k8aN6Q
x6MxCHMUxQ6eg4JgvHbG9fZAOFlr37lN0Af5IohlU6vl9+wzSVdrfQShlgkrgLFG6GfQDEcPEkGL
6YyKuSLVt00PKdW+iQ+SutHHACjmZHg/sAqzB6zcNcDHYKieS8NzGb5hrBUZSXkDJh0iL+ixGQCk
GNc3kO2ZL7FJJ7KNJoIPbu8Az0quxi0JEqGz7tcobrslI45CCrPeLU3eSGYmimbXDOLahPo27AdH
+DerUyTe6Ug05DapOqsbnUza7wdP0byq62d4KcI/kxNt+PZi2VD4lVBp0Cz5sceO3B7ysp2CG8Q7
mUOvSelKqnjY6OAUWTkwSFwfFYe0SQRUhrFE8r9rQYgCKmdZqqA81tYWpBaftaBX5daEe68uN1aJ
qySrk+TzsFXHEW8SYwrSydozCvq95iscj1hhVN3/Feq7qEApKkbBItiwUV0Dx/oPFyvBnDpxWr4q
bXNHMN2sOINB+vkquDcchjSqDb2rfS8npxx1V401C7oPclwoazw/VfYfZObJuAk9nf3/vApIiGas
cBpEmDfXpduZCzipC0YPh8Bb4Z8+tf88g1n3PBulS5/VTdh19xrMIB9q1sjGNgKo71UUxRnXToOM
n8lXAjZtW3GLKSgGOsbeqLZkxHuUXqUr0+EdAlpXawTfkGkmo+e39+MBUs8xhyr06vbdYGU1QQ+h
jX13KfWPwH9tyAYY4wav2eIkHPP6G+493o5OEc28jw2tynaL94ytUcgmKAXqsHkix8A2P3JeCZcG
57Ik+W0UW7gWsguHgb+kGUk1TmqCj08AU5bGI0LkaVRuUPc2n2SGc7s/MwSBexoYdkfECdMTXzG8
KelYfJaVSuSOIN1A0Z1GskUw93o7eWZrRNaP8+lqYoH4GH+MMnsh/f+BxSb4ylJkQTqR32ymhZt9
GmGsm6JioUrJsifq+2sfDGDlrCIQO6lzaQaQ8YeSNGl3vuR1raICvGr7j36iaYJ09NIz+nJktb3w
DU151g/s7fp4eQ9JaCa3MNmWo8E1pvKjyMiLUq5uU48umyLaCGIwBWk53TwMiynx8E61L1OQTsIt
oa24Tq5dJT97xugKh2cvtMupVVx7q7aVXzehBaFInF69Mdti2Otf6GjsIBAY9NieqjGQeNbLMYab
FDhfU0aqFl9WsDRNtdFQAYcYOCxGILVsAxl886If5fiogzBJ5NALinBr2fzNZGICG6+2tQxq4qPi
2ESnq0Y/BbL7AGNKzonpNZFZalH/KKCpltcMpqI4o2cduab/jzrIH4HP81trOmNnhuj+eH6X/3za
xiwTln//vlahWkK+wMUn7tQCF71xN1i1cu2maVihkLVWLhH5RKtI2PZQVQtikZ22XE1qzbSJbDpO
PSoBnLPNV2gbgGjhh28yZv83sAd8tFZ/kbiekLBX0ySUIYzFl4k975wICGExmw0PqzjZne5xiPIV
7nRvNTJEcwEJbPf6/QMIQThBJze751UUuA7pIJyH5AUaqb3KkQKuwAvoxwDxZzjhbx7XCC7CfqrU
pKxQl2+YdXc7Hrcsc80OVKXcl86J06VGnZMR7rvoYM3i8n4+FhaQ6ADcnXyVX9tvWwXvNEbFkf2Y
bGXaECiXrDnNQOcJwL0uHXUPUjpRyrAaICGy8ayHbyjMTaqYUAWM0Sz7X23/lolh0qT71HWcChQy
WgRzjsZ5hOKVrlg67aKSHENDF8V5tAeYWnIDi4+Q2+OpE3Jeu4tJymiQLid/ao6YHBk611qi+jpt
Ryo7i+e+3W8EUh1jgg67IyIKrocPlCtNvJbN5qeKeE0KkHMpPuGmLL5ww2HNF/IKV+8Gw/2NLFFX
rlTDQiLlOM7MsMpmHQVPg8b+hsOfckT/LCIuKmrYif1i3GPBiC5VHref+0iUpSoPAFFXdJ8JYd65
wRF8/AIOyT9LVKM0ObxSQmR2eRajWJodkD+nTKLPJEF2z2W65Pp936TDpuYlRuvg+D5gY2jCc8os
22YdI9zc2NVMxmtBTjhzQSUcOS1reSgXwFizMfcv9bJdAWtGK+vvtm5CdccroAskYPdBaQBhq9CN
1oHmNeF6GYggoTZvRNcPcGVRw2+WJQhqFrcJh/qMF1PH3kruap1j1U5EKAl2/qZCWGAKds+u+5EZ
pfvhF1ByHsrtDj9mkNEWjZzXw4s/xsOA9NHr2srB1ongm8pI78WzoVbb349vSvtZtgpSu3ZFZPf8
kfsaxXxsMw5Zz5HmjO2F21X+mK2WUDNAiW/AvaNMEUx56/rGYsfn8kithcqgOYpKwgL3BljPJsaL
c0UbqHnogRueJtf7pX1ea1iqpuVJhrYxQX+QKyDJbksdKftYlCTXSiJO/cKxFL4PhgyJ5AF6U3vo
xN6IOVkAaRLRWUkqewGzhg7HCjN9nnAwMkWgt8O2i2aAUXw7WiZAb8GRvn8l/obXZiCkpPViDDI5
OpotPN5ZPvScpZGY0E4ZpAMVjrwhWhx/MHI/nb5Xs0c/pEXsEEnyJ2NjjzpdiqGMtdaiVNbOTKay
R/gpo8M+iN2AYfYpJ9riFrUUzj3xpagUBVJYRBRIeuV3f1D58CuA6ttc8IoRGBHz4KvI79s+o9K3
zxcnkFk8IR1+a38mJ7s99HKhw69NHOsYORzPTFqgSAUHN69/Ioe+f0poQwLB6FXRm6vF1YdkigAP
XntomVYf+q+7PCdmvnTRLPc9VKqvQdiYtiKmCGkP79l/H+mVwka3cxsyadDf0Pbk5TwlI9W/dTpX
bT8P3oXAmHVpM/78yeUoRc3bt5tJLGmHt6LXZMeZdXhxXv2yyLSY9cqh/LIFvUH+wBmcNjxLz8k7
sQXFbuGRKgDhUl5v2JpjZOeLOw8bG1r8zSd+xEdbC+Y7/w2a4UO6ErRM4qzIP0OhJvACrqxP/N7U
2vcdRiau8VAoGJe0wAjuvSGdwZFbaSoe9PdodzGCOlts8SEsMr6zVCj9SLBx/HBuiyZdrBOFjcRB
gAMw0q2o+NKGhXVGIHbvl7JotAjiHdIULj4mtIeIUQBYyKbUyyGRr4Mt4mSwS133FgTTjXASFaNr
2h2JSuILlcr1csastaj4mEcShZyy9GOpj755N1hzZvM6uLuI6RzUveKzD/4J3ULe4escO1eihy85
uogDU2HArrK9QT2Mld+9F2DsPso7VPOaBDaUXX8nc2mXN13qnYVKn9cSUkxvTn0pEupe97uUSMyn
mUNSqSGGC+Sc38RNnM1LhrlO7zz1Yb5aVeDiz1TtSSElgDw5HeKzg95QBGWMYyw7LkyeV34tU4oe
OakhXuv5ae47FWhgHMeZE3TKtQeAlb+xycgyxdZAx5yLAyCHXqMCbzFe0NcJYgQ9q6p6i5sXRvLq
ipXP4EOqe+tQdiEiEMVWXBwJwKS9+qqT3Yh37GdK0hLk6ZRf6WVeoGPO9DCzMXbywf5YP02/Y4XX
bMnTCdz5BhPlC03lpy76vaJ/1lhjqcjN0TxTqIiICaztAwQ0u3UGtgI2Ear0IKbYYONI8QQk0Ens
kT1pW+261FK3iQ84/wIdnJlbxCyRXh0xGNeP5w2xCekhATv6mfplWEBrM1pdD4gGsx1T2ZbnRph3
ieFGEKZtbuZK4Z82OJvM/uc0rcR9fzjlQrp4po2RPxd8sQFFJwPOOGPEZtZx3reQrSctLuaXGQ6p
GKyPoPefG3lIjwlGtNaruB6JjkdHEoSeS3wa66AOpJx+uKFFNQ9OTqokbXwcEGQID0r7sZO20EBE
faG/RM0rb/2N30JoP6sJPZUGqdfIh7JmZOfEqZLLeMKEVzReZ7N1w9W0HbzilkATcpeoPdl+HxYz
Qj9GPJ+iwlBVyRXzb5iBpyEHdRYVjCCucQBPf0TyYH1KIG2NzzYqn6MHdrxXsvVbcGGhC/Ac8hzg
RcuWj0EjAAi+jM44QN5D9ApgdFU2RwuALixIjdYt3dd9JY1HuK+q5JlSsvouwZqbp/Cq8NQny5QN
Dtm4WVASLsGV5j65c3pPab6V/cUd0jpk2JXKm8hgMRp+7qh6lG6bmStiWFc0iX8WlfeTqRZJSfBL
FiHfM8kFnIv9YYfwIbCdovHz39n4OU6c1PyyqvUGXHubQ6SD6ju8xlqXjCG3JDzUDPwWqc81vXHP
O3IbbT3zLFCwTkYINJaTC19zU8B43reDWhh6u7xDbkACDKr/zDK1USlNOgEphJ5bkNMW2ZaydsV8
xcFTzUYg3d1RszH+BeNkQzpmfT00dRlQM/ISWxgm1Z5l6fm/mwKJGhZqg96ilo1opgpQFYOsmKC+
8TzfOD1QtE1Iye3ISguzTUyz7v7MIinLtnGXp7ivN/vGox4PNr261nRCZtGpRh1MwTwBEX2r4QGK
I2WqwqyWO/kDTlPuFZMWBTRn6QLHjt/AZe/AWNNVxN4D3AedPzVcJRqTWnxL6T18XHTKdBPNzBKD
7eaPT4yh0cwIGzDkyIrdlY3mYCeTp+PAuEFXcfyX92KDW0Yma21r6g+hU8tUw+Y+wHk5nbZVhpC9
sujiiADCEMop+zT1jr6+3Nnob6k7bfuspBqSL0q2qVlnynmmebYgLFGBovIxgl/63cQZh5VSDWVw
0HOy4irIHltrdiWpCV8TQomVbUKxI+adzXYTWLRQyRb07RhOR6lVSDKICKtsWRSElBwL/jQE6jW1
elPUTHk9d/SHlyzIyWEOxbtQb6MJTWf43tgAh5rd0lDEBggPS+5kZqD7WgCgopxU8xncn3ImU6O2
w3T/TYwPJc+KSvQOPjJQdC5AslrV6hpP81z4v1HyUpyXeqr4uZrbfBfumVMXeCzcq0JaNwajyRsp
ZmpPm7QKQ25yoKSfRdjbjsA/QKvjj2hStqbUXrHy8oFefoAvJdHlRXneDeLsrQ45fkU4mQfEJMSx
eeAfZHrg8unFWRoxD9O3/Y1MZZWeKluKW/Bx1jKC+phAogppyA/78cFCrIAX6PoZ9TfZHnPRN4ts
WMzdQ2tu8J6JgKBvwDtbz/pPBTiZGRDhNMFc3i20o86jtRbXFfRDe8qQK+zlPbRocnu+IDFlhex8
KrPbbM6Ju07sI9umwuKHpdXGS+Eeah/ggyoqapNvivwJmzMDbuL8ycvR8mA0mEWCMCofF6yPKNjG
RiksAo5yGv0VQl+h0UlC6c3qKRmXF19ormtG63xLuhuHn7Rnisioqrvqj9Fr4Ks09tP1Qt4UKmue
P+umPbZbzb+VMHmfg0McgQXEKyFn4VpLcjIqOya0kZUU1kQYcTp8X/Tgp05IU2rmXTZJ5e8bEifZ
RK7rmursx8tGxapUbObydPLDF+5xxAYIYfocaHqz11Y6nT9u0vqj3db28UL9sC1q/Ng3uffJa78N
OfVHN3rPchGeMg//5eL+IH9ntB26Yaiz1qNmwKgx3AD5iQdn2PdWriLDy1UroTmkehMwMt730Rwj
en/YPw8sbRlCBc6g51giJKTXf774KcBZcsWxA2NvMwLjaWlyG/5L0jzWzV1LVIuGfV/elfiT+xU0
uY4CmnHtza+Lapz2aRf7BRf9b1n9T9c+QM6GFUoN5EDq6IZotb3q1oU8JjLHJqYcBk9WhT710tO3
1E0ujurDQrW5SBJEmgwoyk7hAVh1QXc5uBgz6JtJWk/pDkAA/Bq+QfbDEBVuu1c10kBMwt/EZaR0
+aKuYtHb70AqIySUoWYoQ7er+7TC17PTTFMxM/CKzl94N1HqTcdwYuI/rX4SgGw11ilXb/3m3Fze
H8dPWiZrQoZoQFG5T7sBJAPmHjl8hvqqLSLrRKHbgnKiQ/rY0CbgH8lPLvMXmX6sOLeZBC65A/I9
GJTwi9Dg4ihGpKYuYMuLJDCSsuUp+lzczMraIfQ6ueWTTrL6UbK7tJ+XQwCMI1KJUrscWNRre5Yd
6N+xioOPUtMNoRH09ZoxKRTcz0Ekj3kgrAFjBn8q5vyF0F1pocAKjMM/sbfNrIzOfOkR6zaukeXW
9JTvPj21UzupKYsPLP8XOJrK0mvrJkVR5116Nvi0XpLmmyossXtOhs9T0627/5ekEYEc7SlQXsAW
Ylo7J09m8kk6sm01yYVjSFGHht/y1ENO8gjzdvJB33kvTE8iIcMEytVmRvBD3zltqdFAkONmUoUO
AzZR0APnivvdf5sm4vdjqycQgcY+wJRHhI65MQSsSo8iBrIYuucEChI0FPrGxmPlT1/52b7Pk1cN
UWrlgRuBGccYRtKUhHMBya2SCNNokdLw6mFg9xIZnnJDTl00iJxpsyO8lOAg/0BFS7s2TUHImJUe
CRTe9VLOZeT26rrIj8U9bHVXbIWDgpaBDohtsBt9B1ljrHjkYjsQXnz7Q1ilCHk7QYS6QRk5ZQ5L
f+yxV2Z+G+LE13KrhAUw2hH6tHabqwi5VnO5f2JjrD4Vt81GFSRHkKzZpZOCBv4SgkwtknaHOYYB
9FZAptq4Q5O+3bfwTkxLpow5YX8REFY5JPK0A7PD0cQ4way86JsnJ+1jNKqvNwvCmjkAaWdqs71d
gL0O4OSVaLYgd4pP9F6RBQmeLenKombX4/FQ7FpRr2A80PL5oJnEnNb4LyMoQ3PloLxdGbMHkqi8
FxbfXnbcoApx0jA2QjVvpsaRjyUx/GwEJcyZ0E/Q+4LbOqLzrqmfOVe+nj7KgDmYUgTfBRPAVbUr
k7tuUSWFGz7x1YOpDsI0FC3lup72pwTtVQWA+wm7MDVUx4lsH6AqNT3ICCZm0TVdJ+128dIxX1vY
Myq1sk3+AmjGaWvcBeGRkqP1KK5rcrNt4tSmI/6K5Kx4m8nEc3hguQNkYGshC2kge0cZwjIe21DF
do4BJM5zazufSDYD13QXRu0CXZyHwFG40yYVczFlkqbb8v5k+IOYuaZ6A0szSswmYLX0j761nlG1
Bq8Pl0TV2f2juHaMhEAYGX6L32zsK2kYHjReR4eUosnhaBuhsBg8BJdrVOH3KwaFyBIao5FFFMnh
6nZkuS6zV7zm06zTozI15g+Ju5MpRu0mi6oPW7+7sX9esPS2ji5+yHujybEyji4xA3sJVCqSzpKD
at+PyJPk9x2CvqciDsE0lQZzIzRR/20i2KwRs4w7L3sQAlGnN5MtU4eELkywR/G10rtyyC5OYt11
xFS4Prs0YQVyrrf6zM2QDTjbt7a1EpU+F/hFAUVPw72sXTNlPU1ayxUzkYENma/4UDJbwsZQIt8Y
C3AunmbYe9WQfHngVEAw6w9hQ27vsZckFcO7Nh67iK86r2uTA0aQOBTBycSm+TI1W/qbgcq/CC1H
ztkLokR10eaOU3O3LwtdREEoTq/EAZTwIx5NzG+fcCjt25y06G30lVphZN2bWC87nukxg9+Ua3DC
o95VBtdulxY6Om5WumZLUKs01uMQtDpAFbo6PAIC+jCknFNHBZWDakeLGEjYG7n/g1CZhkAkX3M/
5FygpG8o3JyM2nsDtowehVQ33wl/jJTZTnZWWcutsHL3u+JYDL2gZu3iuA4pBc2Y8yMseEogvclS
bKPvPMBUwqyvV7T3FcQMI1tx+wCWmdeJBbppQZkfU7kL70xmdq6W52ELfuyZ+qwLSsedbpqMusq/
M/tuVojIKsvMvRlctwYRqD5m5UOul7p3sg7w9CgGAMYPKCulv02m185krAd4WYyO2eBEkdan6Rw4
03HWOjbBUWjW8GA+sLnIVudCcMR6iv5xE19J7Zv7gPeCmCpjSOWwUOwepCHTtdjWkF8YFvhar5xz
mvutthI6K0mf+rSjkqBEL0nbJ22RekKlnKcVoLR+Vb2P9VvHzDFC6fdepB0YyrWyDRrsmmSF1iE8
8qCMYLrQgAY0lP58Delzrr4BCOKit5jSRgXdo9LE5u0812Ai/hIH42zFasSwMH1XTuyNWuL55Mg7
6Zqzo4KFn3MO6g24Bs6nIrRf6AE8x6+RpBgFOCIK25NY4i2m6uVH3vYAU69k/XJMl6ej7kkY6hiH
wphwR2ro1y8skbjffJSK0+KGMnM5QcctsLLmYwsl8SY7eNmujIJRjLP9uSDrWY0/IC8VwY+Gc+It
q/4xwUPTKbv+qtwfToO/3+1NcWmhmMe0U81p03n4YqxWpfKnYREB+EBDcq58+5kXgfB89dSSQxfN
XxR8tiJ8rMYM/HaUcKy9y46zgufqkKwdsYtsALXa2adZkEF/DEcdBYhI4ttEc7bE6QaJF3DtWwXp
sGmmq0d1zLHEfMvE6mWu0sZ6y/7xyY257bKPrCEmzyjtmXkjzDuh1Vtf/WsLy1hc9nbIF9Q3Lrva
miaLg4S1LQpPbu47xrrneE95dTM80q0LwAemLIvvWqMx2Is270e/9M6wIP7GnZcJLzENSiI1de/d
ev1nQW5T6axUD/4v+kD7PzHwxZ+KUpS91nReJnYAqBSQErrsAlfQ5f46Keb0mC11W36WzVXzkVcp
l2cVJQ8lgdeyM9IjPWPp7ofeSBWFfyDjL2ze5yGluzejScM1P4OufzMNFEOQEKprotdUHkUmleEw
jWLkzIpX03lHJvnOt2jY95ATNI8qq8WVq6uS4WBLlCgq48/lB05LfexrTS85WcxV1mztheNqMTcP
o1Ix/pHsjZcYC6pdg2lWPjE7MVUnSmMWI0V1X/uOS2cEdzEaZ0begvPI/iIN5osRcNTdnJ/ZtyWc
U7x0a8hns/8bz9deSv1quRjnE0aC08+aL+XzXdudiIlhuaF3IurldVij/O6lWdsgOtyMifV2pC78
4TVctI+hDZBhHjQLIUpjpmQVr2u0mD0XbXH0QL7b+ZEAXfOqPU4czQGnKBnLSLhTd8kcqxNY63mX
7I+7ylTERbl5y+IhAZAh8vi4tb4bKoeWj2gmRKxZzZIlq+47Km/PdRJUAtOraRPUVcLNNk6hWD3O
2Nxk0ghdL37mit9xSoFQWarY5CIHafKsEWENDV7k/rxPq4pvV+tQzdZBnqgohfGkh7qqha4euIiq
LxcjHeFSz6sATMEQupwtRZfY+KZTSUXu7fIZcmD6P/6U4BgW/MPba0BFKmhzObDN3ZhHLsWxm1FN
iUDaeIVyMZ3bCO2IQ6miLGrcbhRUHLgKpSH7UIdMkgwVoyyPPd3RkbJAhG3BLoSstCiU/Y+DG7fv
zoEscUOv9iiWDUSM/SopS/a5G2a/1S0Hol2iRTvebpGecobEqzOTjSM4OFevUICTr9Ro55YCkF36
dtdraHlSY9N3Cp+yQk2qakBGibpmgHBp8kQ6YNSXr69mjDtaJvvCDiH63pvJBEN0lxf4hcMLut7E
1VU2ZXG8hkj12OehOqGMuA3tB28uzEgH4D0b5xb7g4jguY7MeOblG1aSI/hJSIXxZKB9bi6W+Dqv
6ALAP2SXd2yeulW/71UGcsGdPYyz32H5PugFHQ6Oh/GjSUrkOWQSdeqimVRhvg26MygrNWEpICbq
/uEmyfDpx+dnVqxCwflNNEtRoxBXkANHbxNLdlLuT7iUH2XgNt4i93hJ1fDPqrkZ2p+s2IuNc1oY
UPvi2j/Tol44Ru5V8pf53d/cl46bGemxluBrFZFgdApep5ghVrEebENcViWUrdhywLB7UrQTeO17
7McXG06C/Tqxn1gh1b/GF+9EKz5ubT60nKCZGX1rGes3uuh8N0mFh176bclmDBdaA2K7NQ4lpzQ9
ZXWmIWyma6yxeQHoGIolGXrWddmqrx2YnUgfMaYGhBfAClLNF//Sud1Cgg5LCgHuR8H/uW1MFWOb
vg6Znsx02p6eiGiEvEQNnf9vDWOPVNq/AsDY10oz+83jGN4LWvJRI/MK7eOyK3e6KeLGp/B2SGnm
Yji12VwBnCZ58i7gAYghLO1JrFXy0jVPrhQHwcjE3ohrlnT2UyXHUEQVvivGVPtwB/TEZa4+LGaS
pKYYDw/X5PzY2MCTmMz5MehhhZWtWWIFM1CMcP7iP6XSp7aqSLQXGhR7x6TGJJvEWQ0rFJZEPXDF
tI82NS9qA1pkbsePJLIKqltKTJDeV4eG1tN8PTzdPXuxxmZoRDfsMRX2YbZ+L4ZPHQ0luJp6jjvU
Ngnm7RdDwYUQ/vhy/jCdkvQVt/Y2rcKQr8ZQLd3uuzaxVa5FGespc9Q/MqmkeHzVq2uUIxGzr/Zh
eBn7AiXR8maFVTzLK3eoWcMBFPTk3QoLVvMOWLufVmTNZ6+Ia9+8eAA6mppjESDcFeegnF2+h5pV
vIURt11R5sFsRO4nDehWoKOTN0TyPGbL7YPpae8klFg28S7KJF2Mcajhn6wsjIZhFTa548UCclvm
blx4S4qobqsCQf92Rb4MfbLkZ4AhCzyrvvPwcbG+l+J7Yux+qsdd9P2UAGiJvIYlOpjF6dWM+uBq
IzjVz2C81rXSeHhVsookJa3Tlex1Z168Dqh7NEJM8ZepST7LWAF6r5FqOnOZ0+Z5GiCbquOLrSPJ
tfNtcKPPd76ydE33YrLa8iF/VA66RY7DLrky5jIvLZybUnaGC2vGT3j0LXD4JH3//RoLis535ncM
TnIZqifrp2BZ0353OGpAjVuvGqr4GbDDiyEwnLFBng4TsE0C2yqm9wY2bwEgrFHinrkCmSmvzlMh
yfevEXM7pOV/O0TVDkGhpY5YNzTE1PKys4UwkGL75rWKk03YKAk+keYrbFbK562vbU2yhv8VYkw/
CS0XSMDxpXVFYbAYmBWOVrY8RKsZgDZuCxBDEtpRFLy51IclO1NWj/GnbcKv5z2AOWAOhhU21Cyu
jROyq/0c28c1WrwS3ooLK3J4pwt39k1Iv5XlGrtgArEUYORElYGdyboNvYb/Xe7rimvXmoPcNG+0
evybgjXq8vcT2Rc3I4eemaVkTV46HPoBIq1KTC6sRxZ7eJJ8KdzbBet7Odg38s9OK7e5syId+7bT
Ib2OxMjNp9BOhg1ZdPnRvFw9lAi/J+bauW6GYoWYvEhWVBG26J4U4UcPGpmFCDQ2qiw8V0KbtRiT
69MhK/SChe2hGPq+4/ixWSrXVS10iU7aD4mAN93CsXFe+N1rVx4I7sv+5mTWSAR1LVa3ddoifdts
Jr7S9/MzpxvsmKitovDhvdWiKOea9WBXoNYUgIdUE2W0VQ85/rGKybDRJHeDUQxiPyjuaPF1GLIX
iUxWGtdH0s3F517a0e7f1cumlEkU2//FLH5nrkvJ8qO7h0qxLlP50zywF7UzOxQ/gdFDU+lvqlTg
3ZNEALFIclgAvbJw/ARbP3Fu7TXIIPA3jUpl1BqLmNkr6xoMNl6JOvxhJyTgPk3aSEwtYV3ZwqpX
HNyka1P5mUjI7gZ6RPuBW5fe6HfY/k7xyQeLBImK1SlivwTF9L7+NTC8kz0I+Deytjgp4lkbe4Xm
c0I9VOqPiVor11NlC/122jb3TRzGaFv54qzXSs8u/yuUoNTY3eNH3xciJwY4rsnRLvRiMCN9Okx0
hf0ENvmPWbFV9Cyy9ezAPeHhFzdPzEgXXdf48Q6qipB1jdsIJkXcIHTvnMROyT/EvvF6PKZZsnmZ
1f/+H4JM5lG6Bz19SfsJ5gtfZtAgIkbQdJuOBmHfMDzQSEMR4/f9MfHdRQXIo97wyHFyAh29KYjJ
gwDh5P3Sw6SsddLhVAbSbBerOmfHIqrjq4XbesFMgo/mHhHb/14DS87MmpkU26q/A1mi6x3wBNqa
noqbVpoifLXNWeP9XJucMB00xbHi7R6lvDkQQmw4M7HTujG5H1ZKL4dpDN6OTLBB/fdUWfx4C+oO
E3gOoTrYGTN+5OvsG84jIHDNbxiZOEWtsFb1JIfto7D3Uc/m9VdbnsHeY+ezmE0N0Oa6zNxImzae
pENvCvooWPv4ec30lkE+Al0YpEIs8VEe8RfBIyhVMDviSEAGA6pTnoC7JvtwFGYcGT5zAegnA7Na
KFafmFdOHYARcXUYcjpPjElmdWCXS/9nbmxdwJg/2rsiUP9xBJxOc7o4xi6U2AIW7CFa13RBjgNm
+e30Q6NSxyNXGPKnbHMkwO5yX5W8ar+Ya0jqkDIFfVjzW5MPbcYGU30AW9VzquuCXlzumXG7Hhsj
/+7/nD40ThOnon266gmOX2aLrLU5ZQ5G0SGjIqQknP/MMe8PFbRw903PBMuN3+ZS61RIZxwiMNEj
wgiW1qeCIwYPk7M2u5SWcdTPaxTnknvhB593/8qqWWuB1vpaCR5KdboYrCdpDW3uxelg1eYwP72D
ZuEwRHzPpZQVe7HPBWnZt8BgJ+ECCf0tMQALsyYkIV4iJxei2aB9ljkMR2qKp0BDWln/0BBcAPcB
OnPSMacZfl0BonHaMkqIUDCDAD9S1eocPizy5Mao4oHV5Dbj8KS5B/s/Bua4YKDgOf2Z3PfGEbf4
4P5bPWNp5aEgnEJ7ADLgXYiunjcPiziQMbJWslDDtsvX6RDDi03buSFJYjabG/rHLYSXplRtunGL
IM6UAk108zZS6dT/ggWpko26O3uRJ6Bzh7/RlxbIqc5byRhdUKVdd2s9fkWdcT7FW1GFQ/CQZ8QD
J4vj59X7FDAlvkDQBOCh4Ktd32YlEap8tL64SLGkhTdeBy4SKbvFgIFQ8gdPlLXWw+ewnVE0GNKI
qp8OckeBno4kW/mDxkgHbPbJ77ly6vMmXcJcBdLVPE1ylRRUKa9nBVq2dbrs6liih6+xvpyg5Aqc
B8QwQgD/xQjHU2+cJYa2InBRGhh5pJTD9S6E3nmwDq3rIytsHSyjvPIjArv2Uwy0rYvp1oAVjGko
vSWIonorBa1peBGWX4IdM6s6Ap97RpQB56YC35yVwTja3T4xFj8a421EQbcBRDC+AO+30zHWuEKe
SkvX6Vt2/jaeYkPI2uB0D+H6+/l2GOw+/UHFs6ZtU/PM8Z/K5ZLX7ljTUV7Q6ijK1ACf7GxZMsaZ
4N4XEjcO3wER3i9gC89zT+HreO5dfpINluVvjsVYjwqUWJwd3KFaoZBy775a37OU7UAPX7vZP3HL
crbeF7QW8A4v4NnBUH0Ab0IDskDq9gRSyCaH3VcgNQwlWhzSBdMQWc/QKs0BjQzvKnyS+N6H3KpV
zQLBze29oXjKAKpW3I/FLSrVqdsF89fWf1XvdEZh/4oWUm4Ki5YuzRiToEi/95RGORmlajgIMkq3
oPFgRkqZINjGEcKAD5o2OIlIpISpotxklkTdiERl7DS5VrLb4D+PUvb4DA/01hlUmsOzZSqNlw7d
ZRZ/aqAXIPjJOl5+VQMuY/Wx7ndGRMtLcNxxUqMec+keoRkYMv7PJjB3M5i9sGQO1cW4mG4TM25F
kkSoKLjjiar/1spms4bgk+n4LzsV1z/wo1NXvsMB0weqCND01gXEVVMImVQjshet1zQZuBaukFnJ
PON0/LvoTedKzpPGawHaWPg1U0+9PGj4zU4CoDcUt5femNBwrCJEnE4jPGxymOUU/Yamm0oy4/ld
MCJsvmM9EgEZESUgaD+fffiDI1LqDL9AVmF95WxKe9yr/K5isrBvGXf0/waP+bYW5qb9JaB49ukt
OpdyVenZiuJx3KKj1KdRxrJB78nIUdmRva0+G3DsZ23Qo8ZPZWNO5yGHgEjfaOFmN4QvHU/lVCJH
XSxrZw/dk2JWOyvZNeI50WJ2r/81wFjyUxaZVRLvI0V7DfkgdkII7+939vJ5SpUgLTrxCwsTizsL
lcQrS9q0WG09ZOx3njJt/cYc/QNM9+PO3yLRUr4brltPC0m3UDM9GdJSCJ9PQ8rrWL6irpQW5QBw
O2I+XY4yY8P15vIcFbbkouZUvjxUx9XVkrjCWExZ/rTbudqjkjmTiBqrHjGdN1cp5+p2evmgqmMD
QHV7E87L8WXTrcxZTAgwVs7UoCHuXUVYbDHk5uCEKao6l7LAzFJWL/FKmYvOIUajxPvXEEozNns9
BNJlBuYMbD9Apl6JLoIQgTGiFwRe7ZeCf6MuogvGCQzjpkmTiQ9+Gm7hXFJSupnfC84PAa05vc7y
9f5+EEGyzHq9yQI/bY6H8YQdsy897OIxajxFAijd3zlxbwJBZsPvJAMpmuGPRfQD4DUNuWIx3YIW
fTfhV/oPfZW4AE/tcVgUzJRcVjZGbBF1ddIvv+CyrWf2xaxNR9oLVv8CbxfYKpJL9m253sEbzabP
cju3uLiSzMvGmLr4RozcCxTJl7ZBR5NG1f0ZXsPFdm1pEd3ySbXbAI4PHNkls9pY7vzr5aLAHyNb
0CRUKxgGUjTwMOd5XW8aCah8jGRsrBQNA0Z4SIVnu9GCL+NIMFxolUq9exmK9rMJKWy/PJGNckwD
NFWp8VKO7Y6ml+uwVTzxQHSsUeKti8/uACsH8zylSXl3Iv/6jlZCDGK7gswqrVewzWV89FVwqQPH
fbbbO/OWNiD/K2qfKHttC8dMZ+nRc0lKTLc0sPweG8Y0R6c2rmOc2fKE25/6XHHaSyLzZYREHcWV
YWu+pg/BxtqshGPaYpi8XIZWF+IJXytrZC/31NchHQULLW+i0CbnEEA+9h8M/aj8jwqRVu/RinwJ
IQLeFDEi5zxa4b0YCa+WvLeuqCL47EvdaITpTWlq+UOVLpVkxEyMG6dOLHFsNCP1jUgbC8TRIJ9L
GmXtLmSJn3QX+uwwm3y3acwIJ5rOgz7756urVOfC2TkkuQ/lXp6ArIejfS4hXkGTWSSWhZDIxJCE
QmoAA1I0e3wPnNrzbvjDPqWlDQN9SS1uz5jq8wSeGH12E8XEN6lzjYIxe/hX8ZHP/YLPdlAGGxJk
ZJMAtyrlSuTzrtZb3WS92bvKB45/j46X69Tr1T1MaZtvuTQp5yKWAsYbUQZ+s15uagCyDRj9oRH8
1iPwpM8YlCfsbVBCzYSP5c/atJ2MUJu+8tXaJFKykNUe22tESyDPk0USqZ0bImbHu6BPouebfcsG
uZIxEgBI048eYrx7WLxuYkTRkPVvMJbb9MdF5u3bnNKlnFD9+xGC8S8m3Fc2+FgElqUEy91n5Ybq
TOw1r1yZ39jkl/O4rhJi8xOSB5HOqtbxqD9tun3+D6DprhsFdzEoNAMgGglF39GTJTQM1iKdOK+5
THUdasYcpSS9SrWBmhembID9iIS3NXAtg/OYvaNhDqdhrLpA7DtEApvGVIrMdhOfMVYKaFFaNsQE
hxM7XhOo5PG4l5dSyfB7fob2azsWXfOP3prwK5wTmTHyROPncyRngFIy3ooDfl4yHEwPLBMGCxbq
W6jOwp5zVKpGpk4kPr+aqNSIAn3nm4VlAWg41RTAqRAdmDUQYVPIKpNsecZ2oSzp4eltrRH0HcWz
a2U9rEXZ/ZiUmtBQawsCfWZp8yJdR6CrDfj4jy1MnB1V/A5zmLEb/WEgxGPZJXay3Rq+bfvk7Bx0
tFyKPRAT45YLEo95HJcd5KGEpo1IhKM8JX+2IpGhxmOSfDDV2O1bJlhzgtJA5dJrYsi5RjJD6CE/
WpnMY6HNbSpp7ReO21tT9it7dnovzxtF/MzgAMlEb/OAt2qrPzv/aywa6LSopuPrq0EVldix+sq1
qz3c3sEnZGaInoujya6dyHybsthG/h/VQKjR/rpPaqhWN4rcYMEmyqyu3BpbwwFq5wZyleNoq90S
guashRLt0bnMxfEO5qiMQY66rG4UPSp7sVC/LeCl5nLmMxSEucuOgejUsZGfLMnZGho+p5sJzyFF
JN7ywECElTStAVTP7S/gcbPTbwJOyiS7UXw1iMvyt7MaKlxzdXDBlUbFkJtIhYFHVoVumSiy8yCj
iclvezf24xbZdqwunWM5xCq86dNqLbAXg0ABNUPa+a//0lZzSbyYMOOfluwFP7RkcEN/o+N4DzCb
xG8OpQEj2f7FSTGhEOPpHrd9M0hkK5ExAp2JgvVYlRhab651XgK8m6fPgeowGQ/PIhyu8IJRY+tx
PHHqG6rWCnHYGL8NhTMyUSnJLQXwXXRqAbtJcS7mnOvVsF2/4odyIbmSpfdbY17sJHbQiPJGrCd3
ZOQuKVYFdqjhF3p5TZGvqOUhoN8DaUp03hRll311EUMcyNTmuPGOyOTEn0bIfU0kuYQW0N+I6LOf
fUgULuStLV4/W72ARcz8s/RbhIU6V4uRj7DIXju9jFluDO7I8RHLqoCHSMsqs9rqIvZGB4NZeTQC
+/qoZ41duFO9K/7kQ3Y+L6DsBZZqgWmf5RH01hT752YLFjZlNJwyPhLCnG+RLeu2rqSr9faLpdfR
tUb/hYUHutrZMnpqC87l4bfNzXYU+vT0qegW5e4VV5JQDFxBjiiwhdwZ8PtaEeJ4jFbYgqY+soAB
6grjqLnkBN7t9Roi9J3iU0wUHJS+Ii6HRqBA0/XaLPp/cwaJGbdXTrE97nRLMogiwAzbqj63AjJz
TDPpko+CRUSDRNy+eIoEjxHpIiKmfI1q6SrMRJ80RJCCv3SqykjIgovlIwAVz1FLFZL6FnWGBjQF
mrkd3+Vv1OGn0yFtsvCP+zxnWUACG6zKyKluXxBbtqDbLnzl2HMKp+xcMDoJdoRnRUpQDtx3tmJd
Lsm+0JF2xwRWLE9NCqh0E305XrfQ2AxeJpnYUFQfuJrguq7B9ZdM7s6CDupWsVFPD5oRBI2ZSp1O
6V8fPCEtUBQ+4rPL5ePiyInB80dSApT/U7nUzDJsxcJUwBWETDGZy42EjRB+80Uyj/DmpZf4ThOz
IMDJwB2cq6unTn4cBC7RUjfEimrVzpx0btR/mDllRwZEZQG3+pEsnX9VIfQOk1og39KrlMVa0qEw
Q9zjcBcfNctK6pMm0O+57r/xGrQu9ffP+nLONKd4ePH8NIbSi7ympIMEWmh9uv160OAZAYwItagJ
XQ7nji9yU9KDzevRviHDa57dUF7QXdJhIzhIJH/c5/CZc2zPsf/P2h2DxSi4UrHnwnTmdK3VmVNK
tm3MBekTLwDyYWcx/3l1gf+ajMGg44g7M0tUgFGz4QUXiUy4eiT9y3XfKvjA+1B2vQPQY03ajiyh
kr1TkgGBmT8XjKnLbx1x8XISL2WJS4ahPvnK9mRp3PYrCfQjMShqH6rf9oSlqhUoixXNuw6+h6eK
+we2L1pRaTiafh3d67PMUlrM4vm0n1GrimeeloxviQqBVpNwyQCZSN8/N2o1c+sJngtiqIcF6e4G
wN9Yd2gXAXdjy/OEFPnGutmDtAs5yNSAlJOAh4e8v2ZY2E4IOw3TTkEphyPpyxC0Cr0a0yzoonS1
Az5mAbxOP/4nHLPtQqyq6b4D0elq+wV+zwATLUSmWEz1IXxobaZ26rbgfiydqyZGtWFaQtC4vnpZ
6CG5w4VxhreHR2nV/Fx0HysbcUwuMQTpftO3UcOAAolaH5uPrEdVYn6j3+4TPm3udNRZpna8o7u8
dYVxeewqWNl7LGKaKbPeTO2U4PA64iP0CN1H4e3olu73Qse5/agsiS2C3IjbicSGBYgOPw35Utfc
2I9cEdvfgio9ux3l+ObhgcAR8Dta11vIlCezhZKy5gkKK5xvzQj5+w6AbrFAFyFopNCGGadmuPB9
njVZRTXmYSkcSD9B1/hoJmppBc2GwMxXcP/rOzEpejLYSMn0AZTyNnlYCSrTlE8W/EW6y43qb8RU
kAzg4ZP1jGt3Os5NmvEGmjBi1hh6LGvjAC9HtyR4+xYtMsf8WGInpu9qRYFHx/CTqCx2G5WeN2cQ
+K39L1hkIWAH7QaQE6CNRSr4Np5UawOBGCA7cdK0wzoZ3ZDf66iRNq0Sc1smFEk4XUbkPDEvdvsJ
Ge9oCUQmDzqeL6QGVBnmpKGZg/9El4VTgxM4LjDItXNwcJOfrEgwYUMiHk9aJZc+us5s5jhECFap
e4XaizYOaMYo865IOb81/lOMf+nhG8bRLvgrTfgnydd9ytRbpi1c44Icoy76+SsgEamGi4/hOY6V
mDHAq0c1pgfsRqnzBfoYVkTMSGMaZ4YTicJPe/HSDn4LeQMZA6DwJBRCkKRGEhjDjCf9NxA3mTcL
xid5XC5VmHbdkYDyYJhUR8UNxREGiBSCTUyOyKmQT7VtlGxD3JTOB/k/Nbthm7n99ls6qLkFsGGA
xIrIJ/76X3cSlMu4y/aTKFtTqtpqW8FYaUeRFsdQPLaAcIHXVQZffhsK4nv28CPEkTvUt+ngvrwA
VkwSQhO26bdNVMLCZBrK84gLw24CZtZ3MS/DbahWTe7HGAhBxIFMMSYcl7PRmxPAqr+Ge81TBlHy
3o32LLOfSgg5AXId45Skb5VuDtmVVyem/Jr/7FonZPR8dnAVAGfP2pKz+D/hQDBurZeom+v8ZYrY
IKCIuSPGK+SX9W47aEQ9rcTGQoiHaRZUeBjOFIr9tp4zGtNLRLvyaO/ZcGb2cCbe/0/IZatrF5VE
AeHPztQeJipkpJ/jNRg5LZFY9QJaE5+9o0f1sWU/OseNFAGIjFjJOazgKKBP5xDSuCM87XiGP7Nv
cOXVDUEPgbfwnLii6SaA9J0RPMd4KeXk+WiR05+bT3aBOMPylV7xyWA28+KoQWGYPSo7quTknv4a
7zadPJU6h7x0+9uv6x0f2gGmCX6gySy7+EmdhKr3RJ9FL8P7HVLmRdhqtmiAtd0ZDbx5CW0h+Msi
VjIf6O59NmoxB2b9ASONYcvtDzM2DxVXEEwzHMczErtYzvIgHnmLjJAa2ALjOHyiNGITCw0k7gid
xoBOmVNPEfzrouGMuU7Q9dNkEIHJJOlxFko7xsspQyoYIoZ2T+4RzUQsulNIy9wzxFDWfKRDxIui
yzyla5g7B0Bc4pGzFYhpLm3344oncZIGhLi/r+kQgUjzxkWVpfcfAYaWRVioAnqN8/jogzHTz5fj
Vqp22bid+6WmmvNJ5cScrbQ2/NKftPPxIB/Ul13swJ4k6kFUQlZmEEUMV7qPcApWDOVOtSyWUD2d
DD06JZiljTCRwIxMDg1QQtKavFE+ZbxSvdE5oFENwIEeRiNXn13amQI6ilM8ZWU4S+3ZleJ/uNpw
XMz1L2ZGwCkl/rMYidC4wWlVBoJOJjyBCkisCycQE0OwssVFDDUMZfUk03WiJmLOleh0ThS9QRVb
LaQq2+GVatNpNtglM3nGX+0vrGVKjSkOy2e7OeaHYGRYc9COHSPv5q2WWmTwd/xZU3wzBgqNzTi2
wEPlStPI6EN9np0euQn9kRhT7R/mvP1E2y4DucIj5pnh6hMNqUAgYzVjL2obpyiCTzhvmEF8eWuD
8cTyHuX9z3a0os0qW/hJDpPajyaV4lGYK0Hppo8YkDXwNh74cJSu8fswT7pr2wgswOqpkFX34+nO
Efs5hH1rIn/OICD41ITsXL45BN2U0A7UwK0AGLtACDps2OCBRlLM9WfjpWDmTsc03Gji04arrDZQ
aRkVWLWSfxNWeN1KhvNSkrxsxi5Yt8D1vewqH5IhmZs5D86c/RJiFnpIHUh0gi/KnAmwt93mhk/R
0WAqAc003d5hV81+yw5Ww5VQ5LKzIB4x7Fn6amY+LzK1Hm/djxh9/cHJS/2JJlLtiddCNTa04ufZ
Ubqgg9Jv7xDkpEzjbbjNKHpJQyHmFPbA3B+alZP57SASqRefdHmTQk5IaYlMIaaiz0976dm/kZuY
f1XWOBw4zMiqksC7G9vsVp8muojqurPG6QrbBb35pkQCEaGggbdnUO5kKS9JLyFtf5L73E9ex5TT
CnrilyeUl2RvVf7kBX7zcIjqOoXALkP0mc0jZjKft1Caa8aoJFNl3faeatxTBD7ur8MkW5NvU3HR
9iU3IKWsmgV3uH0ptUGRkiCsh9npXnktD9UqqQJErguY0DIsHRAj5kxjmbpbB2bWUqewd2G2Og9Z
AnukqawU/HMsepkEPpYViI4aB1ypocRgn1Gz5mTTg0Yv5MyO2UAqAjYYxakYf8auhi2nGrdlzPvq
xFkOL8n4NEZ+b1I1KqbI8ZqcUSflXo1++mVZK7rg3mIKd1pB2n1L5SvPnM8wW939E8FB/VhTZT1x
Abnrdp6Vmk5UoQpwNtpZiIudPdMNdaZhmHj/lIhTnRlIdOJfDLrL4s7MNI8tdXezk20ph9MNqxat
xoH6ncOjAZexoSv/2XuIU0gJI2OeV9LW8d0xojmNXBppME07etOZZOhpxcRV8cgMgTKTtKrTqQ+c
dRs1peHGPnTyax2O7kVppfhGv2aYw8QdFaQHJ7k9p8htbPs6X/5kp9bzMM7mYtbdWB0FOfOGLlYd
R80HNwMP5R92G4lSee6iwDBV01N1CwGm3engktWD5a/+sbKYzEto5TJzp37fzC+6rH1wcSZ5kxpu
pDlu+KAH29lIfOcPrvWoC2N9CPD6i3I8cylB6rTePaxN3j5peWvgHy0zzgPYXo2+j5GMnaVzl05O
gS5ZuXnCuItsQF/TLVRjL2YEduaFqqkNRCecRACtRgICcTmdZhwqOiUttR0431mrq8t8Q+T6eba9
zxKUy+vDgkW9u8LiBOTK7ydx5CvhUCAyMdkcT8tO3DdLXvxSw3ieaNA0ycFv7wIPEofL2MuG07V/
R6zGOZm6ZqEdUnYvIWuSCmUz5/T2KqlnhJZAlbFAPPsqrFT+FWM/qR8kXJWFFzgPE2H4ch8rrm/H
DxQB5/k96cP5wYU8e5ohNmEkESxhkqsdTFSycWR4ST3W9kDGce8aPaas2C9MwlOSY5ER0THdDZD1
m4OFow5adqERkPd45akHM8aIN5zudvsqvAf185l1stjOOAHXFxsfINVH0MZ195+8NP5/FHtj6drm
HLXibsTyUywVUuNjswS1sph0utSsYtmMSYJBcfbOD9b812e6EfgJ3IBJYsyODsnoBsJGoJ0pSeWI
/gux9uHQB0hyGVlD2yJiJRpRhIZyqiXJ+rhqHJXhqwvXsjx0FhWnza4JoBPkcr9t0CCOxCu0x+aR
Mtllg0pssk8GPbSsNgHdsDbV+M47QQsPWxkCWr87K44o96syJmLxciaJNz/ejn6E11hfbeLg1Vse
3iGsFA6yaAMjNmqjMqxNE2PVBdElwUi896cCHAeXAPQtkVDHo0aKyzNMXoHoEsTHxwsQ6L9jIZ4a
y465AdbEpoB0AMKQllDPxJkx8mreuijyS9Q4jnGWkMYpufEnXvaLwC3XWGXFRCgClXcSZA+J/5Q3
QYnowfi3CTn4HYDxdjz3iEu32D6q72DFJ1fgmOcZVJNguGcXa3bcRYNScDuq7jqFoELWzKPvvEWl
ou2RgeclwuqG3LVAhJtuNBHtv3gL8fYowm+CD1Rf+dZo9roAavtCLLkg8yIu1exIlDeqUEkNZ8A9
yNUM4NqiwLIOeKIZo102u6K+9icww5dvoEJtU9FGRBjUMTicPr0ZilbJk1MGLlQvp/leqZr8THzT
S0zQVFnYcI4CqNRczTwdTTCvngKxs4dqGvKcGpKEakmgcwKinNwcSuhqyo2K+y+5o6qfoDT/LjDF
sMtHlsvP8uavEXYuZqj75UCHQ2TSNwr4CLdHeMaj1CCKFIN6TzysPng2s4w+tkQ+ITKLHH+bcNYi
ef8MvNvg5PDJ4etdOiVtmIs+1yczrctYq5U1XfoWz+j+nljA3wJYjS7CQQix1EUasnt0OGoolU2E
kjfP4+/4drJmz/8Xxip50g/f19djB+oq8I08DX0pKVw8B1ki+SQdSeOKkw2zIodcldt3jxA5DrFY
2fL5QAwQonWJBC8ZESpq0bzDDNDcb3OH1JfeVmrLjhLDJPNtDgZjcfp4DwmED4b1ONDfrHvmPsRP
20nGMeNV6wyFYFnMHgx9kO3RTKxyEeNLHAL/I+AuOrE+n8SGQ6SzYRKM0GP1Z+UqPs45e0JGFR04
3kceJMUrgUW/G0ImHK1Vd/w2H3tE3ZqPmu0UYP7JRfVehTi2eOzTQEb8cuAzlInX0TRYJd8lb6mR
DkVUc/U+txc374aFA8qlCr6erWvUyvpy3ICTWveAV9wdtP0e0ri1mzDUU/RmXYWTlc17m9+ovurH
A4ODbsnKU6DOo0BP1o6JFlDL7dxJvB2E36JWj8lvx5CU/CSDAOlYo1brIFzV+nmaECI6TYgqNrSA
hLz4b5k3d//X2RaduVquqZmU5J58BDxPDJkJaSRkEGWm/CfQh3Cf8zvAF7wIAyUr3h0vEivhfg4A
hf/aHiEBAdfSJEoci2tUN1vQ2+sn3xb3TuipG777lsaXRUvNMG77nWCGU0TGEvY+jpkhxjy4AiGX
a992saf0Pd79jk1t9K/PJW44eMqUntKnhddoio46ljaME0MQh2rEfBN585Q9JP8OnPvDD/LSOFg+
49dwiRMDDFH3Nj6HoPvVHoX29lIGkcvQqz+l1OjipcWZOKM98jOpmssA380PhrPe3fMk9fog+BZ4
f7wNGTnMuWCYXFOL8MUi6UkzeIX+HcBf3Dxko+syYKfVALOCiqtazm6Zrl9EH9yBLj53g/HkMob3
xjT4zjlThIjXAVcTbHJRl9VGal9GdySNLYwD2jAVwcyaAiedWFS2C1zWd2gBq/6+85CK13Q/vDqA
cOdXY/SqUC8qdXahGpH75t772y4wR5nigxvDdOk4za28PI9Fd5Tle0cMGWAoBCGMPAbC69sAh6iU
Jk+1LyHCTrPY6gMLRSAlc+50q2ikZRaEUzOybGypxgkYJTSjt676xlSLEe5ihy6Rz/JQhQVhMpoV
F5IuFZZWsyLR2wln3gUQxhR7uQLgF5rsYOAVStPY7Vio1MJhvCoybuF+6U4oAKVJvFLWgQuubgpo
JE3O79/GKA7KNTzR1gnENpnj+qcbf2dy3V1D/T1kTxlFalpHiC6gt7/GcKeTsM7tNeuQ3MeNrlNf
cTWy8C30bWQK5fFcXH0sYW/T0npHfGHZaJsDQyPfkcWihLFJq3+DCqU2ffxFTdOXo7Ruan9TBK9Z
wefxfXzGbR5RRYkjRrZTqGuM2N/+orGAZvSMT8VMA9HdIM2/A83wuvdxuDFznNY51xAkiUOyNhdm
fXlancasZXkDRpuf8YZExiBe2y51NmHB2qekd/bGNdJVqY7a7UWX/+kHnlfCxKtelasJD4Be2vuQ
6/xK2sLe5VVDTscSzfgAdFd5zZzZ3PgYT33ChnETVa3YhJWlmtqwmJonp3KdJBZfcfGcjT9dNjEm
YURUfcAbN1r1bZ6FMMisIocqrX+jmZRsW7BzaRxTqzfwgUC7WhAK6Rm4PorNcQ4iaOVBIiGhlPgX
DLoDOVg/gX0HHGorhjrKsKTWGW6L8zRYyq2PI5t6gLzZjHLxRrcv+pHGgYbyoOekxhb7hvWTWvtO
dFVsqyQ560TTSWHDPnVCksQlxKisVwUlIvJ3gPh5+2wSJI7Vp3Y6Pg8T2bc1FO11V/Tf4UY9SSG6
6+d0JNYCTPJIzod/0MKiPvbqvPUfYq7bHzjoMwlv3e7z4U6jy9+cino+qWdvtDWqNEaR7KEgAIow
8Td6CgKZIMOj1U69We2U6d7ZpqO3Uiv6qnC3C0mS0yVaDV9/PPAlp/AZ9xPTLi7fk6RSJYXYq0ep
TiLnkWaWpwkMHewXw1inxMIwOtPax/cYU30Twqx+rYLw/Q0x09uKb57eshbwMUhzyxhYfPek+cLg
2m5EuZKWkHYyh9pXiOoDnsWf1houGukUgbsQfX+sile98zpj3sNLUw9M7y3Bh62kE04kmU8SmSlN
v07jq3yguPS/PrBv8tQqiummjGFKkzWwEebgi2UqdJ405RU3ZVzw+YU2zKaAtCccYlWKzm6aP7tu
NHB6OGhu6ug0WrvNrHMaJ3hGC2oxICBKTmIyeH0/DWvXDxvnrUwWdxTgN88FKTz2LyJr59fpswlf
NVG9cGtRqCMoiPZ9TR36kmMwg0QBc5R/0A0e/DUiUtJ5WcVbzBf77x4A4FCzVnB+BD/OypQ3mWM8
LJYKh+VVAauzV47T/dRG831Ta+YtYjDjXNYBKJrHRE5Y2lnl5oe/qwyIxx1Fcggr9VJhZMhYKzeZ
PjceU/MCdRnA5dYu8HDWkg6MXL2ALtG8k4ujk+9TUKQGlETHmmGTVMXcLafBh3QxSY5vjF609XBs
91Uu9KKJ419rYebOxUYfR7mS9zCOL+t/wwGt2/mrTPd2wZFZh2NqZqUq90iQ6cP0ow6SqtYMBXuN
1DditC89s1acEuCrE4afT+g+sQPgWATmF/l0IacycAZVnt4pv0DJGU6kv3wTOXFuMctjkHVKI5Y/
5s2xqxnsDWu/mrWu8ifh18sd8TcfCrXJUG4MNZ8htsWzikmhnzjURAMBHHT3EhTv48IDI1QUEoQQ
DmOnHAubO2GEBfa9b0UhAucue9uSBhPyIccwBm8RnHQgfl0NTqfC+9YIYhCOrWEts8pWmpivdgLC
btEe46NQOWl70ouKdqtk4kgA6qeWXq0iUO86z733JAnsJc6i4tlPOQB2AGKzXBFkLNEv/CZx2Ek8
GI3oano3ICDljKbkur0YPClMbNvVVfeMN+tMBAXcZNQDAGZRwp38q9SQ8QpDl3umLr4G5tC5hQqk
X8Bri33JTOOPpWn7Lw79whuCPNf/ec4rxDox8b2V3YUg7nU7UPaYjA0J1pArq3aRdQDhl5Jv3iXv
vNe84FmwIWcOz0MlB66wnniHQuYWGYK9yx9hLbykq9lV5FG9P1TttxFn+Lq/D1NOba3Ds59QMvy1
MzOwT22uLRogMDY35O/cw5R09XlVEq3KNOm6gVuezCn1zYMD2Rx/Mo1AN6TD9a8kr+ftrgTPcxT/
7RWvwaq3BhSg0Ao26nGTNA9DZ1gNl9v8GYaqhjPNY10HrC22WOqbqQagq0tIfyn4IixSMsWvaMIT
KUgErcIQOZyqnKY+SO/DpOegwKx6wSfVx/k27FLQRphIVvGc9gkladwdUWXqgD2s/egKetCOmXPq
tcSUqQK9+vnhS+uBs1VqmUg0pY4O+aXJR/DshH4QMzrFA6GofrHwD0hfxverYocSHIvQNodRTTws
Y4Ri4aNP+tuDP8ZWmh/pp0ivuejJBNDkipJuTFnreZcOwOWqbY/Dli3mdMln27Y0LziQwVO5geTw
MhpXRphwHO6zcMJOujz5XX0f90eloKMfbKnz3vxfMuSlEryFA7F8dlzTFh44jECyAqWx3nWFSOyV
mIeOeJt79AiJM4uyuZuIfpM8bktCmSnz1OLIt9FeqQcacaCKb5BEcIFtjI9CD0vjqh9utYWIgswW
E2qza8gOU2AxFmamIcCXOLMY4mq4CKMIDXXccI4zvbEA4ka+9dUCqwNe0HiXZzV+2qQYrnUx5X5Y
OCvnpNgcASrbHFsSjVZccvmBSXCMTC5gJGKphJ/aP2JlbrELCoME5tJIOlFph2/EqywqdjdBukwX
mqttvfE/g91uW3CnO3RL+zP2wn5tuPxo515kUqKVLzEW7bpYttXSYQtvillF3X31FBMSKeRTq20j
zqyQ9ypwTHj19S12v2aV4zt6Zr1C3nKIYagggogacZHMJn7mls8ctKuzAp1TcenN/bNm/F/fvQaP
lxNBtNHhwVdh2C8OPnfho/kAXA8yOuzQsKdrvNQKTqnoqk8H6Wv4q8zrAntfSn2vKkjq68ub+H//
51QAIj/CQAuQRBYLSJF/fRMwyKmUZXHKUXKI4eZ7+pw9J8ohcJanY+lW4qMh0JvzXVhoC5Z7lWEK
TKnkS8yOQFgxTlw61dJSrj7GvmygcDVb6vf16hkMoAJRRfgQ7aaRJ62YydtctsqIVzAQyXmNOFIC
Oe910RZ66yGHYlcizhGj/6ocbD7MBpb/EvsW+nGdVVpj+S23ecXFoEC4AFChxCNkuGBl5/O3F2rM
XIoMl92JTqSl+d8EtsDWgvHyxEiUljms6xE/39CejA2F0wuSIRyEwCywkr1Gz3FuOLUdoI4wMJS4
Jknat4S4Qgo1Nk8ipJTPFOTj/idqNWeY0Cyy9ncjsueNC6EpE0W42Omo6Gab/IxQCQGRoyCU+0ke
Fi2e34adQGcQ41yq5scVxnhzqNSDAo38Q8LHdOS7fm254LOL/l55lzs8ce9Cos+2MmXCI8TiO9Bf
5/glGv4mUf+2wKT3gLhucLJA5Z1Y7y6MvHvNCUowm5qThDKDIiPWX3kjkuoACogTZNc8Ng3pYwu3
mJjPHBF42qSQzNugVwssE8Q0nvTDHJiI9Q6GBXxCEIrppIGo8NjKx0DVAW5u9CrFoKlRlIE8Dl3h
QGBEUJNqHs+uEhhpznLyngJtrjwOsj9/JspUpWNuNQlA4ntHAKvvRjgUDxkNHFNjQnqC8d2AROYV
kl7Wy3u+PwjlYq9tSfhGrdTZ25DnGI4+YpZ7KEAo1/IrYkLQX/ekrzAgOfn2DmHy6wxSHg9+oryj
+BuONgJPURzDS8PqwITGBDIRtLTGMt7ar+z7kVO15i8dP3C7A0fKpO4E+whmA41LfU+1GFL7bd9d
R09NG/V/5d9ZmeQ2ZPBYMYZkYBkWTsMnXNZBcU+l8LqxqFQkAUKV1TBemSeACfooL0sGGzErEhgW
gRWKlWDAFY0h76s1k1QFB+zojSHUJjHhugWWxpEs2yOnKLNonyYfkbvU6gSwKskC7yIZFN7mvvnT
hrFqadu91ScTQ1/d7NxMCustyJysVPx/4YtR4qvRrMsd+e49Ow5s3tz5V4ctJis+ZyXMbrClSMbQ
LwZjV3TVqTwxqMX7f2sYS7r8nlGyH/BdDcC3qc/5fPioiWd3iEr4QZISkAJ2fRxqjnoj5oAhcKew
0dJ+XkpceiGWuth9zsii42lLyh59IaO2Dx7USp8XKLuiRsV9CNIsdRExCWgNzyG1Nq/+PHNb6qjg
1EARt4EEb07PSshnNfRzWbHHQxJ0igH5DaETqhsdTKntCVmX8/lHS0pdio0VT0UsROlMGwTIe7yd
wctT7hNYDfr48q6PWdPEyDozHRoXBVYk0pJ5TTY9GfWFiVYIliu/mwUOmGN5usu6aOZdtutx2+ig
ygL3Dg8/IP7jOLcURrsZ/FIrn3qXPRWSFYce1BLrv4Ft/WNc3E6zYT4mTu0nWmmL2LbwH8TxeIIE
kAS3st04+hPiMEJoyMWK5nyjUC24qngx/FIzLYtrL86/PiOvEmW8Afu+UG3eWvtt2GFqPQCxRzYq
6HETqD8a/ipDZcqS8O6QABSRgKycQTjLTngzgxfTjNLXpxnyBJGVEGHOYIK663NBQg50lIWmXlKr
FwpE1/XfLvoifsOXtvHsrVPy79a8sgpZZ3YFU7tvbt63XJ+80YYv+p9LXcPrvQuQz+yRAYuZ8ZXv
XWSfn6CPCGBt4HVFJUtqFAucCFqLmJT3jEzokyVJki6PUveWUefaZfEBmDQLPUBd38ekFAi7503W
vOJxUKV6BsE4CxYjr21DauIf7iaZh9K/o7bnKVzBqPbVBQ28L+vPfR8qd+hzC/xXESwr0axjBZEe
HiosVNENotV83JWB2zVG7K94QxnHvAuZf8v9pMPVGu+Xj5U3TVvarAIQPZW/vR7iCJu5ED9tiItt
AQDMjh8gSIh8RgK5kt64qhGkw8OuuQKt+5Pcc+JstL4Ml0lehVD4jtp2XLfqyPBvRgUv3I9T81Sq
+uCjhX8M25cmQCV3oq3tkEwhiU4dMBgTiL+Nk8q+qOesthUwDwseul/I7sTicZD8/jxK1pRQdKmm
JayIz4AQ4QcwM7NRCQxfg6ZYXbbl+C99YRMfZhVwbSpJv2P9XNS3eIqrwFIdegmoeMD7t0YozBYR
bT9gwOgeLZ11zX3D/uTguF3gSIYuMnHHofvQkWIRiRyxt9aTpECRR1q0wKiqNCrIxytqtDQLETMS
BueWQLTSVQoarEbUrdmKyNsakAnglu8/hQRC5I2nPpgdX7E6omp1Y40S8SOKUaXCZiutZFJaTbBn
/NvHijUM1mj0BB9Jc+MJ83nEa5Zf6PVEyjkcpkC4H+uPQoOnh5qP+FotbXlxUzj+StFTuWlUE02/
9WeSqSTnPxLNt7JXQHJQjyTtXyBm1DgnUi42wsrNzurq42rhEV6tDd0Hi6oTOkZK7STz94qHhtq+
NIOd/kLcu5LxU1wfNdxJQ8O811AcchUSO2nXi+vVXa13G/KleLMtz06vWJrXQXEaWpWKTV0jnvoE
kaHz4gdVug4tMf4s1HoEG/XJVobkcdKmTX4at3mNSAR6rVmH2I3JcyYErtbSY+NcQzhicxPW5gI+
HzZUJE0vwmpnd4AkWdkFBDqfU5XVJuNOsxeychlUGFUypMWxTOxzmONn1qUcRm0bCJgAMqfNIhtE
jRqGJyP1UgD739Vhb9mgHTT/2A9soQVfxYyFhTg+YIJscWdEI55UrBLKp1zb25+VnYlz5zKUbcJq
rz9MZcnnthBDA5ktqVu53uv4XRh9iVuxD2hNiXEk0R7GgcVp9ahUiNX5xEQnTSxBHGuSQCHH9Lj2
AW5DJErKa5AaYvplURHv8488C7sCt2pMjerP161XK6kB4yxVTJWYIfoaySr+/jdeuPdRS3feSQjR
Sz9E7INxm1f4DCtmICajjMYwJhJ2r5kv5GKJeC+2/3bhLNQePNTfk80K/CrTQ1cmtXdzEWhuWCn1
bD4nW40lVIducpVWgm4nelcDIye8Mh+agnEu+GWgwpdb97CvPQFw3prY+guFaaFq/6CbNF+P9ZF4
lYaSB4E9pKDlE8b1ivmetLRp77W7fRrCtgxkQ603p+LrGjQ0ngenyQ8ImdCXK4YSDnPjWV5MWBMk
qNJ2uDa2FNDyleek949iwdsC2Vc0VrEp1qHvhO53xPDvEC7H7IkN8piweM7Bde/bK93GEnczKEVd
WFpv53W+jooe5XXY+jEbVgOxrzuX9J3RsIIyUI0kYi9h76owfVGSzRVahp9YG92K0U56HQr93zuC
FysuOhPdU6759lx8IMBCCwsIbuipbAHH05MM/T64CQYobL53BkOIt7gnkxswjI7g+GIeTAdLlnSH
Acb4aAFcfq/h7KU9LpW2LjG/TTbwRzc+0sjPadRssJITSfBH6OIhTVTCWVzLJWfxWp77Q2N/w7lB
wV8FL2ILPedpuVrUvsZfq7USRJIbr2CNyEiux+1MiBuiJAGBJ8NKdf2yLw3l5KO5KXFMQPlAhz+o
ElkFEOy8BaDuJ1Zc5wPMH0GmTn4+8ZZLNulzcKBNWPAlOmoi9RJDfCMkS6RYm1gl037Rr38GYSKZ
FZQk3TIsbQZ7Jo8Pj2mnsE6vxC18wq9XuyOqPUncTSYviXj40R5VE73/kduhe5s2pZnR34MnVzki
6Dg5TrTLJIYKwVzpNY1qlyflth+DrVP+a9gRm4LwgaczMP4/ezAP913bRmsv5HXjgKIRzVetsnKP
JJtj6zdd2VsLeqgTJqwXVF7YrZyteSdZ0w2xkA+4jP45nehDYLSm/JIhddWvn8N6u+cUXHWDBtRf
/Tsz/WJKFGgJfPpOLOtrbsh7enEm25tbvnulbYESvDX4wXUDJcov73D5lAyoOeeh0SBeAGnjfp/o
eTx+ymUSVnXF6QSV/tisiwJZ2dpGZp7gKpW8riz3+j6WVa6R/qBiH+207Gxr/+IyKyy15OXKHJ0H
IG+Ls9p8Q8jhOIb8ZqfvQklbxKSwz7UK3a/FMl3E0hbWbQ3JpbvtDCX2oltdw+G6mEaRsChAxAR+
n0POTpH/TC8V93w0FclkZoCGDASj/we+TqYSCJclz1+Q+E2bPWYVn3gX1Lg96tREx6wMphHeIEyj
IE0O/ZXlmkqQ320HMfOCBbC0aqh34YYNRl1Wfg+wWsIgyJDwW82jlM6BkQYaIacqFpAG/RJuv4On
72PbhXwFL8y1jcNFRLN/oLffDYE9IZscEqOTY397PJ+z1960mJNfB9vTFCUGUuzX7f7YTzp9JneC
XPIVMQNtkUxcP19mLoGp7U94XXq/m9EG3Ui8DYnKZUg2DBaC39ZTjkFJ3QiA/LtiWcJLIKy+Io0m
hd2IR2C14eYnPTSpMpfqkHiR+joZnBFovMitKf2tZaOz8eEs2egLbyyFOwYoFMUsYRfondSbcHYA
ulhCm7N4tS2nwZ3R0to5vzBFqmdk7EYyiPTXjYA51Ct+YvN9c4o57sDTGmGttAr9rC73zaU01Vs7
JkiFQ/2sKpejXMZL6rbOYC+0cy0PWlJMsy+mmnqef3IcZP6S2ym6DLKJagd77yWxX9lJQiH3jU30
wUIO+ZRuM67sfPuR89Ai1JpWZwIdKhmESS+4QhnvAK505yzDbD15zIgBWib3CIJ6H2o9uQ9z+nX4
u3s1wSIiP21/1+p+eS2WvU8x6O55G28IEVKD26UFXrgwLSu7gjZwv19np0CBJiJgBGILuAEkEMWL
/m8TUO5u7+JMc1hc0HcG+Mq/p7jniyjjdM6i7eulsHMgIQw9rtrTyNv2aUtGsQdTx/TmGQmBhaOj
MSOrGw7gmo8z6af57UQ/rT+fySYp2JC+Y84XWF+vo/TXEzqH8wCHq6a4Qslo9vVBzqc9RWHEVoBg
AEj2L7Xy97B4b43d6crTR/4U2tHi/hckpOimYMBCI+EMV+KEkHCtRJv+uah8XY6FOgG3swyEUB9+
n4rp3XNB7/gBqKzV4OLWa6Lbmbvu4ZBPoMXuw0tsEQ54BrDYkCbnW/UjNIv0AJkfMMytWOJ8HLlv
1A3K+rvSpgZD+Y6Tcu2umHHneL8gQ5FRH90qkxe8wZtUnruT2t0kIMVHy+ewZN3SzP3RwYCrUzm4
ZG6MUqf9mk+yX149LArs4ygC/K4sXYpglN6rEgullfY7hAmLwFIAdIi1hsQRB1o/HuKTAPe+rkB2
jtN+Hqfq+NvLkEQ6Dg7SjpS2E0a+myb71USUVD0BpSosiV9b7WmkF369ZwkSPwJFvb3LJbpvi1dJ
rDvwnS8VFzdhacO82motMIaad1eDX1pz0NESWKYY75DVP8jrqNY4ZZo3Wm2JV2jU3/Nde16iRWgR
2/oWSkEsHqi5QkyM+Y+ZVO5Q1azi0TNMUqdSWQdw846JjtWKMGMdnAvNCzbdANAO7bNPPrbMFhck
BdqGrDMO2XFF7UL1V3CdrwV+Bz8HEAJhplWIpvrRo48Sy31tit08/EltPg5+8zNWPgAY+8DNITK0
RpReJWkmFJVAzF7fKpz7YWBkKTuvtoKbsMhNtZiZWjCDUK73DIGsMWE4h1qb22NvmcyxOgBGSdSV
WHwGIK1qD5Pd1/Nzst8swk24u3nZ312DkeZx89Ur1O9q4ioqeRYFjE50eAY4ErX30NEAEErVMf4M
xHQhv1rUbfxnHacoDsn0WCT8EyKcYX3JmgmWZhzUZoQbR3FLfzm8redggwTFK+BzPioZwFP1gLbU
VstL8fYKEPkjU9hFHJBMwVrdpyM/nbw00RmPG7M+mR0VJbyeujRn7AIHePt96Ydae30AGJXnHZWs
auOS0apwLQv+9/ImpqNVBGdxoFw85LOyFFN8MhZTw1+njJHVofhm/mU1QmkFYNvp0UAc65H0sO6F
/46YT8H0Pp8hFyZrvDCAN/1ns+mtBi90j2dscjOj9n+e50KoTApF4Ebiy/vl3EngXUxAuo+zF/uh
YB4g6qviDKwUZ4bfKOfhZ+EqoCvuze9Z9S2oXIUJoeTM9KrQUOl1PttxHj/clX1RbsooSHAjdfaU
ax1te7M8YXQHn+GvMmilAPoNJWUxrAx0ijEHsQ7055ePFDOwFUP9jLFSDnnjFkZBk8fL8NBnh0qa
2vBzB+XouN5m/ZIE0TEZQd458WBjqHvBusHDZzxljf4agJuN4LbrIuoPiqP9/0OwhEvvF8wGVKf+
3B9laun0RAv8JCzBNbqhrEWJ1YrUWAdkfuSPzf/qQIgRfHciK60PJZVIZibDTs2wvcPdHbi94R1H
9dwk0iIXcImHAdMvGc+WVpbDKZ1onRHhxuBR6HXuq4vfKfsRF9vVpJ7gi4EwV/3nCLd2JhJ/TSyC
j0sbese8Xdvi3PwiJGPchYv1nOMTnUUWNivdsYRyCLqRcWrQys5NpA7o1fqamY8NvpiJVhHLVA1o
VgKnlYAtr8ijs80cuCJg+8HB45FlwQ274q9vfqxhYUIVVl85sUUcqONOztju1Kcdx4FQcScs5RjG
XDUpZpV50PvpTEsnpDlayC30ZNOyn3YQ1IGzfviMtCk+w+wHgN/lWwCxQyj1Y+oADQJqMGlNEas2
Cimt+DdLv13rfiHSftb7VMu5rtOwPSLDuzCK0WPQSgSqFztwcIVo4mfjNf7LD25X22AGonTuVady
sNN2VwBlMxHJXf9FcsEQHtliDrojhHFZVokiq1kDWH7cZQg6Cssn+3dYcFBbhc3BpNfDXaRsauNk
OrvujsBk21/XPrLJjneWZt1+zOXNkOADM863owfb8MJHDyxsCiJVirpDNX1NBywhDlfm5BDNaqO8
36a6HqTta9jhbgB4DFPKz9Z61gpDLTe7oWA9+CTofb4whmKDL6v1za/Ux9B1eGdCf8oIiRbt8dUO
68ysFjaITrIs8e5E6JU6HtdN5frlj7pmKDkalws5+kcHt9ymfwcVVNxau9wbbqPOl3TfdGCDssQ4
vh/Gpvazp8tyCZRQZvffFC4DpJVBkl8nAN7dg0tBiTSYsBgCbft4G4mp4Qnm9d75I+IgyMR61Fpr
PbwjcRFi8WmH7nSIKQ/bkOkmckyfRPec0Xvn+vALffXIRZiC22Fu0NDWxb9F4TZfpQ5zg5EKfrHx
G94iel4sxZDeVskGkjiActWExR+poHhPAcPjOPf87QtiqL0gD9OmS0HmsmAfNL/COKEFkVr4o8v0
GovNiCdeXHtiTb8oqR3Zps8CifLsCZpdurNu80mFNPfpPz/rCxxNxNT08ZYI4LtAlRx1cOtDUsrJ
hmdEi+alABWJ+ibe5UTSAPRRLVnqYB1mcjD8DD/XeJhHix3Q5Q7LIV9y9AU01Vvp1HysCrHzle4T
VZRZx9Voey1zkw4VN9okZNHNPI7Eml4fqp48HmkDG/q68JR1itPkd598HQsHzbgixFkcTWZ4LBov
735opFXWrMl/RY+HJCA9LFGkIoF5kEjPjswBTrZUMV/0P2982EaGcn6Q6Sk8/w4vCfkaE3V1MVkO
oRfSZrD7QsDSbeG4IE55wEs/IqFwqpIf2eL2rzGfynta/mLN7l2eLzm1HNlqCMFNrsBVka5Ecu4d
G65Mk2oFDe1PUPQLN6Ke0PjdbSdxo+cR6oziO1hmw4XlJnzy8Bb3oPefwGpdvMDJFlUUL/Y9Ei2U
hdee496oqS/ARPBbNWuqZajcuOLnqs1qbyGUcHLIeXZw0sxj7ZqWde015ecyUxCc4HVEsx0y9x7H
9aOTH37Ing/jerFPH/JMFdxE0u9UCuYiB9pBRqKMdW4KMMFuRqiAdko/jG/kLSpfTw3lLf8ARgJj
Z23sIKMJ+7UCqJNj4t0L8WZTRMo9DRf47FPHJBjvxq1Hth2V/xQzcqh7SIZ41adqB/pr0rfCAj9z
9xfuHBqAtvjzOyedwylfBYPjnwQjX5faYV7sPCPTjNftgQ/un57cxE7xSCpjQeDiRjMOyAIRqzhX
JwIEcRGLHtaBK3VOiaWlrI1N+FzX1CzKur9fXk4mW47UFtakQka/8W1rtdeyl9Y2dCYfUHfOoSgx
EcQ073Lbcd0BwuKnSuqtZan5qsCam/q4pvaN6gKl2t7AzoRDuE77u1gfPGQ9uxDnrudhVJzRM4BO
C4Up4cKOmJSQEAT4mDnT2GOMUClqiyLv8wDgvAOsSyuJwZzSBetlGVBBBNcXfzfaiZoTEx/EpIxD
xxgcMNQ0Ap4xkpPZC7IEy9ILjPGV9eDqZuMtZFHk/hi/bHzTN1vIJkELB8PsaNHHd6EIT21yPHwu
r/z7zUgeU7cWCAgFMYPPmdHtfF5+GhYnjqsCMvuamdmkT+w2jhu3IO+rDup8AWh7dn7isPZL0xfd
+bwaOj66bUefQNvTwolnaqtE8N9liQ1CEKGYEYZjNpxRQQKNMcln6e37Hs7fTXNZRpto9cfk4MZy
zgvEmsqfneLZWlJDXCOcLWNGHUkHDShxFQHBcpdaqIZMeSSkmDbrYY4t3oby41ef9ht4HyRAHzcl
fqQk0ce+LaqMNQ19f5gdkf2hNqlha0RoYFqKxMaZplmlcnThquDYweAni3zvFDNeqLYFpAb/JqSo
djee0tsrQg9O1WbZVBF8PpniYmo0zyx8XUVcC5d6Ix+jHZLrPjWVRdSesr5kjljIPEumBrPzyFTz
WT7zLV8myIUwVSQTXdsv9JPoFeyA8BYZVvFDCqQPstXu2+6Nv+/OisMZaPpSFCS2LGe6zyowC6e0
dpmUFc4a8O3tFyziKh0+Pj6NnzGI50eyo8LCTESmfhcrZO81AHKC/IXpSfPwGN93EM32CPsYRCMU
x+HlyeAQpcSooCYUt5YbbKs7ZMYGDE94X2ooXMqg45ExzAEhYpjetQOXEeLqWHZ1PwxT5UmAdtZp
VeAK/YkRlSv4Zxd9Koie7IcW7NNwOn1AVVntzgLKqF1XZVcmauwTfScYqgbuvwaHHrqs9e1gc4R0
VZI5aV+GgZ6IjQIdQJPubTgqlWBew6sBCQS3hFM9GHFDlUR6loJn76DdFhWTSkZw0w6gdGICY0RK
/AHNJ4RHbPr3zS2Jr7HY4WmjN1GuIm4iTqbalv6Ido6c7He7p9j/QuueHLYFJnLbUrBKFyZcw0ee
2CSZsrdilTVcbVApZjUeAnmnz5Qwgl34U60vKzSlLuFB9UmpF2cjmxDzHAFT0+e+Xr7ICu+jDHfz
lxakhhs8S9YJTWUN5/5FAjG1s0BxCC91T2O8ipBAYdnnXQUWqLjRYqylsz27nTQQdXatv2cq0Tkb
jJWciN6heGPjRk6ReKVjLBWacK/qnlcjkMKhVu9DhSEN0ikNW4LVxLhN1vhP+sNYMCy5oxS8n/+e
qx+a2rBv0Me9XNI1aLnhFtajbJpOjyuYEQbQUe47RwS5CfER+DiVgUkhDHqRocWyED27h479na5g
atIBORFYuu060mCSyoOELfdaXYb8iEw4A027TAY/qYRU6zgzPnhBzx6f/ndD00BD6S7JZgpV7llP
+t6YQFHXJNHxqIxX+oF6La6sxI79kAGEnWxoiFkTiSMVoWpLX9vwqWK43Teo2qD0Gxm3hTCWTl1N
X42xHh4rvgBQOWN4+JYzA4GsMHQgjGeJQa3DHV2X8lwqB8gWnIYEi4SssebWK2aWQJjpyHHGp+3c
OT57ZdajtciMGEciXAn4FBPnE7mEG9kjYbmJMZgz4qCEDH2Oz9Ixkx79xK+7x3tLvoUV26xJBTu8
lFqeFKvcyl+3ZxUEf3ysWkvwnOUH3Z053lnLgNBxLr/x6rZK573ZyARhKe7P3yzpxYLBxE8pfqVz
BvxqRPkt3QggcYe2fFmAjuEQv1GjU0s7/PfZnxe4+yn38PKx6hRlOjrQj/BTI0q8c/2C+fZ88iwA
eX5UucWzInKBYZBZg/fQEhFkGDaL1i9jKftLfjQD+3BkdRkMnrSZGhtvRHy14az/DFIDihF55+7o
GWpcZqkgJTIG51ab1gZlBCgkvf/GxRcZrKmZdZWiL92rG576fwlAjm6c0lvL8A+GxltRC+5YjrEw
dCLHuMS4nI9hyBdHxryyCfBcvqDM362fxhRdy6fpRHOag97KMxcvtPKqpA1ybkSs7PVj45kZlhzc
1Vf9QIx8RpqjYspa4W0kR2kFsxZjOIcXyB7pc8lrtS5FTO2WpwOqSh69kk5rKC7WDtJhAtgHj62Y
0DFFzyY/va6s1kk5pRQOOZou0ZToftkARfvu1553Lnq0F7w+3fwVc1Gn/ebL0bzEXIllZiV0qtgP
NGGGHI2i8Fcxky+mqwx/ICkKrUNfPRZnHGZLkwZfMFaNYz5X0OuAt7sdna6qccgUHHa+EPa/mHWv
Qp94xHQAM1GHIzVhaYSKmoF4vpEMkkejxj6+aCLTfzJCkWQEIjltF5SEAw5VphcGzbNFHnVXy5PE
Zmp94shPRTwp3771kWrYiWSfHVCRX7sj/JuhpKafYR4LU/UVV+hkZmdKKhWNSW3HgnNySOjUb3R6
C83a4A7nHsm3saOctgoWGjFZYzyZUk1r/rx5uYciQihy14v8Xk07Kpnj4PLGXwoDVdosMPGdRspR
2fWJCXtOPJGHynLpUj7PvttF/uOpI7ZAsEPbivrYYJSo6UzC5tAd+Mj49RRGZQUGq+R3VZm52JuX
88lV+vbBcX6NxNnw3yuOwTU+r4O5X6S4oyVLspxhlq92DTrBsOvvrKHk/zsGhnt5J6hDOhm44zog
cvnbL6NiZ1a7ZuVpB1vrEWhVN+2odqBphwyqpkHwv3Pm1Oe3KWdjibBnd3gHPELJsTjJ2iYc7ski
lhZJHbGFhzGwyzrx0PjmDFX3INHi+MtYK+lnSTc8xnjm/uM+78eLYtv+OVij3w3xpUBalpvDkDfm
K1jIg8B4/5XeC5Yn+ok36onhKSlUWKCtEqNj73FelCpe6KtBJvtsRjBjHnqfHAQiWHawBpU40MZo
1zFAQJG9wrb//+w9DYwycjfL/J/1etXPMtUbh1aMoOWrguh1DxpCiVJT0mru+orhnIWKxsQXKSiS
4r9xc6bwr7vQT3TQUi2JarWuGU9StkRChMJSWjCz/Rza/l7HHAN0n7p2Lyr2rieUpR5tGekFBq30
8nCDenhls/O1vo4bYdKvNNr0H0r4+whLpcGIcWqZfjNiI+oh/Lepi38Z33bOEosfs0yE3Eox+br/
ejG7vQwnwmKa6abfK/Jhn7tP6CNJKV8Px9NEdJ1q4b9IBpFtQu8yTtTNwBX8h9QKu/k6YuqtXrpt
x1EeqMUuUwmaau4xl8Q39astXY6GBe9Q9noKx7g4KRzPvLdm3VX7yfC/Xo3R3qzVgb8rRLtP3NTy
ocwvHdTjEJiM2gfQVkTC6CA0+kaUPOKkdGPbNJx7gmEySfZT0WHwJaVjUlxzzji4EdBYdoNLspY1
IQEwpmC1Yz+1FiF/bvLoT/seju1jDzXqmOf7vJspv9JzKrLi5gAfQQKL45cSeJCbdmeIvkb1jZQx
X0AG5Ndjpl3ui03bnx/KeLbtMcdHPx6wYwbiJJsvdt7Z53F7v5RODcW2PeG78IhIRp1EA/86V2M0
FseioP/NT1TBXlTHu65yivRMM5XH8TbatDNMeVH+JwafdbO/fsuyMBnRFqosuCVmP047iWbf7c7l
i9LppDZ7uO0E2kGCzrx4skL9erawQrt9xv1KANk46TQ8P5jBZsa+XMkL0ysQz/r0lNgZM4JoTyw+
HpSHibMNs/ZLxQjyniPaQz5mqkJ04V5LF5R5d2PXFGhRxa71q2LyqweCUGq7hRw7jA1FTZ5dyQmR
wwDMvdseIvo2j0g2KxaZ4pqj7aptwbdQODUuc7le7VJDc5LOpP5dXyzYTPD1h6nbt7z0Nag0Q0vy
H7rSloPmCHk6NqUIZcmgydtFVdoG88Qc7hrvnnF4hEx/oL0PX3OrxpMypFwfW/AfF2udLcUQoDLI
mEF7rK6EvvfzgMRxtSF/bKhbXWvP5h1yvRrKgtdXdVRISFlsomRERO8k52KC2fzRW2dUOpKmt7dv
wPUmNvKTBz9RuNOT0KfZ997WPUS/G6rcVQt5uL3/vBCPZZm4pkfJ1zk9Gjk69VoHUSkw939zTaXV
A9RrS4FrCLMZhmHGcwC8U9eLqsp83Z6jiYY/lViSTR5DUeVbGOYWlMUHaPx5m6siTDsy1jE2tHLv
8FPJO1Q2jII656h4roWeQG4nC4rUCQpL+b/K+TzKKVMUpCJz/GYGpexTZpuHIL9IgCUClxOwhw9i
WDZOS0dTNR92bICY9Y++EqmyzMLYdgdNcz6RjnV/ZkKqoWpvT2CeKosIZpCShihlYdfCeNUhRZcQ
lyrGA4P5vILj4+v7GSKdB6gqMzlxnuKGMINYuIh6C5j8DUDYvTXlAaEgpf8Bn7znyzPDlReaYjNr
PYVwGElHp1cwf85i9mPW/iUnhE0kyW/ZQ569/pbuHfd/tRZbH5/0/29Vu2lFly9ZZW+neC0YJG93
qB4ZNWgz6+hm1JLM3otsraQxExi0B3xO6W9n/zR1qCKz83y0j2JxM04jfYEy5bpRRkldVjWz7+J5
kTBsEi3yqr9nzE+a5Iism1Z8O+TKpAt7PLAvLvmHsRD8eEhJmDr7JqyBCK+h12a1ORPbT7LjfLNW
+35xRxDJ3S9meLT5P7w4HP8Z5rGV9G2GUpMs8Q/wQrUAUrgSkJzbFuGTNMoCt5VSTzBKP92xBrKt
6bVi00ZFOgUmJwohZvArnTZLtZ7YEwU8e0gBe5avDUdqjRExmdbMkynOzPnJB3EltJ3D0sZ0o+Hi
R1CQdubIff8FN4v2KJ+7SO8NrW1uI5PhGPa+/mGH+TwBrvvkNErYNnhVaR6lDpO4xLWGmzROqB0V
vri64VQj5AtDuKV7EDGAl7HiON2GKDGbnxHDH1hZVS0tfcAQ9rZdMkGtutijp207vVqUVd/lkDo+
yl/y64fQNx32RyYkPs3m9FqAhGVle1D+EQhueqsDmARXYChNIN8/VSPtsp0D1q/WBWX8+aT0erYP
VfIGhjfs32veb1Dog58U/svB5KOmTSgXatomY5A9VIvNifFM/x9R2/XgWGfzSiRg+RNRRmAY4GK0
Iid/PtAAioS9pJAr/5KCPkWq2qrzxzVULHEsD2gZe7rxON+AFQehniN3tnsGUlhiVP+pjbq4EqfN
S4Y+qOqYNUuAIydRDF2JROwGG9CCe9UUMyR2FezLzr35VXQY9JlHp+Yn1X7MXLXTALJb43UhLFOm
BDsTzfXIm2qL02TxilV8KTSHTg47VVnnya3lzQU+GBm4elkX7sTLKaxI6u0LUZhyqLFvJLajw0yg
MOa7eM9fHJjFe6ctogsQTuxYz/UqP9L8uod7A9GwiwtmUIAGu6soBJr6ikP0BLQsL6r/pGoapqp7
SA3CPdG2/33pYsbrzLIGNT0GCr9FKJFk/+IDgZZSbKkj8p4nodzdv8Mjgokl3qJgoCQXR/Wp/ytX
QTwFnkTRUPtMEAVCh/e9yDDnH4nfD63d5Pnk1Y7Nq00v22zlQIkKEIHxokKRQC0myTYDjz+yPriM
fOAUrnwSdmNG529LeLjlXC7YD19buBFPr/Vf4UMjU2D5+QdqpTEAM7l0Prxq+N+RKEI1WTf8qRob
eFTvKtkQdUnZcrc80VQL/a5l/NJ3e05rgT4B+ZxPJBItxdPN2uy8akKwKwkY8MynVubhIGtg3F04
HuIXyXzC0FwWzus/PCNuDJnr8YaPN67IsKVPsYm6COeohU+VLY00mTmRKrMiwDVxE0OglLXO2Ucd
UxR911336JdHujNgANPxsSMoigX+uNcUi4gLJOlZBFDVOp4hjQEYBsxPkHTcBlRmTBbYGXkvMw25
tQJY8k2CWDA1GJn9oV+C2DvcHUfmlSjFehnmcG8u/PYURgO4ADA3W0CbqaOC53ixpJjW+C0QsRep
tcwOLuho2fBB7yRkfO1Oee8pumbE47HExbBVyeILZeybx58doUyLeFz9AsjOpa3mdO7aWGPrRdwe
Sp1GhnMY6nn8zJW/sDkVrQhBsaoW8SPBg+L5gaZiposVNzQPpIU6KknSAIO3l0ztBJwmHpDh3/t/
zwQJ3sASWtc3WfiZnCvnC91fSI0WykA+sTn5PieWszZBaB5LpNZYriR8SCTFFqKf3CF4Pxot3/06
CS2hMb3VC8rkmIQRk7lmPBh6ethMFRARh7FWx+c8YwShevINNIjmqQRtIgt+Yezg2FCp/zYwr+tv
d4w9T8rOVLyS8vliEp/jgCy9IS7ZIOVZeuHgmjs0CbslJF44F1VLAPlHQnuzydHqDFSQTKPkuLG0
YqqlNUPm+deDKQGwYk2FS5FeNsTwDtzwW7b8w6eEedaCpJXzicXl3y8ogveas16F6gEGtgN7U51f
eFBsWq3/m1/ij1T/H0JVZ344Itc90u9I9exdTlqnsc4EPmnv2BMKbjK24miYB4z0KyR7dHE1/4lg
yDKouEnGkWkbyCTcASyDWnj2nVrFgv3lUzal3kej49qU6suv3GKJKcniMvGLsATrQiCLUm1rufj/
+6oTTqBYvpHk8u7zwerWzNhq/iyGcfvmP/fL+sriA4aj1QiXckhKEogH6SMBsZbRlv95c2aaThnE
X+alMHqgbrU0x318bqoRpfNMPjcOX8GPFdCqykgX8ctukBZltWBIBTfLSrMj4YabAyYKG3y4ac40
J1gX3HPVYe9qBe9R2q/djzhYHFQbLMYJLsyNHU0bPFtTNZZNRHLb83nc8V0OZixvQhSGlDxYK+9t
NJcMVAp+25VNH3EyQmXhFfYGHZULOnkf4avI9P1FCTnpoZLU1brm/HrwpMHBE+rilbuY2cql/nn4
H7gr7im70zaxOeFwWBMUa40YTCJ766BRlO2H1sPy3mOWo4nIPvIPsjhpiacsism0IVxhwijiVVQK
cXhxWPGF5tk1LmkN25xw4axgR4yXbwu7vWDP+1wAWOnoCffWfbTbzNnm1dQEGy63J2Ic9bu+tboe
GmSNC2LsaI4H/Te6CSBnF9aP58kdUPkRt7Ze2QugR23TN9dWxHSccVq04Jyc3K9G7HuuK27Yd+od
NiNHOCFgneUWUs7hM8pBe4oLf1QV+7qIdYQD5Xiqz0sYQ8TtedXodv+Kuy4GSEvq5pnYMD5DbNzZ
yUBDJ2j2w0Ay9YSdPeCQH+L3KJliPAZ7IHXouXjiXZPtX20ECyLg9n8etXH+FcVu0xbQH1ShYQm/
55vpQG8kgibMcx1K9yXMG1W9zS9js/kNahAxQ7NW4TissLCAB1c7xdGAHzhSbZGLASRos8L2DHRz
zUYazopx8IQ2WC8oIPVAkQK+Nt0XINftlP7kYyZhaFlYgtHQvSzuf6SJd0Srvj8pC8Yzrzhloa7S
gVokq+/Ag32+HCYBfZXpkYAb24o+YT+ZgUVBuG0dN/YV8qK8VNpT4tPVd6ae+yNm0Hf3LWt93NWO
3DwWxHOcdP3GE27MoXumL4/fgn/KQOuDmXGtIwUr1uoakSExv0uKL2CXnuekv/UE1PdvhbcPl221
33/TXlTpWkYlXRb7/XJR6QrkFxHCbcrFVj4pOce7rmw1yGVw0pYS6uioOqbyjyZZQD5x81oP9oqT
7CX+/hxte0gbaQghURqaxW1kpjWP8856PoRZ5VQjKqRSRWA3Ha5DxPKFzvn3YrWGf8DXKIsZj8TC
ZVWmFxnG9Jz8Fj16KHASrd8CB+jTsU1gLs7+A7a63VMC2tkeusbCdOXykKttetpiATXz93cPhHW9
u81eWrT8bXlEVL+W3Q0C2WpIY/5QMm1oBwrlQnXlywkxjfI4Y5ajqTEO1+m+ke2dOvIJidU5iVdp
6f8MlUTS8djQHs6+M1j6J626BZRxvbz2Gjw++lJYxw4rPF/urNdi2aU7c8sZ3B0NaLRW0JpOezJq
CwIIaXdDHGi7MNh5juicWul4/2/h50AdCr86yMWa4HND6drCqqP6Zc6Q0Vrd2cPAQ66EG56Nm6xL
LC1hrrxHPU45XUCZT3szvU57L7oEtq6f/eazhJ6YJWm9sAXUkS8JbpXI1k9mk6VYdMvK73+ApSBv
gLXWwKTOKzWHSCFfrb9MeJXAIOMirIrtIG+lr8lR/ruwBCDkU26nzp1XjzmcIb8Cx2T5bXIMAfK5
E4sIRyhZ719e1pEF5RBUlA3FNiEenMcrfRWy/4Ux9vHsoXDImXY3Ge0i5VqxYZIwi2E9cppWHEH7
Mchc77jnXXxuL1VbnJp4nmJMFJqlpKUv4J/x4gg8Obf4YsgMT5wpAY7TuVVl+1W9IfEYruaJWwZg
OtExGaf6DLJbg0W2daMCR5NPcy6xN2Bg54tuhxevgLRz1YKDt4TlhJlgMLRaqR9R8QUAe1igSpVo
YR7SGipGY719PD68k9Ue3liN07K2n8YL7eJG8NJzUHfEoi7kpCS6eTaxklb95nbZz+veudwDz6p/
NwiqyDFyu+wL6pDp4LZShvbnF6HZJO1agU8YX48m8tJJPKBuhnj8ZLluaZmDRj3v0rr8umNKtOM9
OEeoT6t1NpfHM7NFufJE0dcVl3PpYUFwAP71S/kEhHRKiqF7RIdC4Y4H4XqmUsZAPO0oIYE6CskL
xsqBv4Y9tkNWhcJWwOBC2/m5Qw0vwVHY+4VMYLssVMqsfpf25e2zZs8t1Ft0eHkfkTUgXHvPErk2
vNSg4xQ/ikaw8k8CoE0dUPqDtyb2t79qh8s/XzXM1h6mX9dZOlMpvJ4d61kXUFezNww+euYPCYBW
nZ3PUFk5peOn1c1bHGAPdOeyWNekVdojkFkdUVDPJU+/TGJiBzsYawJ6KslS1iPe/zUxrraiNFbf
gLfzU1sOWB9zcOziED9kixyPEglb11DfiFBGu4djv4+5G4T6LAMQr1PHeHlnitj+Rzgfut7pYSfc
oOqNdyrLpCkT8yefyZ6LgfGL/qrdrPDVEla5zom25gxqSfcNq5nZh/HfAMQ1WMAse66KiuzmtBt1
3n2ce8YiPFFrcX9E+9+M3siny5Dn4uIE3H5z4glcy/eEmzPDH40G+RxVsX36zc5289D2rBQDU0df
hgA/kwT0r4kF74U1SR3R7a3dl5v+QPUxKppV8QJxUS1+efQsOWd9zpKgOi7dCa/X13N5NTxtjF7Y
G+pWcoarWt4lo+QTN7KmtCqd1fUDUZjKT1rOs/fN6CUud6TazRqPV3NX0hDFu5ZcAOhp6X+QEHxt
Rypkwc2ene/DQpDXw+iz3zdSR+/V5GslF0aNc6PEM25mwf3kzdm08i1R9Ix+ts5qNfiFxzDG7xxD
Wk94GXQc+XmUgkMlR/C9odosdDMBtZkgODk+xvKK7j892mHtLoZRdg1895SZJM4Qq78PLQ/CBQbD
S8N/fNObZ3sDjWLx6dq49S8bJ6j375JXulHgB0guSWeUr//Q8gE0jtH/cCxTMDi1maVC6ILIqGAO
2M7nYvKnXCJEi9zzt8tOqPMD1cUSo1BSROlpIjvucqLw+u1kBnixyJ5i3MUUioe3hK2JKR/rtmtq
hVp+KSgp0qFH4DxgXXBOIQFZ9sF9MyfBF4HX4PjwP0ib7+J2B3UASnaBZpyoMZANZFAfCx6UNsNd
45tqHF8+AHsAsDaO0P/8lEb67M0Tm1k77gI5P2lI8PO2i9f3QzAD1cLi/XBhgsjCeMweHf075hNU
9wQv1Ah3HAuJjhoaIa9KasGdc0TUmdgEXxPHesd0U4LZxMHiuZzqCgyeCgdnugfPdmCfEIRvjLXP
7vld3gsB2RHV8jafuNDla6c/o4Yoxu4vg5NWKqzc7WFSxOc2Chv/TAJTaoujlwXkjKT+VnOheqGi
3cw/dXVnXVvw8moKY/oFMm1uPOnJd+CBiRZ5PnhJ3066xlalMn//BVxFnK0O2eSU0QxEJnoXTzxT
UBTPQ67Dim4hF9QlI6m0VBpFi/c8BSqugmtF3ErzU2a+XcvkGuczXduq7FqhKWzSFk66zm7y9M/i
tkrL20mjlXy0nH4onFZy32/iNyxNXEBzz7mw4/6kZ6EYPVyCWPpCJmrXsMmzsZOHSKXaz6u77lF/
MGgY+ESel+oCvAsP7hgGhuSolOTLG8QFickUmszk2XXSWvhE8I/g594Df+avByorzB3byDLZEfz/
OGzHGUkWnBRiqhaXz5NFmdPb7dYvtO/OLI02GAGWQJZTXdo6JCTcRGHcV4GFxp5W5u9FI+O26g6v
UU3hfybB1oer4QDhm02W8rrmWleBX+4PiCk/DK/YjIEBfpf/QoPK5mNePCjgPJApmM7n6g7zL42h
c98vx4tRgeRM+y0oZ6PElEnSS7EgIrFuKH9hPqNUd/gt2/KKkerJzsGtatYZsRXG5ZKaewMDcpIQ
bzK+UvNP8YVedjTUIhMLsug0W3RPzbyCnTldkRkuiQHsxGccPEXw8CyTYPREjkg6nIqDgyAb50UL
zk4SW/Nl7TZatH6i8V4vtFetEID3azbp/EbNrWy3GWnE6VD5wvL2dpJCDA5QREYpGuCEgvj8N0K3
SoofMJk7a5S4BDJEkzi55iE+V9jrlLNNlrfRWmKCVT9R1aKPy1DWz0UDGlwn/WIz5/VTwMOoRAac
UHaTSnc9UpnQT3T7pCCrkEp4ycbpLokJoOi98gIIF26Y5BAu4uZ1AHyqhdU9rvspYjen2Cq9smS9
QcJwInUXDDABF7Rs5nmKtVo08OUrI+yknPv0vyfYyxPEkIPCw/9gbgyfmGacqhxcUoi5Jfme+K4n
bV5nPEqeHP22y+kMi+NLxq6kiEqWGnzohgGuHVKcfBrl9KUXGTUYEhqt5Ughe44ngflFO6RuhUR1
PkKRNiWF5qkvkYgQKNLAC9ZprxU0EsX/qMCYVZ2ExJi97RiSM9ugjC32LjImtP+YrKAbK9sH7gqF
17TObmQBGWeaPcdzx4czudpWwFE5asl8Dc8EWpbohRhdfFjisAxVnZWMXrfV7ylKUR0uA16GKex2
wcKmrKYL40Yx/filOjtxalMAt/+LYveUnNvUzQjprvdZxhmpkqrELBYcnUobe6i0E70g6A/4qjH9
cIt2T2EjtHpeuGXoR/A4laKklRLdOvT6dX8Ce9M0ElMX/LyE8r1SB5egxtRmKI2zWSzBvFLCwkVL
SNbtQO/sE7/yN6mWfhOQh4cZy+/wcGdWNbJ8/9onOkd1UqMc/dib96HFs4zztCg3Pzmp/2Z4qfrj
wOVxdDpDiWunTde9wdXQn/jCFAU/o79nFXaFwUiD7AC2MNRh507rTF6vKxQvMye4ftiRAuBTaNWm
rr5euSi53/7HDDELB1dp9JIwxwuaLjsV3dB42baEuCrj2Ozv5p906OtnJgj4PhBg/KyKMb6KEIRk
CbhIioe8KaIFUC1ENN9KkkP7F9EeScjzzuHKwv25Y4nFkVqOtn633YRf1qWXaUnF5k15SThgckzf
KLZhbey4O0g6W+YXMBobWh0K0opw3mbOXQFJKWxWtfvr34dlBaJ9xhVX6ExU1cc7C5fVffdmAdcp
xstRejZi+re6nGxIWA7VH7lGqNOlr+4Xk7iqnAKkH39iXqwGMFygUorOCIrb0unvgy5Q3qvQfbq9
nRatdviIXfeZlvRtfwvdkqfq1qbgi1IFPQR6PoZ6oVQZqX2wb2hR5mBxvVoGGBo6ezV9wf6ZJfd6
bSheGkx85ZUbELnt09n1XUXknSVWtrc58R/MIFkyOITVT/ukSCs8RumhUhRIfH+Jpi2yrUaVFM9y
vpy/lfKTrxjTVX/yaP2GPr3w26WMq2lcVVZU7n6tFOX/70UfQXAz/fPqdI/lpWZRTDqi1654cCDD
VJr19ohTY+HE7bRj41qjTle3As1/koFID8576aYgEstpahO9UZm5zNUS5JXs7hkt4Wr3oqUbOIAD
izMnv4yvoWQ298kZpbk8bUS4MkyKOuNeJrpfJy0uaKLEjqyhx2skiF25raqCqv/74FZLHNTJugcB
aJEhtspg/LvqhSS5qNQsV6rG21eBh81GhHFkJ2ASCVTNE4R4qloGHf+pXY6e4XzlVY6wF3w9ZEGz
7JsOeS3SQKSaXnZWBCC0vqGwCbpl8S3TvlTMrEbmViXHM8B5yC1qil39jecOO1ucJ8m3jz4Byzu5
RXrLi9ZChTDQLTli8zAClTVCgY76EFfAItGsuig+zPipVh5YpwJtR0mN4wMdBbGuMuYEhrrxAxe9
lpzYu7HDHxhYsTzwPbmvdbH/EbiFQGjea+wK6xo0X+QutZbDCLAkBU41pjBDObS3Wjhu3FEtaQbw
GVWAyKjTsT6gJCc4NiDag9dr8BkL15f6Y5Kb0Ew9CUOMi8eA9MujBOj31wl9zHnN+yuEV0qdyJs8
1LdoaJ529+jqteZx9AbVZa3NlL5IoHSIhBcyo2uebLgeYTaIyrY1iVoKtWSGDwuCqH2VML76HF7M
cZi1wMBQBCg3Gm1tS+avewP3Kjg+ks8DeFpFHrmA5hVfJJ624yJkVAGImu9NbKOTxFSw5W5GN1Lw
6IbMwIfrWl6XVsIy1H4igkzsBjrbH8eQ8ThITcDJPJTTyFEZQK5vY0uxF/S7Frtyapr8QRP+Ufo9
ky5ZaATw2rqYbnfiCXi4KJhOW8wSG3M7F62UhdcQnP4JvhAfZmvm4VoGlGH4XF5SdmNBZCrB659V
3JcND+jimSs7bM5R8Nzo3tBvSOp2pl5sU78vG/Wmnd4JsWGnUMwMyjNmrf/QGgprjmoAR2D8zmOG
ASkAXIaiCn9GJIeLhWqzMQ5nOk86N0ek7guvzE3+TKK7VKt6X6OlXfjssSrlVXw5Z8CNnNilV8US
PTm/+/GWsBkjDWKkTGVi8HXeLx07WXNeim0KMgdvFUQ+sb7QUEM8hMgkAM7N29VLiHGWJQCQngm7
lx2S/Moq8jd9jG5MATzxVmCc/RmXac2S9/7gpEHoADBX3xYQnmWIn1UcEaJ9SD4wvtayg/g+d+eO
1TRRHkW3i/cYBMkLqoSQj1CNtu5bsGwkwbpvmJ2H4/2r3e8FyHE6cKvOIEgRNpvquKGdmziuz0Jd
e2Md12bPgx4q23Umxf8dh9rJG/Dyjp4NrJSRjDAHswlEiI4CLuBrS1uQrvRWOq2YjDQ0Bf5I/0lO
xLveow944cuQugbi2/fXvU+Ds5swTkAFhLqZUEWBRvMSXJb/Nda/cdSvPpNUyl/dfGojLn1ZqKkx
CrP0LK9n5IEkMhnzevnRMNFeUl05fjPaEV7q5mNd7LasNWrSknfTu5AFqz0NwoYHcGNhCXGlEVl9
s6IOtbUzaAZzPXKfrlbmPD25k45yEPDVeDl6TxJ/0Sbc5NDxs8NQK2fd9lVjPsJaHWULZr6Xgyaq
4Vd9RGXv4kUfCbQpm5hQcEMNlMIQq1DbcJW2twFfCKG7Fzov7voQsCawHcfo3VroVVi72LFgwrCH
/sOrMdTU06iz4F3oqmfU07yPa8wuReeoVU8E5MKDJDBhtfkqETGFAwaCdNluMpTpxVEAypILyN5y
qurUZwSId1kIiIZ3rj5z5YgBGdkSbkdzhNttM+5Ug7CW/mxfeysWBOF+GRSarqiRJZ7wuWkM/BKc
796LuCfihptjzhEULRyMY6pJu0SaSXo5+5+QCtkETMoo42NZt0gllpQsnYvb95sW91FA+Hk3xRQD
Bq23ePPKbyepSwgIqTvXC4JMhKFH8Cpbp4vhcnx+FW84Lpdk2GlFAK8pfdvQ5+aNI81udrZGa2MM
h4wavGaglSXe1+xACYXVEf5Rdlqgr6a7g6yTd17ZZfUCAscK8cTtS7cDAxMR8wBc2op0jTiTLSVx
5OCqqKTBNuQQPdDetry+wkB/q/9O4D20czTa5W/2+Pi/Kf8NYhb+Ujs78bRq+eAU4R0xffjaxEVt
A/OTq8PVokf0t7U2NvxQ9okLud44r6R2Swr7axEiy5GJHmrAQXjQTU5SORnzrLLiH6FMBoglFPvh
oyqG2kH90dm8h/m5uUfVFvtpyKmzVkdrI0qTE7AQgvEH0ivImmW9adEJmpHa2syMTzzxuyNwm+fu
cxJ6M5OaZbCfPoAvus7FgeLr5QYcKx9VXVzPLDOzZVp700VXPFNUQDUo/KMHnZceckMUbx78Ucue
Xi3wK90fFitEQuosOFCIrnADVooOeuKABbYjy2pauMJ9Nw+1PFjsL1PDA9alx/1PKVYt7dQgbZFm
XcpLBUsCu9zumaP/sC1xjeuUCSAKHulzCky8gUiuhSPeNrC0FQ9z1Q/+QFPZvJqfulnzvMFr5QUX
pX+zxJ06f/HfVERo6rgOV2e1hbGWOSlJIRmEJCTM1S2Bi49aATPDYRSCxQwIE0Yd5T40iqOc0xg9
j2SqOF+n3UuO1Lj5U62+HsAgXJ2tlnHsltJfwfAc2rhWesMPoFebRKSmhqTI0MT34YiQuOqwnwx8
moF9pYIDZ1JMzZaJAufKgqW/gpFuIs6vVhzYzk4ZDgAkH0Y4mQCPcXeYGfFHkWe0wSEiMbBt5S9i
LAeE1mp3Soehh3RTjTWS/72dlnB4Q6uMIfzFOJlASrzJNRv8NXsQaMDQY9Fp/0pM9BxTIPT5hQ0T
fuH7t7nKI4W6Zd9dJ/46CB8ePVOTSP+9ZRablfg/fIl9KEelYoLi4i/b/Fpy2WjaoEC6hGFrG254
+zcbs0PtJ+vqq5VxE/YgccquwGkG1LkhFneS6U47uZNT/riRFNB9ygwtyrPWc0nTaan9j6ij2qin
h1YLvCdo6fjHS4Lntj0PO6ZfWtZyUKeVSTzeOlYWHE2TnedMgnMxMSeJeXmP1QP9SQrCZ+Sh2q2d
njQHpQXR2NGQA5fRGOnXN7K1tpcAB+9jtFxpm26LZRVNsSD3WLjtvSJTRNBNNAL+KRPdq741TjbL
6G92IGXuzoBQ4G7PKqEE4fxNzX2VycYXte9KP7PiCoRAmSvi2wqEwEQ6plU2y9XqUY8F6c9Yoivl
uApIVVmy7rtv4HsiR9ND54CxdUjsu3XfOfHrZKEEdPp4W/xKq326g8Ygzc+c+hKnhY8A1peLYobb
wrDN+v3d7NaLHYmqdbDyr0oFci8siUTEWFo1gyN7s++ZFV72BRsnx8i0K1VqVT9taT1MupO3pr7k
UxL0uluKkuLNRcvyl4xm7BB9U95tfKGco1/Pfd7M5bjAAXa5m84J7K5ORGucSFHPpHaiInvx66+8
XgvnOPyPPBnb/cottIa3utflGANwYJOCZvVX3bbuCPsUAcwzwHEeWFFXVyudrE/twgB/aSqabP3A
kEaNy/Oku8YzG23RJiCNwB/cs8lUUPUqAj8fkxmOZ7SukcRWFuG7fum38zdn2m/igNI48W5UnvOt
zVtsq71GYz+GducVymvWsdi+F7w+XjrQRUXzRN5jgifYyWD7Mc6pO4MHvQmZ4f5nOhVHOaYykGJj
bAwR497uE1EPoDO5LOFARQGN4JX8gIP6yQoOm4WjC5NBs8IbdpgIPtr7mHDHHkzv/bU05CuRVgkB
kqmdxAbeg9zOqIRl3l2hHJaHyYg0c1P3joRxUbQMrLkPgLJy6g2TJrNMEyFhkJjYO5LPA1/DjVEc
jc4WBgBbMD6AV58lxmWFRvQu6bjDt8JFJ/Mc62vazgcUeWgnxOB4Vc1J5ql9BkLojYzAdWRImktf
yqxCeoGGPgZvqE0FyBHlTbN7ZRa/yw2yk2HtApzYoyQKe2rpuaUr+aqA4WErLBxjHjGEjh/HMrXL
HmU1PyEs3wJ0KwuGYrM+qG1gD53jo56H4qMBJ2KGePVnjBF6bw9S0USACBt7vzLtoRLihFuvvd3i
kQ3v+Oiop1xVXFiVB2rUbQeqXfUjdiY2uHgoHK4prDO870ryQ4Bo8RmTZMeiqYxrPEZFY5Te+hbO
UcUpQ1qt/XrDH8kMhbTPre/wE0Y1pRwIPYnIZPimWkuKr9Y5o1iBIziE0rhRIJSKi+N+PlD0MQq0
KFBKOpgT5PzGMRzNIvPBgea2l9kEyLMKXiZK4334yq08gEpd6Smxf0zMmUPwGA0UwxDfMH5sxLJe
kj6jmwrXDf4NHw7fMtPyvvtIbfTm0/sX8WRcnXoaIwdtDAWKE5TbdpJ7TxpolYFW+da1WbQyH1FH
9iFON/uB4SSxA/z35yDgMJvjIn9l7yNRu9ntf9eW01P3hvrPLTwBse3snWMFi6Gf+ZCpq7VHVvKS
rk/8902k5ESZS3EysRB2EG8/55ia2r+E3nGXcrISG7HeW2HcAQAdqn9GSpxRFiZ4VcxVbeyiDRdw
5NhBkW3QfeTbacL+42HS8MNKg8t+HbSqIDNrYpQkw0U3zARyuZYQn/GNzuLZjM0HfX0SVeg84YWX
XB2zH+M8DNHGzqrt1ek3OlodDrp1DvrXiXutlz5KdCTRfzEhbSpCytv9hksAGhebujt89wQ19nrv
tLvBwy6s1zogjGtQSKsd1uMUDbqY6Kki7i7b6Myq3G/IWDNyG1+B5sdRgfQfKTjD+W6CgyTw+H5j
0I5cJlmBI851SRvejKWlAHxBEpIZoJHFc7lN56hH90ehamUnehcX8Jniwhr1rLOSNm+QtVvK8Q1K
Lv7BOGqW4trDb7bcI1cdXfmbT656rhAHOZOfWaostaEdGqX7nOp9F/39ZadWr8iDCUZuh6saULBe
9Q0umXxD5Yi4g5f0bzdxs1uQrIc+kBHWpGF3CeJsG0WPzHSaBziNk/6zGXLHEtGAj8zmHPnx84JH
Yp+5CnwGPaJCRK7Hd2QkO/apI2oNVPJqqgYDOK1vaV9aDRwPtS60qbGB7zCGQXiuRkdiKVbiTsQ5
2l9afHnD31VPJ/IhZy2rOk+oCJk62C3EX2pWvLfODdm327jTR9bqwDE92Fh3JhzHi6u4yfCRPQWO
5TKOL0wxZMm1gfmiRMO0PcWeCU0Yrqbk84keZ1XjgIOkJSBUXHKsuC2bJe9gBNJgMxcWQhGrEsRL
XxxM3D1vNH2VnM+gjAwed9OqW5OGoThvke5ZvrG210tdjU1IW90clycm2Tmn5NVjAE9T8qNdcZYO
RP+K43EHI0Cs5dP/UbmJEV14EatvRCsGalHG9aWeByBGTiII/nbWNZ2Y35GnpasZpHjWtN8j/5/j
df59NAXUH1tu9MuDbn3jNtVmzE2oRbwRO27BBEsoDHG8BqnAt7Al5ye4mNZ0QCi6f+Adx8BiyPuz
l3stc3ipwBUOoCAdwVyTogFqsZktKucN7CxCDyLjCeqCIdXbCEN3wRoang/KXg4eK/odcgHio5VG
DmTP8wL90gw2qym9+NW0QZCW7AlBLX/O+9y6kyVpDKE66VXK/imRz81NqMpl2kCTAo4MzDgdUej6
bcd7ducijSnfa2gribwe71P3Awx7y7EXr+Ij2gjlrk9d5r04eEI+6MJnBXV6kjKLt9PgM6N0p+lx
gxgS5Qp0x0AWnq3UabmvfsJqi4kW8g79wl/poXXjgF1mWEfdZXD+wx1iUZJ23feQiatyaA5KqPNH
KUH9LM0TeuigsY+iaEaltEyDeOH8odKgQdppfaWnVNYg4ste6yaj93sklyDcBJsbTWourfSpLyU6
kNgGHyeXFaNyREsu9rL8HOL0GFFdF8SYwdEL1dFWOpCBsWluzBkHD0LKjOVv4MGoyXbz65RmASoj
6Z7Q+8F7ykNF8bneN8c7MXqG+oZAb6jzPH310Z1xer417pbQ4v9c8EvdFnV7bnGlLYy5m/6dXHpA
nY8Tl5ZxJTM9pI2Fn+XEwQsMCdcTZn22z0h4rcUCKP9tijHboEMcwLOJIKUZKTl2WV14yBsy2y+5
xj2iIv8gZgm3msVJHEle4mc35Zn/YdSZgTOQQ1ZyxmD3w6RBkVCzfJDWT3I/svSlgMEplN39xfDo
oB23hu0vwKY3fASk/fBGYFU1Mr7vQzpX+2/VVNp5J+o4M7fSo8tWIzCidF8sTQQgimGPd0ygweMp
XkzTA840rOfD3yGM34R79KLW7RL4CjtwYMbypEg5bvOSYfRzDzdCaXGTFcICfFLQojDlEr2u8Dg7
W1V4zCzFVQnjNBSPcEUq6BKW1mYDPKqYxAwqKNXK8tC3KPVJYNgNli759msQGfvrY7KNqDf26wKJ
eLKS2s5SafVQW+e7oFuhdhdYthbi9yxQ1XxuU0mkYsGMi/lNUVCsEBM87pZWyQSxxmncI7RdMRox
riCbt6+PaIJy/2r566ZuZqbtN3uv9xA/uvxJu+TrEgsY/DyZbWLjloinSpqhI4Uy2dwB/3AlCHg5
oMo7w7cgEJVDQVBv3vg7l10YTHb34o+Dag1Dtxn+GpgqnUIgLNipgaWQzKaBslG4NVfZk4SYIgGo
ED6PpVXSx1dXJW0/GePgSqgXiqF2Q8Q6dweC8GaZisyFcg9TFDpCUcRIY8iJzbomQ+5dRdAtoJIc
ok+Qlrur97ej2CFYAJLuI78wnMzuo0VxBX83cMQ6FkxqCNvBOf2fCbaNXUzc9qqv036mJf6gC41w
sbIu/pM/1MdmyN5JbQmnpOgWG9JrXbswnmyJIN86rJTOXEpevi3ne4iST33y/AAZp6fAkxcbDkrf
5EVI49ylfsUP61CIW/wtmgtVis717qICm7lYpQ1CevK2y/cTZUBzekcryEkOR8L3gOV7LoQtaDnl
tnIRDnPK2Q8tyS+sRfgvy7MQkQJgW8KmLU1yHu+GLa0SHl+J1RBw0rBSD0b2bcmTGASE6xCptdrR
ZSgK8/QEvn+cVV86idJRFEdE7MU+IKvUXI/uaF3YN+9/X2zitifQYLvEJqyP9FlXBgFDkMPPlsLK
ex6o2JFfFQht3LBWi6u3o2ir7GqrHL00g2rt7JJOu4a+Hgj3a9BD0PyJ5hOcobvdvp4wawcc3imC
vFdKDGSxzKhqwfWrSkMLX4zRqtygkWhr0F8awD6ceql+KZrN7TQsVWvB+b9nhlSN8gFz0JJdSlMf
A9Ohb3uj0obbz8/BV32hZch1GmTrGA8jyN4e7+6V3YuGc315BGGfU6EgAIPb1X7iMJjbVh9zmsQd
L7n+YBgLolh818xUK+YCrwHz+WT/0ASD55r9TBWEqO2WETwvK9/VGphGAqNovtP7M/5VTw322Mrp
bFdbku/7V3ggVErdGAyfASNCXaghpsnMY+A/3RSWV81fQYvsq+i7ASlJBm8sCOfVx8T7W2biF+DF
wNQ6yLVQ8JYD0f7Qxx1jyty1iPys+kcWOV+LNM4sCg2KomYnJHs68xX1P9WeWrvfJUeLL0DPUbcK
kzy7QkgmwXmvn8fHD11yJvm9uIdzBrIDjrzCfNzvfsfKyi/NiFDciA8mFGSgUoKP9KmA6sjz/05T
rXKP2Z0G/SUYiMEHutyYuzPnmU4guGjkp4I7tDelnH9yyI9DbjaUCuUvvg/pEnjhN5ZaNe+g1HEN
tXu2DpR2UTZ4c4fHLjLmVwVhT8kh3w47xp+S8z3XsrGVsIz6g8JqvcWXngSBWPdYBNNYe/k4wUX+
gGpidvr6h1dK1puDHzY5oN5x6C5YsYQsOFZtShPSn455ktoapp79HgznD95inqTIT6RxXKIf7g5t
Q2HyV9dToGpxKNO9DpdKpRouOHSTAWdlaReFKUjC/8Nh3DnN/mOgfQGGYKqEe0H+jdXNUSE+bl10
QSP+H9cAZOQLscsIPJ1OL0aRV4ozhR9KrNrS1uPBywr1Qe3z3CWYXkgjj3igpxtUVvHN8qkQPfIx
mGn0Rt1OBCj488hE9YPCIudsYDJKvVLak5gFifIkKcnThAUFE60OtPLpRNEPeuT84UKN3nHn7Z6X
wJdlCockZNjp7FWFkPppcpXWx9daQnrR4WXbox1CBUH34TaE9GpoB+XAag/pnhsCUHj/n8R+0Po+
CPCEOUEWRo5vjgDtKembdVTKcQUNAu3mwLQyC82cLCwxKs7sciBz6+vg3vWIn14TM8R4NNNApSN2
hMV9YNvBl1n0zW13+PxXyk/o9TMbKoWJzisJsq41xP9dug+O6YLx1SZ9j0xzRmi3AZx1/heCSD5L
Zsgc65iJFRVmMvjHG/3UwaW79R8/dJiY4wsP5UxQQ13XpcCxVLw7ceVyeIZJGC7Fn+ubPjmQvMYx
mnGv5AWFz+1CFEgO1cFLX1wnKwtSFx2pKEDHbGulgJ3djIdAv/U6jME+GkWt3DuuPMsPbWiN7o/7
th7ZiyHYXFCTwqFSh9h2dhn0nfIKXc2JNX3Dhls/ypOjJXRAnuKVNABtvj+BmFVGqZxFyVqSaYcU
kvdDqjFa9zF8lk0zWUD22Q/zJ+DUKgaiG3EmcodDpISU6qOwPGM/0dIY5AM12DX/+hIH8rGB1QeE
Q3Mt1sAK3f6ocp8lhFOmKbk1HLKb20VHIYuqNChHeU++0Kj6UrvSNn6Q2WnXMS1W50ycqdEXFDrt
ZH+vqEvLTvMt3nRMpY5gg7MVGODgkkRUARGLLiqZ+FYhMV/ARxJTXg0FrAzPRh0OKw2JoQHqYIZZ
rZ71WFi3iCm7rQ18/Bugmz5TfNObx6ySP9vNQ2e5VUfaWWykLByNd2YpB2AvO+SMASCjK5BN8FfW
cQNhjgWApna+mEs5HeaebmmPvihRUbE5F2hgPxQghbTZkv24weaNsmNRtWk6K/CWG2VWHtV3kFKL
Eru829dZ+mGfcIhDf6oC272Hg6MwFkPxM3Zayz+v8vbN8vW+lrPrHB4OUFHaeuEIDL8W9Yud/Acp
shId3BodzgeNlPG/JGusKS7vs2Gw0T1lsoM+NRP/hN7/VEdpz0S3fc54isQdMXf9YOSzLk1DZg+7
qNFHQ2PP6yq93bdWqphoxaiGIsrQzszukTMk/zDS62i2+1YF3+6+mlrHnEIlFyJX1dzd5Lvkoosk
sTCNRd1iqBf3QUTptPPukwAOiGB6pOCygnxhbg/9+sXYamNNZvOwVHnCOAQa7bpes8OLOQtPSmq1
m2z5mfM1/trGTzPVTZeY6m7PVltXjlbReePSozFVmfLBapCR3KsKXuJZATL9XwG+bQKNzLq/b46U
SfCI1gb0+UUKerPaaG+mUhIHofy7FaNzpmHfrmYp5v/kyjyM1uUFzgZOxRCgs4Qp6CS+zKVCdZvJ
GYcNlL1c1padbFKFMzLwWB4MG/Y7C13kz6pDgLmo/yxuKvoPTXmuj6JhKXuH2z/RiuxtesL1OfXk
y3W1bPGET/KqM7Y4x6Kw/80tKTTbhzwhaTMjFmYfUZW2WjVCbGtP5trHmAaYEM+GX4GgNJVhL0T0
P54lvKFHictsrxpCFnU9M4XRlRz4c6ruNiDGUwwBcQL2uc1T4GwOytm0sRwxjD3nIKGesKJgK2IU
x0BPU2WwICW/vhkKOfM8WqQcJPCZlbpWR7To/+mHKX2DcM3m+cMgDb47150XNwHuCmMlKYGBd/EF
mJX8T+n+9wMl/+CuF9gOxl/6nnoZMTTXEFKw8gE/YCD9vZtjdafu3bhbyB2rpBzaNPDb9OkssYaN
49C616f7OmSarF9oFNphbkS2G+MXo1+5oI7fSoTYcErvAoZpFu+DK9ONL1HrS3oHjRRBFWjMonoI
FRL/OSNvWa5cYD+r2r3QNqlxifwb988HDj8qtAym5YSmku0FMGGly0jaGzPn9u2kBJH/uFGugRqk
hW4OGRZNzzSHdaMvS0+Xfe2DVC+IsDbKDLpjdHxrgGJwy4B9BqKyIV5oH842e6m2hu8RQ2K+znMl
Z36PYk74qv9WINiuunt0esIJ1EefSBfTJqZbll9+58NHdRKzVZvCtjkpX05wv3u4wNRw9i3rO+Zn
UCbyk8kG2QRBfVRA76t7/o/e9mVxqXG5fGqQHbRsGsm3LnoHY37tSxi9TmdANMh4+6vpgONwnWWg
KpCyVTpvYV7OBarEfaMI5EIaEp7kyWT7gTAZKFXIU2KBLz4kK1s50t3lyoQJSzYdnHcG/tBOTiIX
2Eu0exmy21LCltYjBOHpWnxA4rvJDcy3xbk/qNaZ4Ms+18LIiAqYSeOnYjN100N7VNPZ0OLY/G9n
FH9s4qhouoYW6wg/HlLeW+DdPmxtVP4e4ob/GlEfbuaMsV6Pcsu0mCK9ocyIctDfCgoWpUn6hVcG
GVWglt4yDVIY8ZehaqHyEW5CNcZ1GsBJ/MDyyzwv31MVxQYLl1ten1DwtMNGVG4bNeR09doCL9BA
cduxVZKi7OCSI89QqILruMtR3JRczrlviyNMBr/5xuf/cVZ+jiwSPDEzJcG/UHtI5UZ4lOXFQbSw
4UpEa36qDHIiHYjxuZxihZ/O3fJa+nFK2PWZiv75qPbcUqkY64CQqkv8EEooZcIgmGbHw24N+j2X
buXl4Bgi679J8Gu7az07MNe1/I9Z/p/bo3x29aiFKXzjNHD/z5qaQeEQE18Mvt4iuW5jQVtpUN0C
xrHkFy5zMohhpy+tylqQ1n6KpopLAxdImtoDVMApkeFEcC+78Y3E2KCqkiPDOAOqJ3VvIqffqwM8
ZsMNOmTVlrjhuiuRZF/+alyOhZ7gkl2LEgq8ubSTIA2VMVWl3wJ+XPmdweQTanH7TEq5O5hWuzeP
T2xEMcM28ksuvgrofo5Bv/Kow922wppVgo/rHhNIcn/PXO1Evzw4AveD9vg5pby8fSiRKukeevmt
plOlCTLnXEOmS0FIx8lgCvPTAI+APVDQRb3gwzCq8DJLrfWr07wmZwU2PVIu24yu4a3/vKnOR/fb
eEJTxE5axy6We0u701g8MeWVjQH84DICgV5sCeDcugtHSumv20iPZx6F5Ymfw8hzVz0au9gIKs+p
tlD9xAdWLF3YieV2Nzbgg6eugADWKmHT9Hy66raa4JBqTLRwhSEiNlgjwatsYKFIG/yeTak4zSb3
OUwEfYodswC2v2bahDFczAMxObHuCE6iuWuRL3MawmToiGKaUiMjHqS1Zk9dZRuqVnBpEUbr06Su
A6lkfwyOCi5+vc3okc7g+kS18XzE1j0MQnSAvfXq+4aK8qg+2q8HX2ElpcWZpEcCrzjrj3NTEFWI
hej5N506GTCx0v2HhgyC+U0glr4ERZxqr5OiSW+rqGqcGdCBMDaMa1hTicQo68g69jpQFmpJUt1a
MKcZuDllvFstedVTDhrqZLJe8iB+7mBEeLL4XL4hfiFzcKZJ9fNRzY3CkN8JokXER/F3BDFQQlZe
VegX2tgBzdUoUSvEPf3zCVXrjhJkQ5jyyoudlb6VAAehEtCIZcoNgJvBHivP53EOgZMv753UkUNH
NsfED8gATkqwIbmiihQsXPWzlizZgjmxFLgxCJjX9gt2HpCHumWh/P2XYBDyVCnaSj5QTgL2CW2D
t+LwOBGmAtVX7KWkpqjfyG4LUUecWriXux+YLyFpiuaZAlJHHPNEFCqBzCYF87Ivbc/WSNRlcP7P
64RSoij4uWAHsf8iQZxdDxgqiZcUlV60Hitl1rwft6NzJpI+mL7DMT7X/zatkzq0rtTFfq7RXO5T
Tpitu0B+LSXL+Qz/C/Vg1kDmjKHTu2L/lp6caJssL/ewC9JqLo/qAHxm6iA1QOhJhkR+poZuLDih
1SjCGQpDKRyn4VX9Ek1C4sIDp9CkJ3YC4R9/XmV7HI/mnU84VFva3Y/K5HAJUs5MEpszbvvPijEd
RCZ6jodkfrja9yfRgDkgkwo1JBMEhsoeBuSgMJ1AANSThKXqi43GIemXvMNXFp0+X/BkmAdwMWDL
m7pHxtjqyZ69QKvhqSNxp3XuiNnWWdNoFHwevJEgB0t0z/EPZHm2U1MrptZ5MJzz8KdJqxv5E+Nq
3Zl7pdNQsbagzbmCZBDflsggJxxQuej4UBSrP6osLNEztql0exgZKJdG6bzRl3H1JPyqWc5BcanH
Qhs2ZGZ9Do7IdGanbzJ8BteGwZbYbVLakui0I/QdrAdIlWdsKwtKTq4ylzbBpzz/bxK4Hfbur/2E
u8nKVTx/6EREIBsOc1bCIvR9h0xXpFYNpvkNFe0G69HBgVjGOSyPzALBobi5GL49Smps3bFO832Y
zpwM48OXdNJUOlil0AqJgY1J7WHMF15wFj+35Zp4imh4xlAtRehjteFXDenvhscdEkldJ7lT/Tci
D8vQzoOk+8kt2shLhIu/Z6ZuhVqsqpxmNVlBjYktV+uc/S3hBZGmoCPagVKv3EmvvCc3S7g5r09w
zOAp34MNx4D2NBadT5YrLTgICcJinVuPfEtSArfKjRUQkDiyKN2uSt3LCvNx9+igdl/9bdkegw0d
4vkbvttyrZ4cTDmPdwXAsAJ8iLHVD9WqfDP3dcuxdHsu/c+LfxZMAvUvhSJFyzBXrTZIzHgyiNKm
L5Is3VexwWGz1hoOllGRlTDE41WYkboQAEgavINlEvNBkYR6JLQsIX8Sre1GibxUHC//ljWx4wBj
W+NZg5rQS41jXEXk9pAEQhbRopmJlu6Ly+So6FkdO1NRnV7OlJ/TmF/XBFiYhdOEN5H2cvvL73Py
qeVt7hykPo79/wxBy260m2+K1/5Bi1eU/xdCecBFil50OQ00f8bVOWzU/ZZgaElU5IDCp0REwoRM
kH5zBXiAhwqWCx1/edsyKZkvvfWITdnbKPasMy24sQZgpID88PJazwVI2U21tMymye2iOPMdAy1b
MGHcd3Vgjwe2SBUlhOa4jTZLPxd1kA53+GA5F6jkKJR/1skYckesXPTE3xblvn1z4rTGN29qs8Z9
Q5ThE/7BWK4rlNf/Md1adEv3G3M3kKSOfS8PRHBEn3qCfNlHFcADVuTS7iWrnKdNXAvTyV+/eqgh
QYr4wieDZ+TtGcZqXe9L6JAwNnd5WIGGTm7/3MDX9+Bo1kYQxW47IZ2UaA4wBmnbcq4pXCV2Ehac
Um3uGOOt/RcWGQCJ6vV7QlJAt8ib4pNsPr4hhQwBMjvErmBHNcoBFgifRPojo1WBd+AwItc3R+B2
oQvJgRw7L/ji1WLu6rhUEctDZE4gKKmKPC49Or2VCqKSX5vTFsvukLEoCJhIXVvFCekrGtpAgCqf
d9IAfLvdELYMTz88iQvO91rjFh++J08/E5V5trOO7XZT6l+vkZYD4pPaErl95/KRnpp+Z7TML9lT
1rOuZJz/Mkhp6D+ReM/EAt14s6lGbSsvTmxjZ+tDLwEMip6IqOQ1qH6nPnXPvcCR4UF1zirYdxuM
HrLEHb675dcitPWCkszCkxc5A4zL2qru8bxP8uPU83HK46Wj2KUmef/8xIDIKl0PQ3zLFvEjV/+3
vyDHDIAfFpjbFUtRzRMg5h2ykghqXDvTg4j6O2S1xPyUtQC1e2rIrDmznJuCRILhOECb963XMFJf
Z9s/qKZnv/92p94KRAQzaf/1CIIGFJkt9RJ8sAvWnrFl3bo3ZjSFdPQofDkqwrx4aQNuvJ55bFV+
S77wyVRGPa3LO/kcVysTWctaoRfbiGnkAC5w2JoNTzj1Mm7eMHCydx74oORuFIF9WFS1mT68H4x+
W6fZAnwsooEefwfd6U7MPBbbn9LyUUF8TqnzVkfVSZ0paZgXki70Y2bOpbXFrylK6mRngnGCjcib
6MVgscbzH+D05fUFoz5w/97PIXXAioWxHyw7C2cztYny0+IvVkxaPG46oBB+DrjnUD1JoH47t/HO
MtD2E4LD1bu3Fplv3mkH2lRkw69ASESWgFZVOrGaVr6KoQyd4saOZbLvArOkXG6BvVCD3IOu21Bg
FXYNYZX2sIebleO3BwI4UDvSBnot6sV6t6NBXhhS+4KetIt+RuFaPuUEKtLpUKD0TWTflM8MrLoB
qYnQOqhb0Pc/0+c6xKGwZEuJauCRkDwhzjfZxtSjUiEa3IhGIAP/5LlIs95YaRzF7SSeKLi7K/zN
to7uCf1WFnkTT5CKc7bk70Bd0IzhPoL98miM4pxet+r8ktU2tYUG99rur60oUL1vzw6Y6PF5sSVU
pla0rHDKvxAj/1rKdcmOiAKEyKPdEETbArZENAoaKYJ9fH7Fwuj9SZkMknrdt8HV73pThcPBX8zr
asVgXeR5kHBn+QPQ/4J8h1sPaYS2il2hhhHcWd3XiALRp2oSde2f7I5KX7JmaI/uzMxQ/3IK/HVt
jrvcmRsju4/IhNeSdiAEtJb06pPzSO+LfX1U08MFC3Fw6vQMACRZ65LvMBsE7ykcURo+rVBMpwyA
IYxiVTcI6eclSHQtGx/jkwYHLDecgAAvtK+C8kvL+YHBzlXPxacp1jUfDCtyikhUAgU9TwkOTg8s
BrbQwwiYZWNVqnMgCQEqAQ+YH3YqyKNgOI3JaXHwuY9F64G+vOWeJvInEYfMMojmCWsRnQBe5q61
QCvaS4Gs8DeAXAlPv/eVA+q10ii2mHXIIRzAXtcB3zSx4WxRi3cwjV1FMfeKoXkMWtGhRjqniMzw
rX8owV6eIAlfUQvusyFXxdzYTyPhL25ed83R7CRRyuBqqGPAlFh0ZeNltCHYcl2wjXRO9OPkIpEt
h7YtQc0onkOW88jWwmuXsJzYlfeLV4SkU0V1xSSzPiq3OznFiPOV4Z2fEcSIzCTelbm0XvtsfdNf
wcO6RjSRqKd+CLdIpH+IbQ/BaloEL5O5dM3jPWwG7h4139NGQEe3SPB9wxVoUpezIq9+JphLArt9
jIwZofHOAYbL86bdek6zPVeHQ+gjFHPPE5iuNWlwMnQW+WID8HtURfXNp/u26J+2IU4bV98ftA7n
k35jRI8+owiJ4dAdbSsexQV1HUEdL6fIH0EWjmLstxgpoXPsB5NChxlKVHlx6eJm0niaCuUQ93Pv
1rsRodSlNO/TjASZJejOtwSHvkeXAcAL4VInIk89aT0XM+PdJRKwqXspdOicuRSE44dp/p/SUPoc
FXMvKj/nJYaNO3aRC6RUb76bSm2ppOZkLYQGEDbQ/nbf7l3y9E/plps+Tbhta0d5dU+455deC64Y
RMTelWf5L5pVKAarwYPxXp8UMp730I8cipz5i7YSZrLPKqkUXDSH3UlI3orSMQkXugkywbhzCpX4
kavqgHFEPFyh4l0FAZ1dnENmiRSzKy3bXDLFG+d0iRNCptjW5QziWO+DYqz8PmWAM93FUwqBH04o
FI0ZM0jYC5rErVA/AxEfDrVbr4oc24Uwb5P5eKuxbNrVp65Pq9c+jYtMzVQf8FplLl+p0ucPdaVp
kSwoWIvFDSGmH80I9c+8SfD7/fI9PzsKueSoFSRlFYumgk23jYVHeoSUH6Ak3aOwrN2KPBP4ll/H
rjzJHuKlTLpXkBJXAYP7npXV6fzPj69QxFaIWPxiEaGvz2fBBTCiJSU6DI6Lj6t9ZJW+ScBN4Ds8
IJDbj8fvIibYNbnGU2KRblf1Z33ln1WKyzMX3asTjF9xUlzoZowzKLTteb2nd/ytUa/oEfOZZWE+
wW6SuwyIfCbYnJyok5IgY1vi9kzUaTmyjZIkW6i3rGmqEmWVpIpO75LGlJ5GatXKsNIzwZw1h0E0
eTIo7pc9HyFPsha52WXJKgOL8514yDxqd111cdfz/qm1t90RnBFcWLZGK8LOXLAgYQXp+V83Y5tH
Csh3hYZXo19+b6pmkFOcvW33ltAwW2XX2Faoevs3Yk0p4GLvHgjj6t9sEL8wsRnJao1s01DXB32M
qEP1ocnMDFCl81+kB9QBMlBntA+UKTw8Uf9tqglKT7Fjg4hDgjIeaCjo2i5aMdZ92qtnXQYVFYTJ
LCWnWm2l0XvEUOy/8FcFSUJxBb0/C6TAvOFY2BQHygV7SrYLL1S+4C2Kta4GZfInp6xK8qGLvIPV
W8xT5Jb9IlkZCQoLz7TlqYHUDXQGBXpbWG2AsgoT8XRr8RoNgIGxP/mVRFFZRHWxSKLuXe3GwUSZ
3lekgRuqgzwoUcJUEJyLvl067ag666tKF1fW6DzvSez2uxBRIJCknJvGlxVtGdVEsm2QqPgnILtb
QX93vP+x0JoJsB9ewsGNBrFkiACSopSs0INk8KJl+adowDfpCCZMlVp8oXiDQY/tJJmgOOjlKBbI
LFZwwz4f3d0C2PYHXSeSHvv/5S0n5b1qxWp7CYajaVSK2/zNAOphwrAc5Igg1aeEBj5JDsaPtEQZ
jV+x2g2kJMHjT2Ya301CnEU3s3QgVxaS6OfZcLF4NHZyfAU24lBwqHYrOAz3o8K9KdznbkNJ54GN
a12LRJSbjYv7Xl2mxCk/MjXH3OVjHvqHVT/uzxr4U/KCNMurnVxIzf5SS8y94L9/moqB1boKeN/W
IjetXyKl+PioDQFkIOC7hU6/fRl8aYNGkw/7D8aZsnkJmeq+bHgl7s3AZ1Mmmc/MbULSP1nHR4Mh
Xz285vjTNkvg1tHCxzwbvRpsUS6lMp+JTDxbOpAmkBI8HEgAawdt+Xk1FFkbOmGApN5Sv/hIoJcw
JkR+wXLPl6wINxcB63XArPNFPB8kWPECcRSOsRRWPczqG90Io3Q7rjJN3gHZiO37T6x4XQaeD+20
HArz2UXKm8tywtSsUm+sLbp1Sv07WdcBpallXF/HdCD3SxxkAYoEtn4+8EqHgMeAajkEd/GDBXoq
a5WZtBfzd1tNSqO92Lm52GcZE2EVPzjGVucUEWpeinLV7/QTmcMaLVMm5bIBJBQ8PPUCsmNI+3nq
V859/mYL4vaGEEMcA6vai407/eJ/gbNdelL1wSDASWAs35J3FSn1MNHVIO/WKPXwmeAruo/shS4H
A43f5UQqDd86RMeXGHG1zF2Uz+bdzy/xQ03vOQBYFkBEtPrLeeqCqetj9Doo+oZo8q5CKGviyIoE
Fp33R0hK2B27MNNU8jItbYiuhDP9kj7WztRxO91KAXwaU4J6vvO9vV/0ur/FQ9fJL4IoSh67U6uK
r8klJ0gg7ZtLBoRJv1Fog6/uc2BRyi7GAKJRxeL+2bfd8vP4zrVRh0u+hGBYIEzPMGYeUMcwOVf2
zA+MUtX0zIYlZKM0ReJ8S9Gn2qFzBP57kpmXr2uJAb2ZmEfwInTBs07o01b/WPHxvPGPI1sBCZUQ
FzTDBsbdmWpd8W7BJhHm2PeUwxGmZ6WHKYh5TQQMj0GPx1zOd6smXC4Heu17R684GKviOXAjHWu0
DJC6ba9o3BpR38BF1yhtI4E9/yQbvAintiQxByaF2vw2ukl0vpLnuP0W+zum4uBnISqVehIEpq8L
Z6MzeS17PqUqXfpSS4KfCypcC+j3C5eOstfJb/wYZ556oQWhKDBvgh8LdOe9vbd/ksA6gLJ4MrZJ
n7qGh/MDwnoyfvfttcU/9kuCiufxE0ks8MpPDmmwOEjHEfnkQli/fGM/+dgfF0cfhsapPDUSNhf0
LESr41/LP4zy4mU0aQHHM0/xRQNEVLWn+5myyIoN6Cm1FqjaH42F581sjivqBKKgY575VvMS8Huk
dfwz0nL86zPuwcGkwkifv9nimbX111AljHkyu9j7z1bfKkPaApoiEiGP281QEq/eoV9E1CqPF3Y1
ffu05Y1EndscyrKResJnyjY5LAuzI2RALTAkF8jFXquo4ayx1zfmwjGFH9bCfpT9fi3+CUPVNAcX
2m7tM0a4XzJQU33Hg+9zmhddeZ5o9iN/HCR0euxhW2U3ygUtuQqnHTk4wRi0Qqr9d4c3+Lr2VhlX
coUXGVxzL4MiYr6yCylxF8hlzDaCmGoXZA5qDz/Hi+TFlA+UEgGlSU1ncwpEoo12cEKpdeheJIyl
ma2qPHJlxO73J+pbSG5LbEFOKxg9pHd2+eO05Dc4xoirp8AjkOuU8vLT90sYfNHzF2iy15BBKVs8
QwJOX0RONbt7RXDhXCQDKXaD9xWbldxbeu48WUBLC97pSp3SNBrQ93l+j9cFyZ7Tx9YkUfk7lkxy
IJZbatPwBQFYSJCgmtP8qYXmX5bFuLUkB5GPtaS0Tln1n2PRHyp4MEZ2S9MHUi7m/+bmeqoH1Rgb
vzQgZ1oZJ2MRuxOU9MACyDRHKKOouc8QZyOnu/LPl4A9ZZ1M8Wm0uXaF2Bx+LxEiHZRweOfSDGqw
usi+AJURM89hVsT0XHEymKigGvDEcgy2K7KZJ5+z7V4gMU9SrRsInGYssJwkEqwDrpeBm3QOYW+2
KBYh/WZJk//zhrKfGt6wCaxsmhOQNLMNgs6Cm1UA5d+jZycFPNuOGpky4CjHbqM+CLZuVHdgl2Ec
mf0uLtTTrBZaf4tJL8ZU8V0fF0fsD04A7FfUigDspTHPY+Fcak8dGU6F7QbkWjFCPelfMytzTNwC
yie28GzS7wfvPvI4rJUjfeabsNaIn6FZs3TkdMw7hHOzsHxtouSR+L15hzzItHRQNADc0Dwr6qja
FbGh6//jRHlePj2BbhWpGe/VIXMAAeaZCpg11uWxDcCLo+WmPiT5ONBt5TrzwMI0tLhlX7+aG5Jq
VrYB+nLVMLQg3fJGwb1U3jN8qztYDiavkWcnta7dS0aUKSjczQoZT9IcFalHfeq8VhRI1tivEnNa
kPZiu9eps7CSXV6zHw0mkH1bLH8hObcC/Fx/hvykKT55BbIa6LRww0z+DVjTFDq1VxP1WtMV75HG
siyQPU9BlTKFq7ibeXCQEFRen/YkXbHXpy0wqFFRPxyez5YFd9qrnHKwoKm0bUbeUYtOxOccZNmy
MgvJOfQebEguc0YMkHtiimjRM480en4GTh7MTdlEVwtHIDklMMaVfH+vRnlJbWB7Xp/0po5+jhcR
0iQEzbAwfbL1b1yrX5yzcIsPRtI+7gkadjiL1y6gG/bKEW0/vVSyiyXhYhEsQaaJxHvywMqU7mcH
TfZtbnefrmcCWqy8TRCTUs7teqEZSkZ7npNRPYrxz8wX5oX35uu/IxfYvv6YjiRL6H6fo3DgykTk
EChX0tCbBN6mADXbrP1XYv67S5xXbKvkIzWECqxxxm8m+9uaaeVRBVblSg91ag6mDk1xpDaDGtl6
HshMZHvhx8ZXJhh4cxZGTlondmqrLPlvdKhNhEXavL5eduPkDHKG6dypToUIO+C+AhuM9QhHWN08
4p3vJ1LCTIHYAn9MmyFT0WeKzGdXTykX7sK7bytnbahKcaYC1eIRfjTQLXd/58lDTveY8CtngJJO
nqUI+lyBXRJClNthXlQZVw+aVza1VOo31yKZ6PY7szEDuvc1mx3OEqZAFRYM5KypgKe3Vm1seHXv
IxJW9kNoqMKXwBzSpCbzxl9cibnfdXHQl6I2MQRb1V7JAHRL4FxPr+4YkePcL0WvVFLiy3FSEWul
AIP6MCwBSbrhTUCKb/2tgolAjph9QHd0DiuzLs/jK6RRWNYc5HixlRoWe1SPyYlif1FmepoyXZl7
AX5ngxGTtbtUxSTw4K0ijw5PnPZWM/FWad4HbaYVAvsMKaPTatHRVTK+cMh5eeJKEx6HuAHyYmJj
QiKIJ2n5SVTy5YBBDT/qSW/oU35OnrorXiuBoqB5CgJ363FSRHl1jVf+zNpJfimvGftxGuN/qoGl
imqtTiyQC2c5/Rn76gJvsimfOxLLEflGkvqz6G88jkXDwg4NViAKyayaCOL+kw8DIU92IEt798n5
xxijrsbVL9iLjEC42xWLyIvPnJ0/9uaObA4e1sUul3MypKhVcZJgTB8S15ZeyZJfVxnaKqSmQiYM
g2uPOSaWne4Hqk7zT8eCevWqWVdKt6Qqx8OBOctwbfYGcnfRa4G5hiUQkC4ldpJ+2jwLj0S8mj0u
2f/6sq4V2ThgmBVTW3AYGhLwxnC3npLdWcwLQ7GUOz5IF885tNYKMABUSIqK5Ri0au7QDLbx0+4z
D7a9/Yn++7ZKqWqAAAp0o1qckhlUCGP3AE4z7jWUA9jgBCBosAk7yKOMgE2dvCKUX8Q0ZS6fOaCm
iX4xw0SdoMWtp6265o29CHo5ctZ1Upi4mkstxXDIsHqvAcDD/1Gl42Pe9xZjLCJI0zfnhA7UtbI6
SeXtUov0ZM5OuzKpHOBJtRKUqtTi9lS/xAa8TozVKZ4ROG3nrfG23IX1j4huchAx3N31fee+QtsR
/Ig7aSppGKlWTmE5PX5xx/3kamimvWd9giKn+O6vPY93unBgXvweFspzb5321UPQuhvSaipGbgt7
6hjn8vJn9cG/04KLxmlk2L7tIy7HzPP79z82Pm8R/KPoBn+7+dvsduIlO5TAiGBItxDwe+baWrWd
z56PVzrY2nGZv8lkCBoAWKeKi4hYe3AhzBd8zvkH3OLTi370qY0nSuCXx/9EVk5YXWcqeMzZ35d+
LLc+zLaQCGnngC2jejlqbuCxLAfcACiMLf1kY6T30Nad9OAxt7Vqr5PeuwVOMmyhWQF3bMJi6/EX
Ng/g6RSs767sQXmjkVNHxJ6FP9m1PYK9SXrgK5VaF4d/1aCeG80E2fS+BrcUe7To4gWOZXuW4Rr7
nte/C7Gr/bSz/uOTdiPfy2XPHD6A1eQdeTbbIrRBZFuOdY1ze3xMRr0AVusgZWK9+P1XdBbIYt6t
w+fXF3XmFGeFgvb8xMzmsGID27iS4lzWpxiQXJaStm13z/xD4U0FnplqhUVeYqF8Bt6orSBHJVOd
J3EWB3xr7jC7t/+GiSZ4NEwb/Pu1kwW+/V7ms5vh5kWbpXCYKpMXREtFkEhS9EPpRpuHIaIlRcb4
viAQz6iscfRdERoVlgVzlK/NpI522JcjYoTmaaexp5BSSXwdHH5gcI6S7P1dEvIuOJT1K8xooSJ6
kyKUkkwAG/YuEFhsfg7yRUBZomNAhW0WtsW0w2bA4pxN0apWHrJnoKf3+vkx6IZ4xYFaND7ZatlI
l2Y9izHH2/F1GFstS9WS21g4qixty4C20RnXcnNdyiNOD+yr+JSrcjEKn0Ko/gkF6O1c0aMFfLT2
ZLnAQJQyAXayq/f68AvirDG2R/ICHjlxbz+idJJ8/tVlNWxyx0ppXluqMKVVvkizFAQvGQehF2bW
nSFQ18ohmP9QH1WUjAxOUdlXolp5DcatzOAXOxPriQNCyUVuXaX2zjPlZ6wyvZ6irhv1xbnCVFmm
XrqmvqMgx/kaq4bVo8su1MW93rVxgYnyYrfAiE/t0t3gbe+3uyHLqJ/4QNM6e53f0XsekwAtD+Ss
Ag6i9kA77szC/HTJ3MC7ra7tcH1gelNoL8MaX74jlUYos4IJTDk8RJCfypy9pMgRl5NLMKwbuZVL
z313HjyQwoV+Lik8k90em4BnTUpVuV16eVhmvZh7IjFJDUOYbHq9lHxRdKc/5JNyEMjBsfUkigd0
LiQbPArz7YkVSkmk5HcUSLh3grRC3sW/dBjZLqhMnUDdyOGQYPce99AoADXyzEX8lpCmxMgpilpl
UGHtphkToBR/JMMD0a3REuK/hpWxDFQH6yQx6XUCy1P4cbersGLa/tunsHAoRvoBdNmZ7qnu70fC
pDhHx82h7oyN9drlRMgR7TwcRX/rZWip2KewXZrH5qlBJXXS+Sm+vwF61xqH78+cRqQJ49iE6lko
5jacrL2m2OkbjaEcNBXjQlwnALQMULBagsNOpTwVIzwNV0/QbrpOJKM7rigW3R4gy3S6McFn4Z5s
GAh18Bxfkqqc9PlL5e9muJLLBd1dHchVUR28ZlfSYzL4f6oIDxYbUqUq8Fz53C59CqOaGAOWNC/h
Wg22ibmTOc5N0P81GjMtE019xSPumHNC3zoJHhrR5QSLz+BYPngTlD2z1St9W883QlFQex+MPm3J
h0E07kIYE/avqG4BLn/lqJ9omtM8s4MdpPufyt4ypKuI8LFCmzmfbNhcdfho/7HtIpHS8vsUlulj
uJ7ogqWYvCrFRYajZ7/1/XNbqC1iTTNCj7l5uRqtQjnrSykUatCRYUIEXKUg2YRMuGCRpAfWaPGu
nng+ByDZMlhzH8woTS3K5LVmdWluk+O7ayjKwYWmHtnpqcGDJDrAs6TsbgcYhW5OrsxRT470KlCo
qxfj3KafXNsNKqd/nMfXcwRO5Sbq/L7WlrVMPM6dsDXXHYNNIZpuzRghlYB/Y1Lw+HKHEpb7yKrI
53NIYzsrU3DX3MR41LMEwrabLwr1rc9uuw2+a1sML1NMZakX9M0WrxhZpx1sXDRxGEsTKHDc9mpC
0T8k2Ow/RUe0/Euuhv1o5KrLy/vkmF5vRTkg9SMz+DZ8lICQDPytPESR34nB2aGNjZrHtO9SbLn5
BuRORz00uY3e7rPub7Ks3OsOiVg6eapDu+dDQqDCOlr3KGFCp/nF5otB/ZVApY2Z54VjYGCL9kV/
2+bUQCyCwuhg77eBS7A4otG4tk1Tcme39en36DbxRWJGqbRHOZErBlKytdryTC0mHPi9TPLiYCgZ
b/IoNXlReMaIA90LVR/NsWpnUTKKYDxhyZSmkCel8Lm4DNtFv991jJyK2cv9R2z9CvaiUBLj46hX
dPDbv6djGyebAVjOC3QrQxXTZXmh9NhSm91GjEJuJHZKY80uN6OGl4rnoPas1aVM6s0ssxAT/uPc
v3B5NqH7ZdSuOClXyaGnmBdxNrwL+zpVoGwC4VAM9AqmuLasNSJE+lZ06E6w02BL9jxc+oK1Jr8h
5LjopYvSEErxzPUt7HG2JSXBBCsITzQKmu9W7XuLvFGEHh8WV64jaIyU0pFoAxnDCUCsZwYU5ykL
MeSKbInE1e7ZR2y/8NKEo26NHfNU5qIjGa0rE+av1brfbjq8AR6iz/e8VMuY7oEyy0e4FgO8RM29
+VAhd2RaHfdVrRCsRqjQvkJTKNOBDHeQW4WX+wQpLLjVghWis85UI5UGXfwWXA9Ya6GGLx5C41WE
nZm86P+DXBxJT1Hzj1OskRk2kNsZy+XLAooKDJwUXOEYriSaDy2R8fvkTIgH14CC6MrivDyLKQPg
X7huCYjGPys9w0jytpdEB1SRlJ5yTp1WpIz6/84Yl6Z9fmnCxPAn578v42iSZt6mHhmSRr9eF2Ug
S+N3cUynPtF9QkxQIcKEIwO+EryegKEQX/f4O0rNm0apiXg4P4X6MyysduDuYmbvs1uK0S5PfVDx
y0Xdk/Vm7IWhRCOxSAo47RweZILKEa/v0IIYEm9EDfzh2pEz1jE4NKuB+wVoCrTfAcsu/u6IG56i
5v82KIzNf1hYVmz83rr83RNyoxHvat0oLGkaAM6ysCECWaV9LQOYtqrZDuRXSq5BkCHJI00/hZZe
YrfIp4PP2YjnZorO+U8OaV3nx9eWR/+gVH8XFSYZ99xQrgxhG6q3diV63fqMLs1eFqc0VFJWrYik
caZaY4WMrj43DvtJpzWk+vVAXShb/8X3+hb7HzwW2PLdk+Tb9VVhCAPdXMWYEmEL4DSyYbUvpRDp
cSFj+VABKXNpglgefgcqzLNwCUnLXeGOSU+aSR4DWO7Pta8y99r7sFC2RxLHjk7wCKSkBSpq2uSr
yCFev82LwzWLgtlHTO3Xn0mC6BJYZ8Ii8rHa52w3xbLBuk/60gSJmevbeyUr5QyoFmltPO5fDCyG
F81Y0n0pQj1nq4s77SpN0iQHXDhtwLjsu1gm3kRWaXW7tK47drBw7/Q7vfJUcT+Cb/Ihbhrnul3E
u/rym4PvUXqSlEtAyntqRDukIg/YcH5YFgs61+TrpeqistD6WOQVh7NSOMP/8mxXlTlMCeIfaUWG
HXhnaB0J/cAxhcdoktu+C1v1ntCoZz79M7SJO0QdhJLnRdkYB0T5cLdMwMxcWeA2G+7qrZ7q4eW0
XsFfFeGQlQo+UwkiaY8IWJTMDxM7YyygxP0t22b/oBe0p0VfB/3qq2d/tJSY/00ok68uirB59XFB
T8JoTfDfJrYpr01/46qylVLjOqjvD0+JNnMYxci4Y5dO080DiX6DQPlLHYbBbh4Z8zpWB8M0VX4N
ZPYkkFG/4qNo3VSJX3zWFbtzFtRdQftkrF8iBheE3+F+ZqmI3ODdW3JzCoJ4OOjtXQ5KdGILg7KJ
n30W8K2E2t9Kb5S+caPEpcq/hkLPsdiVzmhZDtiAkCLg03XVGqQH8nV7NxxbzSrkvGfDCidv89Cl
djQEigOtB5TlPNSikSsZY5xi6n31WALklfFQgGr6jd/HVyWbw0XkKCkPlQHCnHGnRLwhG1KUURcZ
l9OD/Acnodyg8YO7dXQkVmzNPBhRKFdz3DdJGrdpr5CFHo0mbUM7FB53eZMOZHWWZp/rxSBCquhm
e7PctBSODFsfvTB5Anvi/cg+gI9IfrnIfxgpEEDCDI6LhaL3IY7KnXunUxPhyDYhutIKiu4x6vnR
7yGkpamDCKfKVU6mkdvzHvUSoTFG/x8xmVdV+Yr4Pr+yxQuplhhGuM3b2JL+cVpPnCK8/lgvZbXy
fA35L/ojIrU7sXqVIO71XA6Hs6Di/bBv67COd4HSS/FCFA7RUC2XDTSIH6x2bZ5Kn4D3n0Oj88K6
q0PZ6p0z+wB3ZsEvba6ENztTfk52DarwtsEZ4SuHU4O7WM4e//5UGWiVAFTxyiSXVrKk2ij+5bAk
0BG7kRGYOrF1Nvy1ePwYddbouqBINrQsJt3qLhzlneZaEsGDpdsuRVVqr7RB/PHxbec8DzXL3Jkt
5aQI+wv+E4aKLjatvk3VjscmbEM22bqhlT9ug59Gu6ISEvIos68j012RzANsHj4tz/QFtSmQagN3
omf5H2dttFnkl68rJSWcxCe5EEl1ndlBoVY6xyx3bSe6MaDho5tkuYFV7GMbsvSql4rYIN+tlX2m
V6lSUIkC9t5ARNeMDOmGrwMFEyQfZ0fOzhJ7iiTX+VWeMDPnDK5D3u2VSQDxlanHwoaqwgk8k2Y6
70bMZSxHr0GabCR2h3tBQ9IGHz5DLRndqPv9ZwRUzTEGgUTF1xFu/ljj37SmOb+3cD1Pn32sqBcr
btfuIbKYrcBCwhv88YmM/nBwaT5P8fiBQBAY68new4FONqx8VkiFAiHtNBxzDtFGfg+RziCD0UFu
MqJmBxl0pn+Q8J8/rTUHMjqiJYv1mMdXkH4fwmDEgrshOzNP6c6T2QSSiaZQucG5rlBTM6hkH9NU
fpySp0qjpZSS04T7lYg5duQRhLUqNUNxxcay8Cf+veP+gGckAYKHwnsH5A9LOxpxRY2C6bnpDzcQ
1YyhouZcHSmP2WfzKeYFasATL3yWITovpnSKRkZ0WeYru2azUw1eV15UaBVidhqdCWjG7ZKMkd6Q
rSqWPlEb2nvwPMgUlyB4BX1CnNdnbbElzJ6d2dJwmSAzcPlsbceWSjoOyAtAORxYzU0ralVmUNJF
DmC+H6GO6odMAJ7XCZYBDVLdDKZ7y8nvqURQEJ3RrauKVZdN01zEKVd6OUuwuFTN/mvjjkA9I4vx
HiSRsksDO3Q+oX3dAyctkgBtb1QYj5Y6wGdtS5crYrodx80Jge+pSoOL7O307uy1avUyo+pRYxn6
GesCYQtYXlZYBBx5KR0iLWKFApiDvhKuBoYK/SoVepFv4mDMDsDT2IA1REZP2eszPGh7nxdA/djR
P/bN9JJ4gt/32T7wLQLkIu/XJ8pBtrc5tn6RYD59ipG73GxeT34JjnRsJG2pulQdI7DD5TEwVSNU
ECrhuleI6d9Rj+ifnUccdjwXe7ose9ohBTCJ9ZJKdJu1wtlF1D5jLvWB/HmDk1Edqe10VGTl/wSd
/NKUfkn84lXWi6FpYjxZSqVQ6DgbMJPLNJDjVDdMPg+PNeafjiCvSTy8Dd7LOmbVeWS0YObA7dPx
f2ELJ7d8YEp4PxDnRVadAypDqke808gTRY/zs1cAYp+JHvZ8lkycjn4jbpGWBqNTIIPTd3lkI5Nr
YNnKCiIPmAnOR/BO/uOsISKk15oVrktC7IsPHEv0IqIsQbW1CJz5p52B5QSE2O7cFRUiNueeAOTB
oaSi7QRolOMHyTErZlNYWglg8kUeMWAZvQOIKE9WUiM9buyJXT35yYt5XSc5Zmx9eaeKANC0iznR
zWFGxQdtsfA41r9Lem8QFS/Xm7s5lqoOPk1NiSrNwUGDB9qygDtYThSffJhC1odbI1WWiauk/DIW
ogxytzqPeamdWwmjBj4xBV0NBgcKEPe6Np1W2lLJS+6Ad74YewqBsCl3ovM4VZpWFyEVz4c3zFwf
zbckV7jRgBr272Hh5xkieUY/q6elE62n2bb3v7lCzde/Q1aZMgzheDBUl1jmF+7DI25muM75wnxh
tHpNbHqa14ag3zYMlchTibvS3VPFrQFNVtVvutyN1Q9JUBAhcmp1BeYmsGg2iv/hB8UwaFFl4LO8
PRFWB2FmewBQCXvgt6ct82RsrFRuyADk6B+oUIJLimm6bzwSCl7ZzK8s4jc646bGzGEwiNvfENLI
TsgKvYDgD2WrwbuFrmj9oLv4Do/Lc6T1JNKfpdig4Y5qGv6jB5Cy03gU0rAH/D3zck96tdUP5oEh
G7SANFYxLP37uuArnormtdBMoGcSLpJ9Ufgj7zUM3NWwxRY6iIKD3FxyhtKZesAppmW/3dZfu53b
UuoJJNUZb5POHf1f/VrDCkxbmY8Ob3cFPny8RepOUbqGxprXzUjH3JrD3/6GtRmujM7TeLCb/pBB
jO2mTiJ5e7Oly3cqVhh6/8yYjBxLRLQk25tXovJj+4XvGSKuqcKX5vaQdCBZLe6Jvycqnabp3ceu
fb7RtJzuVxFs+ZYNH/NhURadU6xqXSthiZnofWWXbW1eRe8E48Zz7J9596HdAg8t1YMgrN2x7hgh
RnYhvznSW2S9phmBzncg4C4dUNoApp0WM/0MqNtR+esV7JaKXymtJWqsjJQcEce5Dw2+qVkKBC1L
XR06+Gg1H17zuyfvEoEZCR20EDfdGSx11rjiK0P7AacBY41hBCrrK1Ohg02T3yLzIeE2W9jbaP50
JTrqQV8qi4eKrQLTLVa0ZWdSkHv/CsIwBbxRnD5CSIBdE2IBoAvIhp+KI0qJ/qQ/EoRAkdT+InC5
cWeNKyl3pWLEBjGBjuT3puf1J9FrjXoM5FhgK7uEK+wqDmUKB6tNCED15ZOGp3oKFtadRp9Rk+tq
HaIXX0+ePfJVrs+0hcBZ5io6apsYi6L27Lqfrmo0tclNpzShhprzaNeLq34Tfvp7lbzo0Cxw3zNp
G1arpp01ypQHcwkzCNqHYqxFomOtDJ2h6n3nlPvh4zzSEPG05vfBmD1YsitNJaSBJEMakgwexn0S
vjBVska93eEbSIgoTw19vdgXpkjIjW655FTS4DEcgOnd/0WFhVr7jmQaYSaaoTdxV3EPtXlCxsH3
iG7iS3fRMG2CpBMALllJB3o36+aJaFUZBlh5mfd9KfA7iU+AROWHQ6tWIuyQUMpwue7VWyNyUAZD
XT/qIfEXrKoL56KGtZJvMvnfFO5qt/fmOSFkU2oKym67RvzedEePpP/kfkR0suNUUxKlYG5Iws07
Mh9eDBLNi8nYG828hvu3EMFGvbEhnsaSriOlkdat0wZ5FEUH5dbHFVdCegWwN8E2Qmuqia1F/brG
cAU/1i4eLfOG56OWIgVC63Qy02+wwKw7TZOXjaccuPc7LW2o2K4fX+hux+DNIbT7MqOo3fhrl6Qm
fGd/Of49qjIlZ714MqenRedKRj1dCXIPAdX7kGbp+39Hdf23w7G9Ji8uDqquvYWe78prIRZN39Jz
mxkQj4JGxFkH2Lt06V8fv4vcmMKqtalOkril2JpyB8yEKAIeggYAIOa7eJCcAWqQTjT5KUuONqri
mOLsqu/F5Qvlxats4tDdKb9cEKW3qK+q6MEbWnFR8WUA9gI62pfyRv1o1fbGhJqV+lwH9VNH2mF8
DViydtbuigLaA7v2L2fwI8EEltidBZDtNC26X5Gh0vzcU3t+rirC0npkWNlPb6zpA5olf/Hk5REE
pmN3CvWmdIV8JDqRFCE81jym5plfFT58aXzHirNLhpzvQGn/jTh0RENtaLa+KVz9uG26Ey7YdhEs
Nh6DeDTuBP9SYlkQFq1bwDiF0rLpupr0TINZWJHFFrb7SQqQrwdi1m+1SddjfYcu8w3WuWIii3zl
BEozLzTGN0/8kyOU1zJHcv3CR/Td6ZOdGRYOOuVLU1GKvqfnI1rluworvRMxIPBsrhRyfnzSLMa1
jBZOPIqiGrdJBKWPJlBDZCzBQr3R0Pae+ErvB6bUeQYetBt/jJWNJPYiHXrbPhLZ4eBXo/c9lb8e
8noKHO+8wnc4uFlMjfczm2ii4w1EY1HQIISgzyuK6GDxMgAThYkfhwUAuAcxd3nz8s1dLS1pWAed
PeMvdS2jmArZnpG+eCmmNziOqfYRmyfa1ltjKyMucsIC9Z7+HtRInVIjxCA/twO29k5n11rucOV6
Wsrke1JH+3AzbGCiyW7S2iXPjKHOmBsRBGc3C50786OnLkJa4+n8TVhPea4T22RkK4Axk9gwwW1v
mSTEmcOjlagnEez/0/OaXEofCBz0b3sLAthQ2SWiPyM440RRO1GlllQZm4salv7hiihdGu6p3+/k
fqm1Z1vycvkttNn4fUWMYd60YpqF08Wf646hKY+sxfmdxUtWzuGsMQOemgvAIJMyzHjcKJvVg5ZI
+zivkZMOh4MdLQUPhiCNlO70Kpfs6PA11o6yarMTFPS/9u6qvRH+964bl5Iu+4HxAiDLu5OElCbI
GCUTVqg98t4wYkgFDs+96TzFS4DyezdK09elrcNnUq8bv+eIMZy/8kl1lK3o9DCvwHf2O7CcYuL7
xKmPCNFRI0AKy95a7pkvXJ/rkPyOmpQ9lSvPciA4KJkbvZQ//0YP4QR0p+2SrFk7p7BcCDuEHJGI
idlZkGgcf+ZXuh9Fg2QzYP74Z/G7i0xC0osCkKkHOwBr0gk6XQdqCZake3UMZl+dLI56rP1DP2yM
xok14XcohQp+F28g+2eBcqEPQJHbctDNot130Wpu/hwcYdA6AE6+x/ozFdb+B0jY2dvXY7k925ze
5beIwpL66bMlfvvfr68dlSyTCvdDRtNWpcPBn3fWGzRNjsN+ykAwUcAwXSQCn5tzaa/QNwJ7BSX1
T443gNvauEX+9qV33CBRTZcjMSpWPLrrzKdzgNf1D4qniYXufFsKy40aIhsOJY5zj7gzAuqFZOsP
dsbrjahxV+GZzbutruPAzxn0XVDlDE8ygTMZG5e513mgoukD24yN2748rJ/R81MJ38OeDX6LBegM
EO3djdGjpBlMkj/fVDYtNQg++A35iqUMMB2ADb9SOWxz7YDgJ/r5Eyi1pbirr0abjG/UuENk4b2B
A/H2ARXiPgKlFBzDEa787QOxWlVKRnpvpM7DqqJMZiWvE6U/2IS4VNy3dG8etPOOAIDuil/EFbcz
EaQl0Z/QUQyk3p+KM8UK3y2U5a33hLNeSxNF4ogP5MRzySvl9h9DWiAE77vyL9pj22NA3eEWTqAx
xXA86WLxiCZG4jUnly9QixmsFudx6Fzvih5tkOS0QOiypw14hsH7orx9KU7lwANZq5Y/b5gFYdhL
ZI7KvFjvbA/0Ii08a2rC53xO3ZIbiQrHEWDMZPpTZX/RlptZPoofVYU0px7KcJKLW97SD/EXh9P+
evQLClpf5xIgoB8R0CtXSGDCPpS/PXyz+sepl00rNuwq0tPzSrXCIh+JMtGpcbmdilXkvMjAcETd
XY2BTgWnIqh9g1WMdcQbbWnhH90JNAarTZqYgyyiP/rTxBzShjtPauODlRUlwBO7gvlylTXUt4L4
Fg2J+KXRiJi65JnH/C6nt474z1pupiOIkPEe06s9xT5d3eiMDiyXCfhDShjpkvvTh2We4fv08/SG
0TAnBgPCJSHv9d46OwYsORhIg3H4nXLpj6TUmb68pNSU+buyWXpjQJioC7fIFPfwsLF68RRZtEoF
CumlfN7DQTMbC6/D1EVY12hA6tnELAcQpB/7iC+ZS9G6P89oD2TVtZ6wuMPaniSRXvZHExSP6rsV
EZdHJWgkoLB7Pp5viDhqodsjNpdvHR1aSl50HbRd8EtUlW263kMk+AonJIyHN+y/gYcEDMyqv7pt
dTDkdxgNJdPvMaNeHOX6FJgj74AefCfNsrNOmyg0oMEqj3iYOtuzgFRpHZyuUFlpRgtcaG7CF82Y
JUhg0sHRFWJWYDxvNYkfvTaHGvbGJgQied51IPN5IEe/wIDcwLn9eBqCB8wOYGPXlGT+Emaiclf0
yEgcEbqAyOD68AJRZSmCio5+k+wqwm5FUFW6CpZKAxZnmyG7BMxtUgjhRboeVCSCxYSpcX4lZ7j8
IgWvob6SxjyC8renqmuIWr3GpkSYCpMLIJgiiBCiz1rbgQ+Q9k0ouDrBgy7YF0Vv3s1qHWY0M5eJ
UGEXyZXoUzgNENrBgCDkn260NCjtaDX9KMlxe4PZIAIHvRlvpsicLFErwAzFhrP3yQU7VDXhPWMB
qRs7U25KSFjfmBP2v0ymMt/XY3KHHMVwbAtyLkc3rmdphyCwW3+/JZQC0TqxLLeXGrEHnDulTXXn
+c2j+aUXd/Jd2DQzEmw8kibXxtx1Aw9CCnGuFp0LnxcbNB60QDXIgnWbO8U3ON7kTdlKfMx6oVWV
MjOOpMgSdaS2kjyBjRnAhCEXpasn/Y6JXqPFTS8J3kzaaeKvVzMCE3SZB+ilBaWrVwyECF7QYLQG
42lIXyAF2dbW6RIjlua2POybNTK+CW+PnymyKLSppPjLpyYjy/Qks+TOIhv6f3udD9kwUVl00XmS
24KAFgXaAsxiHor03+hifUwOcAIlpxjTPmkqt5N2sGVfYlwRsRwm/R8RCdtR+9/h4Ak+50PkNuE3
4JYpLv6qPywkTaQ2/JKlOW9mIn/Aqyw861pWjUz5j2C34I74biElin0kZwf8yrXaDiY+6Qa437ED
LV1MZtiIUIa9Sv8weHyshg8hhdfbh4p+wIRT6exn1t0brSwL0gsv7720Pvm5bbYpksZOLM3927Lf
1r86n8A2AYYaXyqrXhQTJ1E7fTelvaCG3dCSynxC7YISKB4WE0+nOlbSU8iitDP+4nkj+6bUMjTA
UFR2dM1m4LS2+51HFStKGJuUKEBWDWytpZlAQV72YvQ+RwWBiLzNGV0OKGehcJrmb3/i/PKoO8qa
F4TFg7N8g4fYHam+T6UrRsMCuXnNV4nW4R92IRA9CuoBxKKZ7/LZ8BAFeV9A9+FYil3MaGYahloX
VZO8+nuzhVP7KWSs/gLLKqzzZpa+dxXjNIWaq/lsy5+aGjYkGAvIhPzmoONuV+ZeKS0x8kayqO7n
80Dh8VM8buIKETJA6AHMY0e925tzzBAlEN0Bu8fCAIcen6SPu70KGjLvhCI0KVcADTxmunHFW3nS
mHay3LjefjfnXNsBRydV2wRGKv4fSMcjC17DtIlhbRYYXajX4JmYv8+v0vuVE8jIkvAUG7nHLqiY
y0s52A6ATOYqE02q2MNXenDmgB6ki7N6H5pvN+UeGKjGuEi40GAB0QaPO6hymg4CHxmy4tbrJwPf
7ycQ/Xczc7770UqMmqKubwVqwun4hiSD4s+1hClnPItUS717X74ERR4sOFe/AXoYW68P8D3Z13jR
KwdahnNMnWWVtxR3BT0cG/l7bq9JgHYIKuVyq4Fgie3O+UgpaR2t5A6G1aKrF/mERcu89klOyOZF
7Et2EgLY8b/BWAemcGtWbjwe8+mFKb+uAujuT9nn9wSBA5xk8h81ywJu+TubXBLSN79+o02av1lh
I0FrIJYDhrcdXiCMhHGIj+RBkNmFXGJhtxTx/rjtlVMueZ+EEXK0Jfn4m/Zyp+wyu+ExatXCPNcK
7xWOcW0rzWvftK7A4vz/4ehWccBoQuT3TdXaEHR3CYqbeW2SmPTX6w15fTvih8pFAY0Nqb6quYDd
Su/rasagdMFgU/PfLy6TOo9Ph/cTsugjy6GN4Qy9Wkm8Uyq7ze8YdbO1L6krv7WPoRtsKCtWzIap
d+Oi5DNGvRfHvvelXNS6FMFABI8XLPsJWhOBKL9HyZWvq2N4PaHd8QpLKPkYH46Nn3td1v+r+tBg
Zllh0mlEbfHnOKFQiRDhdzCzxR/PH9pUhwMnyHMdbacwHrBZBQHdDKjd7WjOxwAp2gid/tgfMScN
WhMzfORPxMhspO9P1j4t6SH8bevO69vUOnYvjC1jNZwYQA/oUvRNu80xZ//8TOrdzepq2T+jLHGs
COT9u36qpSYaSYX1kxoF/r2mFP8+ZAzVMg3yR95atQwqyY5motgeWhqfhN4pVa7eYyVWEK6q0aN2
0UAESRqz3yLboYROyIhRnsiHrsCV394Zf8IdgC0tNF/eaBWun5gmqCpAXhtAnLhHT4gJp7U9kl3f
6vo2b7OqVHB2o5SxhTn5llHuJ2PJVy8FLUnkY2a/MpHpa4qMSX8yLkJ/y3ZqoVRN3qEWEGzccMO1
Ge/10X9zo7blLOZnhvAdtBx9YrocszwoEfmuXgJ1XabIdDrgt2Jtw5xBqHiH5XTEiubttp4sm3cO
b3KJxxUFq2giZpzCk+YAzJoeccvYopH5uSVI3U2E/AIMFzlxzitGeV3UcZfnH/d7y6p7Mgwy6AMi
WTzhIThPdG7KtWH8DSv57aBi4iBXR7sn8AdRmTGnlUfvgDyxd4sjerJyO0szm6onXJGzg3zp3DqW
VI47806Yewc7O4A+Q4fq+HB2zA3C/UA66JjJ6Mitg33TXzv3bdsQnew9GrQiokGstHJePrpfn9B9
Vn1F8Q32q/xLuVxarV/Vw6Rc4YDTYonVpzAVsxUgLBj5JgQYQHiWerp6KgtfbNp88ER+aDL0r0Bs
gSTs4f59xdaOtlS3uL1qgpKVM+P6OlG0dviSDQ6KYBsh2Kw3YY++UZyI9swNogz/WQfkMzmMAwTC
O4YsiMeSznKYrmUTKyLFeYH0r9KpSY2j5IqDGVuY7zbF0jUvmx/812hAphv1RuP5jrZLRzt83Fow
p0JgRiSKQD/R+BEzKhIAm+oWYhXBA+CEAkrto3+5J/dZY0cFi8CaWTHDymVsIZpQ62bDhEtx1g5A
1Oa2MSopNeshFcLfdb913dIhl4S7ONRK7AceSftND8HT77S3CRQRjGhP1Oe7sV4dm63LqUqnlPN6
pDQHNHXeTcxgpYS65Ij8LKL+lpFhDP1qWtuZYulNbxbVyxY3s8Of6rYqcKlhtCviqg+x/quN8oQq
FIA6IbdMhSqHJFCMdf6/QLC0JnxXgXUyDmFSqI4EmnQoUM/8cIN17kduc/sj+FPxZ770ax4X1kGv
EZ5+Zw78s4D9TkGkNZSQj9kpDPdqW5nfuFn0D1KlZ/WUqJSofvD3nvinOczmAHeXUopwpRyCLI8P
bQtPAge12kVWPIJ5yy9B3IYPltOXItKYpbydT4PyCUbcs6roe/eFRPhfEh+kpdeQdQKGrlOSj8Ms
+/jIFGgqXIzkEm3Z4UxTmU93jWD6kiKLPS+Z/turZVg+aVDVuGrzP/1pxE2CAKnEJwdCqM+ykQ45
kk+Vkbn+lHmLkI2p2Ol8ba91aeU1QQ7ja+TyQnEwwXagDDO/x75n9k1rgJhC+fxl0pkoOWd1ERma
N75yxrkhODuHarZNoLdduZ5LHFUpBWQJorEoJOXqqZJdPGc/fTTglKd2H/jLubhOig3zRWV6q8LE
M25bahMPCofpbcOUUkm8UYfwVUQepNcGwHwotU2e4nhW2HHvvNn0mqCMkrGFVU4lREcdqFpuoRRS
gWRnfDurFScpjOdOBkAyG4+FbBXqa+JCxKL+WscKZdaLh+utM2FbpKvr/vjuPPcCdcVB7Th0RswH
+/LFxqdsu8kfCDF16dkvGavxRHHxOPy22phjfgE8JjYxFhsX1vXw5XRi4EDL82nzk0xM8tG+mD0N
kjwyEcRCILrjKIY04PwKnYTPBb/v5GF+Nfs7vejXjvTH6Daq4Uw7iiMbRiOkYqze6/xAhTqYFGLm
UvCA4TLDkwFo3kIqEecQ7ug9Hcv6xfGeW7LyCAHq15EWmHDU2kRNWq6/yBxsMhlrwd6jtfJel71D
1OxYMOWO6NXFiD8+E2JG+fUMqhLu0DEEVY7K606vWBNrB1Fh7pKbxsN+bLebfLpCgKr9+xmZJJrW
StHKnqZhuhG2dcpJ+btlbUbnta3r6kevBaNoyR2Yzbe/1Eix63Lq3MgKluHpzbLw5R2lTCsA4g/n
INrKhOsSgJWe1UeI1htWx5jp862IK2YtdmouC9zFaK+1SHhUDfCwrSluWv4VgUm0fOTEF5sKBST5
I2fg47D2y5iZo7VXcdyrQ/HqldKIU2e4D9BjlLdUbipCYKs/9Ovpl3zYZznAj1Ot5SASZEXIV1HQ
HYuamvF+WPokO6MQZnEUBuwuanwQPUKDdaWKIX0OdePUdOhUUdIhqcGahXpfIUQmChRuR0dis9G/
vM6Herz+VTzz01jYBJ0ewpzgfU6NrIHNQdXXq9OWlLsNgj6L1FxbobppKpDQhN+t6iaSDuIgbiL9
RqAsU0Wq7iXD4jyWQ1TOqwuw+fD7Bdl5z2Byv1f8O75HuwdxLjeGedQAZ8xOOjssZAVf+kCWhFVP
co0ggAe40Nf2GG3kKGaXbFIKQhsNelwkGj5DoilXOaAvn/sSCVmxapugXqEsYTDHH276YJLX2wDL
xQQ9o0ewcs24HaI7SaeylDtDok2MEWwcMHUyJBeRsBowkdFhbnj7H4T9WRnUubORCN0g3fLu6PGz
1YlWfguHHKc4SgWW+2jNUPeJFcvZxjwRc5qNeWVgJuqc9QyDT3MLA2f7TYbOhbcfmL3y+oUnZPdX
ng05iSAkNq3JDYZxRdBmJSAlkHAdpO1s8w9HvOqJeM+q3wrgL9+xmpPO07Wu9RKMtBLSIBDlaozk
Ni080rlkGF+Nyos01nOyU8qc3gaek3RE//A7isg3L0JLtHWd5mUiBkEGtDPQsOmSk3YyiIXDhXcc
rYM2Cd8nmZBtxDpXLK9eUOqkanKs0E2GzTA8xd+kXMbEIrbQNyP0dI6A6Xl6dBXMNJPtXKb1uqfQ
IjjnRTtD8H7Lumz2cPttk2K8I8SWgiobnwDumR0SouhzwRpnFkiIdRnKpLX8aBREVfEhdkhIXMS+
g0gAFBmOpuiH80MGG7WwlJEhvGZN94eC/+ZqW8k6iuWmOyfoSroeacaRTm4xdBLCr+swKSeZblhD
enNEWvA7LobH2xy//6zKoSfMAjmPd3tlOkSc9SAafhAWrpQjGRbSr33D+Y2EdclRcQ7Y4IhIPYJ/
t2ID2I/CgGynmzNIwx5nTtt5ohohz7j1y78yQcT6dGpnpLZHTFj8Outz3bIWmhaHt2pYlOfoQFd4
w8SiYMxLeF0/raMG7bS1JMK6hHcIa3l8IARlDh4oR+tg2PpfAzJ50L1jA6N09BU/kBAS7AFRGcIq
TA0+Bo0zpasZ2IFBmw4KZrhJLHCNSoL+j7aCkUEgkim9az8VVSDkZe7RSbKaUUnyfJ5egWY50NYm
yuhXGgZ1t5/WLl41so3cpCGL+Wm/UBJydaYM9tNke6N+PgI0KpzeNzD0gVFMP/qpq3+nWq5aotsZ
AJGkby15a8dodYR4Vc6yxbfG5nuLcHnVNcVrEuGSNxx9MWUNhuMiAJJhOE5Bf9XqpXE+X5Ivjc9u
rPIcR9Ocs6mfVxmSxW/wLQHuf0YozhLtx1i57Dnm/5386tfTPUBlwbGlZsw6Oc1WoO6VY64vNTC1
JKyFAkzNVazELEWhRM/fgMSiC2OIl3AdHipGPQSXWvpuVdIEvOLrWJmsEh3wnUY2C/w+/5s/TFQ0
t54T4WW/29vE3n+gaXmyB82GRqMVlg3MyXRYUJJuxFOZA8iOm2JqeVo6gQ342txAze+dDYxPdX/x
DhanvG3Ml15xGFL33VTFyZqj5FhBC85Txq6PeYG67wepFvOpmFOIBAXkB9f7sWHWl0hVULnhQS5M
y6d7lQM2AjExwD1/YmDnCGiI/0oFgLMHIhW7JJKrtnwZ4RC0Xjg5JlH3N7VGEP9fkIrCcvwrU2GL
ZfXN5miCB/h8z74U/woQCvg7VwBxYVUWJNY3W5gvj2/iRp+3vFEHfJN3pgT/tmCvNrZALqiNZc/Q
u93KzjvxA2Lq1WAv/Z7ZGz1vTWwx/HmT3xgwlxZviJmcyhkhCcePjFfRV9VzjeA25AQ1EkDJJobB
Ru6Cn0mNVUIDNFfv966zfzeVknjXLIinKZNuxptaSRUy3hKmJlN5fbj+lfrEoLBnimzfLsNUF6yO
bHxXzJpYc2oTWSRAi2k83lVVs3K2Q1ifX6//Y3XcH0DMxLy0AmGd81YlyaJ3BZL62dTu3fGb3gXA
Dz/gx5LoNpgsVnK/r2Ny3xjNVGkNoyCzlKOOaKqH4mtRpD5Yb6SonKv650XlSCwpHCb7J9HVAXxQ
j4dPWfedQ7nfsUnWV4KPyalpNkvPw7DlRSo3T6AUAu8F3neeqRSq5DIvf8DlSwqSIS4y9pzO5MGI
3ohSZ7SxIZrD3U7ZjrIfpbhHP6J4EHFpf9XdUk+ogIMeDnSGH3z8Bq405vIvn452+3fF3anPRiRk
39cTBS2u9eF/fAqhKL+Q8QSK23iBQ5Bi7gN+iXGMyYQc+Bz5izcQHbeTvRAwiXBeVW1OaHsQlK4a
EPRuFFiQAgbkuNVtb5li61Pz/jBVZ69sfT6XbT/O0tBKsghPD7unTtnhVijldciG3m0Oohfk8iIe
ToIo8aODdh2OAfSkUlrpc9Lq0SsOmjuN0dU0J+o4gnQq7r2s46+c+C7LIqStGhmj+Jd1LjQMOlmk
RlojKMN9rLUf37zHSd6XY1PUWGpFz0Q1xlk7969MfhDtUZmF1zAKh/OTM1bq1q8KydhwmE8jKgsa
hQCbqjyr/5GY4Il4KP67MG0i51GkbfQjmasegKjAJhB/vou7Y03XgVAXG09hn4Rr5XGC8R60GabG
lO7wR9xcM5yKuXab54iJf5z6H5ugkw4UhRpJvbzxblYr6IDbR+MYbjZnA822B0ryirs6yAcO83jC
DKOEsvdPpyW9gHRV7tPFeYBeDq/VgbicqbYV3Bi6Tx0uW48KZL4wXNZKBLasdKUAbCZVK65Plsw/
kwR8YTwFfvEXPnpXved47tyY9Th5TNSzbNGVy2cZiQ14SBiAsQUP8hgoPIWUB5SkkidFuMJzqGuC
pDieie1KLzIh1wOtV6LANOOvbdbCt0D5qU3TYygMSLaQ9nQ2p4R6UdtJHF4+mRU6gUYrlMbYgEpf
8aVf1kQi4Bh9t3XH+xjIbslcf5FGcyz5jvu6hLZ5Dnz+vcFb4MI5qvx1DaaHtfjBLDj6kERmTUPn
kdK9waBnYHscwFSn1M6n65T0M9w+Oetd8yhUjpuhHRgkN/oJCvmK2Gu2UZn0+87h/G0/+EZ4mAxD
r48TOjljYXWnys2phaCI7gablNmw5+WI4HdZ3FxL64ZiyixeVb0VMyIwwJgyDVOr1kBSeduDtStt
+qHtwRPY1/bHfqPIHjpKSlGVqdzzihgUNx3rE26yPOuTDPQWCXGuYuRVqa0/tBD1MHaY2MwOGfCL
DjydOnUCKPlCLnm8obKezmW1TloobSME2n8jPSdsbMZyyFTDYe9Lx6yrNzcdIvYIWvgT7+paapPj
0YPrblgLBR8zWLsWCsXWV2nL/QDK+QXsmZ0kOY0pBN2HNqSUmw7YRHaHvmYZYlsUP2rQrx7Hl/q1
djdlUc5YkAL93o2tQZhUKqF5X0BCqcyqx3l4g5CNkVXqkVQeYCQe5AHVNRUZqwT713D9I5kBwsAN
fKMp7QSp10Al6SztCoEEqIEH+mCs+aOl2fDdDaoz26eRhyPyc0A26csIf+3xIr3QNur1kfwJdo5f
qQQ6noJFj2YbiDETVW9S/lu/4r9DBiZ5U4TEM7ZLpx1X8ezGo9qhxm9qD/Ca9pOI6Tvu8n5iqUua
7//C/FfBFkrKQobDoPIPDdCy5IPFKvi8LY6rodmRLAafoo4lq86kTpW/sQVBySRuzlmukhqa8o14
RBv510yOwqtGIkpeSDXDTD0aHmFN2I/SpdjLjj+gT0ZtURDeQ/n2FSTGahniAEc/LuJiem6fhHYi
ifEiuHn0liHKVMwG/BPBXtamhnhYYosVGct/G1jrc06OUkbaE1maB2/cAo5o/U5/MAOoRlrmLdjF
IT9+KJcAOMcLvqPQdGbP3H+72Y4mXkzoLyo458KaWj8vU/yb6mzPvcNBjFcx0id3mrySlKf2lEaJ
SMCkOuME/WcQZAKdFiHF7nVMG+YshIw6SXX5zqGjz4o008RLopJF8FOSZ0R+AQjfZvtFEfO8faso
2VG79CWu6u4jOY2p0TAu3j1YqXdSBI4M4psjRbpoZnH7Rj5McLg84mcFFquJBFiLmIxmWcLoeUsc
blhUQxz7gFFo1MNZ4waljUk+rhZwtLdcDZDUFkVcit39H4cFkSV5JiMzx9KT251MKKq0Vc9ZZDD9
IMo4b/gE5Qlu4grK71RB2DPYX76PmDAuMgenpEvlzJc+EOTQYjwh5VdcbT1DMaofqUeYeaYTmuI0
Bu7/pU6ky6LjgRMxpNEhV81XpLZfCpjtdhUMo9G6z8ILPIKA+O5FmNio31J96Rqw2LVtH8OZMfH2
BY6ANsUKksTUjuJIYquU3mp6yfZQhstO0LCKqdPCoAIA7jQOkX6v12o0jPUmu/Id07SVI56RgyzE
0Y1PKgq/tNyIlwMjJq2Uehjvb5Az7Eba+sPqv/1ZrpAZ8p5C4+ZBGxHq9ECXPqRfGpXcXEjdk78G
+TvX52GKI9JBHCz9JFQHsOHh8m5FCg4Wcx3i2RZFZhH+pwNaHkSBT3QvVitqWdYfiO9YjQBRaDrG
95w2nxEVUqH9MYQJ/Hqtket6gOXx/Od3VLQf8V4+5Fj11G+d89PrO/Yan65DzWPGjgFEHB1s2Orh
psk0w6H+6YkMGWzKRFa5YgRWRS+NJZjgZ6rWuYoE1zUShqfEJDu/uDsDVeGhgNQUKmVT/KbQwvB2
lZ1rrdeLHerCRth+r7wFnzQy8oiGaCSXDsw1VgH8IV8xgQLQds/HkWAb3lECSu/uT3HMHe90MMrr
1ATChUk8x/3B7wTO0GwHiKO2TAOHo72MPqwjhbkxQhgeGac2lrvXlF7rC21oDv5KkCl1LiJg5lVj
d2SYDSXGK+tWU2CWzhsE3T4g4ypl4Yuj5wBUoBhxLwj5qtWMRpd0+Yv7rgR251qfK2mAj57QwTtr
EnvN2mEiqpAnrvOoCqzMbqSijjUFRCdK1c9ksl53Ryj+yp++hxdm3EJTZlq5b5i1RBKtQEaFSjFv
77EzTSV+F6EpZIiXPnQb8ZqF8EDuYeYYq1xbE7201n/FXs/6wM0U1Atwq6Dke9Dv/DeHM+mqwbY2
ECEYprpf8qEzjiW0JTxAdwQwsbqPuvf0agHCWqHEwhbLLd9iA/cG6muRBFHp6AXkB6QSQghyBBt0
BoHzh/0bGZ5SPi7xqTRxOSSHMPHcDZqmwl7pruyYJL0wB1Rz2dLuZhcF1/BkFgmdDE7iORWrjoZT
MqkIlpUAGoRQTsDKGF1xk0HMm+Vl/NuKU39BK0nYpKIrgnXJYdhVt+zWssf4kEKfMm3T7ZIAtx/T
Qza9ZC5TK4Fa1gnL4DGsvFzlZxsSRb71IRPOnnQmqQq5SB585PRgA+fOVf/Ryv0xIzGPfFJJtcfz
4xpFqi5mQvTHMwAqHbyruV6WuJEw+MrfVkpOmmGQYem7bsnZkoCv5TZ3tXCD5zRhrskVnXcppVx7
SQIgghvxlgR7n6r0yfxEOGrLjq9osczVUbhA2T7U3tKqMacZycVTzlRe8Sc4yxTvZDFNreJT7IXn
7ojBIWdHdlu34F3ib/u38UfW7F+epgN/5U/HUD/DL5XbRRxejCwPi0vPbHA5I790Qjkr5AbtGTC5
71fcm4Kgi8f3bErpDgg5J3FL+O9CS08TIfzXevImcSUPFU2R1mplqv/9g/Ha7KA/1fFxhWLKmHOk
zGBEFdIqKjBgK8P0TJsf8jw5wvoGZ+E9XVdW45EDaYBzT1+/MrI2/89Gf/UnhCjLkkUn0Gol+3I4
5jPGvwHPtVgHPQ09OHesn1yxlw8yx5PhM6Nc8mnym00yPD+8IZnB97MBWfq+K+gagDkVpJBER7bM
cfvalFlMw4VBx8G5Kwo3qDPOZCKthc8L0KaxDeqtq2VPnRyDodRG7sAPqWXgX19tCw+39DEqK5D2
cgMtW46R4sNohW/GILZfYxTfChdKxf+pHKudKciu13sLa3asVMvk/ZewmuGKPE+kYQcwzAMBwK0w
LJcCJ5xHBxk725t5nIAkWOYVSRBfffNHJF12WKaUkUEJJMBVtptWSs3Zg6GpDSRz/0v3XrvokIQi
9aZGAo5/FygwCGPkaXztXT5n3H8r0j81kBMuF6FOvqkkYfBWLln0Ot7RS6zADOn37yTLjN8haZE/
ASpt9p7TAUI7pVUUGMkZYRFdFyDd1i7U/W6E606uuorz6uOv3+doU0eShcPLA6qnPyWT4v+1bZRs
34ZiiYCwf3TbSfPb/cvinAR8EX9SoJDvsAW9fBVBEECcytGnTZXaA71yAbO/D8k+4KXpFlisTSdx
Obhqfq4EO5ambou+GvK6VzxYRyw03ZP+p5F9DxS7pVR9/6qdn6ZXWI/ujMRWS0yh6lg0UPsEDuAV
qya8I637ajHfrt5AD2AjRsXUbifKu2G7QeIYL0Q6qQtAvs0ishFFZwNye0TT105AtQlP49ozS8Ns
ZzTLQq+YkI9n0P8n5I2esYz49zsaFGKa4cxPA+bOM8xjjYUbXxWackDIesZU9LpYA7VpxQU9cGFL
8yzf08aoKG5mN0nPymB5noiP34xTIBEXXcAsCyxCzRZTiJsHmloMbPOldP7OIS9rdB1WnqV3ePxw
RcrIxH4dJOOhraWDVcGMmPPoIHmAyUcwuuB7QvhCXg5rQnV6NqZqBbyAm0v25/u1pB4eKvz+yyOY
qw/hjMtKEXdZjjydR2/2qJpyQ+muNbd3IdF9rUvwZJwIV0HgL8VLAW2OnL01xc+TWgg61tgULnM4
C64sObOD2+GpEPFD03dtVWzXsKIyE2TQlL5KObAb1IjNnD57QErRSnSTtyjMajHIV0Q1i43gwIMz
IWmYAkwLjWP8wDWRuE9GndHCnzEuh84UGgRxX7sgjByHD95p721aBL2+6Ytx6qICGKFZxkGEnfi9
Mq7GtLJjkVRe+aaW4YiW85Q9cs52A0JVbErjOorUfk6kBrVsexXM6yMTt6AnQneAM/8n/5OAGemv
Oi+1AhWhY79xeys/Kl/8W51zbgnsLd8iG4gDO6rfmYbCWrPTufkvS3v9RuX2o8GhbZ3tFuPY0MdE
B0rR+3IBPqoLCbUOR0j7rvo3SAjbn0tJUGS8sHJq3b02el8MNX13FF11U2ZrSeCZtHFz4HZHfyrp
YljJkfEpqhE5EN1i8M+o0887CL78OWmS+zT58LZ5omkDLpGwk6Dg5WFvuoHaCh2svgm2dXP1FDOT
1iQO1CuXpiUNSP7jJp8SMzTE2r1uLpUMpHBGzToLL5OPBh5Vth2vXe8SH6MmGD+eNoeKXid/vXk3
nKoDGSsj/0SIkYxt5GJKyrot+vv1sHcXcBgVACM3zntIIYOOBcz9SXuUiRVrk8U9bc/3zj/2Mb3k
w2qzjseQhEDRmYNBqUPCGBgOWiErA9PJYexBnodYGZbEQSuH+ImxsX74Pd7xJwf+afuBRZ7E/Ehm
MZZiZcX7lDoRLZvjE8zuPnF/Z6NSGIfg0+YIBT8f53tX2DjttomAp8dYJs2EuASxQas5NhoMUSeE
XiAnwcogpxfAVjcHralKjW8I1+GntBltpx270Z0kzaYeo10SsTRKOM2M0XTyel1e15I6ZFDdOJFV
Dm4OBNN+5mYId6b+VlEenPfGMMuHrYzZqDKDC76QDwqOAdVlbcVGo7CUs0DjFZnsxGql6ITK91NU
JIAELmA1kn0Wipv/819mA3LujVhTKnRiP9AuyU+EA8lCFYx66XOiKNjepg3SoI3dr9BR7iESKWWf
6K4VzuzTwiTy1WGXE8GJyRWdGC4HFoRT7fIOGrlnoa4VYSD0jMDTtku2slPrcciT/nTYzDQ+K1Lx
hASk46q1MHXqB2Qp3JANbk5NdEOVlLgjpDi3SpWCs0g9kIfWvTv7VVB/XoypnzZwNoHc8L1ZgPmW
yYuml6wGa51Mv+fNPkF39VbSvDqmfCfN0hytXh4RuRNa+rXDazSgweoFL4UpTpMdPkkR4LvGv8ZC
+Kw1s+qz8K9KBIt2IRfnv+23j1IAbZ+9GH9fhSPlryKyvAIKw1FkjZuJL+iL2KH5nnkqEE5Jc12K
/RH0HJFw77YJG86ZXjhD1QE6ehLueK1gd4I/AC0Z9JACLhofgDFl3vxQIdHgTsY8Kg5Ak4N1sXPa
7DIGjddGQqOFiwLEcNKvFjnTl4DBQlNH3FEkx4Z3TWq/B7ViZMmgWISc331zL1rUQO54oixudU5C
57YP6ZNsy6MajUgN767cMXCB6Wu9+79qGRNLvHQgPTjJGSx28Xsoq+0R+acFPrAgiVuBBRQcIIlH
qLzc/IhNrBTsZ/a6NpGid7zo6IcKPBiTIKlhdQ1iGqrDkXC74TheH0IwvDWDgFRazMpsZIzbTNkv
KBkXTj/wO7PeA/OLzvdyLPyc2HJGMRPoeHr//QjbxsFPDssD0beiO6lrjPf2PizIxl+gjkgNjtxD
jKLKwq8Hj5/aGTbmCqHNIqYFT44xaLwtwXpCyan+qAw6dk7MmgvhVg7/f3rRFSL/FDUJLmNlMcbV
Arh8TVQBT15HZRz4BSDkw/EbQxLZi1nZj/h+ns8dIEtQHc4qhsNuazVZMkEbn/vWVTaVboWxGFny
6gAC/R1ygfZ4WwGKyw7qoay03nxzSBuiHATTzBrzoboor0srMH2a6/U5B7bdqOt0LLxoRdCCHQgO
ri7UDp17C2iUzfSx803eeghJCM+foXP4P3Bhlb33TglDmRVgoB2DK82OEKewdvZbXRndRRJHSdBi
hrUSNL72I8yaLE0B1ROFDA2j2glTno6EhEj/iCVuFOw2q0ytIuSMN3FxSIVkZBhsF2vxBZer5tYJ
rgkqX6GFHCICZ+guBxRwoN83lgfHYVSakzWACzOIaqgsMvxyDWq+dDFHhYEdnM02pPvZKsBruWX1
MXaPUpWXniYchTsx4oZiLViCkJ7hZhtVJql0NJD530RG0hcdjPM6AE9tH5E2wZZlSM2TAT0zHAu/
W2qVPZHpe+XaBZJJu48JdJZLd6eaYr6HVXZVqo6wJmegpioc6MoHAUp60xRpXsKSIP/2VgrLAv8t
H9CPnAy6jQEEIr9cxxyWDty8xoSwQB/+ZrhsQ12SoqwrBOoLrarPSyapIfpKtctLuJySg6d5yoRq
PNBkihhJT+UroCTKd77IsQ+ONuC0HW0ZTXPYVgD5RgqNQeQi9gXc20VNPC+lak3FNkzQ/jqd72C0
kkVbqVyEydxVVoG8NcYlpduoZ65+EDpV7Bh9o5+98oEOMONiMaNMP8tYxJPqDKjvTkXV9t90xfQe
mzxMFLZk81rdzNZoOPt6j6JSSUI1ebaIDewLwhT0u6w0kuAO+kMd34ihghwo/5wMF7cdaWlTnW2L
Qz/MpWfpHbvgFPxxfJS4E5GouiwteyaV9V+9YUXtHDgBpymCTHK50fsVWjAbKPtX1iNJRpj+hf3R
IXdLPV9mo5hJyC87wA5e0+JhHjWUIxw/zqefIn7ZuwHpYEZ2sBzom3tiauJzQ7kyCa5OAs2+N5X5
aLIVEkzD+AvlWIRmalBgpRGLltqbMuFcdnGhL1cTO0ctDaswzavdvJfOdtmdlLIvDayfhh0IMsFR
iLdUh5TypIJ5wbuCwWnYhClEvl/tYaudLqivtFwHvW/7z1KaGgZ5k9PW6Q3H1e3ZWFzAALhYLv9K
1+dihI7c/bog+KhWl8eYwGpPLjiOfGg6336J2H/QejS31X3FPinAHk9ylpCwNJNeycAXFM7oh9b4
x5vng8HpTZyhk/f9GB/fDbGSFpbGiVj3MrOrm7+/O7o5jSG8JVjBGz3uwywiRs+L1LHQd+dB37sb
EA3DtVAb7m15jnQYVkxnvM4FNF3/9iX2AP1+ZBRKvt0nF6+zqEMT2/XF4RkKzPxiKPGV1XMfmkyY
Kti/Tzv7SEE9hp5sj0WsKiNie0VcfSovpk2GE7qwbU3mH6PBd9AOId2DWpEWaoNKKq7kqQwPnTWJ
iErhV7PZhTB2qvEz56GYyfEfudquX9U+nNR9o/4fL5qlGtAAuN90ZLJ+u7V0PBi2dy+GENq1KvXk
h5JyX7y5FlWhDeKKej5ZZ0WvALZ8r+aTr8V06HUDC97MvjdoBr/qPaW3OOEh+f/VhXz093SQa0L2
6IcwaSil4dDo4aO8ktgSzDNjV6cOBxUDvVOiRwnoSJPYS7mtVf6bCasYM+PbZ+bDurMgtBxqi06Y
PHflIK4VMLY7+hpQ+iBMEz0BCzH5bXETZerf4V0o27YDh8f1hKzs8zj73QEUntg8oVXdbRPpTx56
QfO0eLCWEky1uYnKoceMzu69rcTiHVn+31ILLchjqyqbmfS5SMv7yFd4IRgdBdtlDFhKa7MWbL0Z
3dJ77hnAXWAln/iCTyo1UKs56JQ/R2MAsZZHJRC6Bs9jRZY56XRnmYfKzfdMKrSApFFCZVssMlOj
btOHMJ6Y0tl4X5Qp1vm3EzljezN4fphW2PMz9ygbzzmkjT609cktB0+Hhb+kP9FsNlNH6ESSzrsW
6RyPFiozV1JptzlDiVx602itWb8eHTvUdz9n8hbjZsfgehXSR++jU1w268Cp1OS/C8Dk+YDgkB1E
yqnrabvxMN9DlcT58oODS/eFcLNhPKkC94t1sfd1IBOauBJ5tLVSuvdkqMX9IwVhZu+secX4y7Os
FpHRHMNuxzDebgYO0SUOCuExAOy1RaAvebCU7bLFnxVxiLS9MIPwx5G9SOoUlSsBV+cpPbU7GD61
lxDXMgXGa63esw7VNEFT5oeOi92TWJ+NlEjg9NR55vt+gkthB7XK9GsLyT1EPKGNd4ePuxpsezgm
ISx/J5rbQ+QrA5HROZOKojfqqsRZNshFXfu638RAlO8ApqREIr8Fbu2SLcGIEO/631/kCiVRaDo/
L+T/9qUZUcw7Ej7LrbDre2/3g3RQS3EibX0tTDhdRQ1dfTMuLr06zW3op4dfsd9RZMASG7sjy9+p
SQ8B2w9PO8C+n0svGUW+1biIT9g1hIM8pdzVYQEz/KlEwmB3kfV+fZwtHPuNqWCHYhHiOOigxPE3
eIUQyuJAiX7oVdoKqbFjC+izlndDjQ9DJy7TyZazzsiILdQi3fkGYq5HfLVt2AuSI36bnF7LjIZ7
/dT4XSkHyrj7YtkEvxP/J469bBfqaRV6xXSORZbZp/AaiH3LFUbIS2NBKP1iqggZ3foQCp/1dw0t
H/SPcU9g9TTLdoxeHqq9/f2TtupHx8JZCquaNnEvGF/WQlC0oEWVTtygSkvyLj++4eDa6VugiExB
SRH7UnjcPWQ+dq4h81YtGtvX6pSpgIphG3o8V4m3DiiBYpGt7lVRA7DZnXh30lowjuPjGo/n92e8
3hzXBo6AiFNKousoMfnb8vbyuNN55XZKaoRYIuwfbxezZJk83pc4/w/t1c8kbxoyHv5bTe59uI1B
ZfvA/HuuR49t9lOvAfhPYoI4W+Fooq0JvRTNAeq64Xk4IRBDk6XY1Lw1Cc34+73u88IZtczoDi2w
Fli4R/xz5Z8Y9MUe/4PkfCLF7qqYp5kG1Si67+vZzImALBT0RJd4/FzjJiJmZ5w2hgEFO7+hdCFn
PP5H63lMEZzY/XFg+DGRgVMS9dy+GkcE2tZpX0tigf3agR38b1/+5AFONsv4dy8bqMpW9k0rV7+o
YWHz5dnRzYHXzMXnb3Kh/8inTPOeawFlGXmcXLOqSG43sOCB1sy0T79AXR/pMlHdPMFGTin5Dfx5
weMcY0MIvYgMth8kBh+kfRlZWz3oO8rtghwyCQLpRbIWy7eMJ4fAp4Z17t78K+IKvDD6W9kc3FHa
7UxfheWo9tZRkQS+rDqBL69WM05kl4u9nR09q8JZnS9D+RmBc3XAaiAausi0cTGvMUrukgw1jK7I
Ze0mm7q5iCzx9xfQLJpy6tSSa9gHmrkTsmKaCrfGWb48pxB7naib9GFCdBow35IxK04Fyb2ewjat
69w3211XHyskVnAcO32bLx9fIHIfRUxauERh/DhNmWRjZP24YNFejDioM3VUKX8hjYtkXRI3UBV2
llp0FRJYtSZyG0NBRx0C5wrElnz8OxzVYVav8I0HX2+0xV0MHNpph5tVX0NQhTnRr/x2w9ybiWwT
kgqTMv8yAb+NrmYcBfAEEoRc0bFMUccom6si1XyByPRX8iEUJXyCnqHGw39L+qZemP76/12ki/Fi
Jbgl7sUfsqgtD8GfhXvlhafKOGG97QBgI+TFRXs2u5w41UfHczBUwU1Kx8i16QGHm9Eu/IIjsDdu
saucS4BBrxuV+YYzcO90pzuvkL7+J9+1C1cRYS2SIwAstmgv0+Ep3QSdF/4/GeBX/kxR9iNoeRIV
BA7pdRSsz84c/8tZTLCz4jg2sDB5ScvQAvQTUlrl6S8Jv+RvHb0TLePYE3l7NqcAW10sB7g4Oyn8
Lhx9of8uW/vYotnAMJw6JzVsF2oOtMPWzh1yqihdSWRlClPNDIFK/k8qlMop7HJrCEK5rcBOQ+Ik
hVReNgZfvCcoJQibzB1HeeUVktKR9RompjbxiQIqP3+8YWpe5XmcmThMrFLHTf5T4DMvOXuVQNHK
32zct6UNOa8l4Rstlxhd4WoJzy32UtTD6KyQ/bdXVcSNjpjV1JRGFSNWtdK7/uwBXyq3vkR1auVs
S8yB+t/tIr+b7ShBn7CGsZCs+KHi7aH2iX6hwSXnqj6FHVnsxYN32igrGwWpxLBdpuhy6sOZkDjn
SW6YIKDwwGifb3jcf9UR0FqbA+Q8Noc+ajoAxWZLSqCJ13yUe+eCCKw0L1LzDWuO+dVT/IpJAahu
CrbC17EtvzuiayLUBnuXNcGQ+FKIx1BXtqSBLYBJbmZUeeCQaZdBP+RH3SPM40ZBcZtCfCrf8lZX
qrhgJxlS7zAw+kxXOfVmYPIAusvbcYJDWjui0HQeAj/KWAMDRJolqq1K3XcAu+W+WexvNQJZ+8QK
8Ke0Prf/bLldrrtZA0EbwXDk0EdgEAnNKdmEDbitxn045oeaa+dY1aoB2hmHn4gDRNhw3IFC9uN8
7m91fI/Gu58Zq6Pq3JGnCprdzI6mloKOiRSTwZxad5DH1rSFYRZY3jBCwpANRXZiVgx8KNcsBbLb
dfdhDoozhBU67A9MoFF/CEUHimI72/M5qAK0rdoDIvjkbHDXMEwdeQh8ce4YoBDi1zkeTDNVK138
j0f8m2CEzkoaa7fNEQQMar5Eic/HfuBcXDm3iLP/6ASGVVGN2CrRBk6rDtl8CyT1FYuEwuXdSRqK
cfaRoqvBLcYX/XKos0jbrz7fXdNm4fpm/ncHatBPn+vvEYo4+aUrdcaB1Icc8609HhbdC8Qt11Tx
Z7JYrSLJ3qukE1pzHn6KLjr5TMTlDHNsZbN0p4uWJcSE1kXU+uq9jgIl5e5tU7BAK9Y+CVKmAUjf
hn2vT+B672BJg5rMBZJQyCtinr/+TqX+3E8lUr9L76KO1N0C73e881jNBgD8yvCo+qBGZeYO/gUT
/8sr8o12E4E8fwmrh93vu3xunEe+G70OXHn09vPOah7oWiIoAmCWcWRpFwlX8fFBy5/9s6cegaFA
1HYriA3Mk0ogdYjJ5cIdVoFOyQ88aBxrRZxnF9R4FHGn9Hhxxs53LLxlOhKTnLa+/CQ48MrguF72
vboJ2BvQCSwAp+ZL0B0dxFNHGw53KyqFU7+c6C+Nd81kg1+/4CTPv3ecfJ2ZIOjYCCvWowJeSb+8
/WUWNfovKV3WVE3w08MGFy/2S8oxWuV0goPo24e41TsXgUpxR7h62e0W/suqqyi6n33J2Gar2GQ0
9+AjKbhCjj6HJeA8gciFA3m15XS+pnDOR+oY8PbQg+vqoe3vtf6omOkY5WMY9rAR229vWJnwBPZD
ix9MLOb5Jm6foyfDGVd0JtpwLLowFp8GHvyX7uwC6RczizXuxY1W5knxg5AjCQ64YL2Ti21PURyO
G7yuwdBg3bFWjIhUCzEbbSzXryiwuo/GnRyUwdgGgBOXpTswE4MtBK8W0np3JMa17/kbDaIVfy1j
ePrDcZL75/0oEMq5guRn8ah5slJjDRLc9n10wL4zPgftSPNXIXhisdDvQnmDqJPXRxK08A3QgSH5
8gowpbgCzhRegGUQQzz6BZklGipg1Wra0xvHjltjqHb0j3gl5k6XidnSbw5eLaPlfN8nVOxX2m0B
2/hXVUC7WSHVsaYN5rl+wiuKHgnwP9qIZaMpukMvirJs1t35Op9i4IpCpCv3ksMZqSgc1qf75uTs
BZn8WZiPQ2vUR3fijCLzhuxte13BnfCK5A7GL+aUYp1tmqS2Pc2GfWtw13qY/2GkdwBCqVv3H1oq
iRkzSesEyBBeH7e79ldh418B+9Fg5/jibyY06lGfaueQj8uITMDuhLm7yXpH/s/oqgbx3NMPGDD2
SpMiiyXZ4OeNR4oMtJoQGc6aQtdjqpMUQgtOQiwsHhvXWB/JUx9/Q36/aBNj/DRi6drQu5HuPZLq
mWKOioLa/INM+5Mih9TilKfLmB1JdwQBlbt9ffvhroCZXcGzd9VGtrli7oS1yJAqDTeEsRKMBvhh
grEB8WHe+W4Kx74QiY0qL0sJFzoLOka4gzL5d4sc6MNRz9y4761Wh2SBHP38Ji+NT6kUERs7Zwba
VfI4M4pNhhD7+alpAcKp2onEbAbSQupuBbj/K8u3u3hYpApgYRh6jL0ViiiL0RGVi47zYSA8ujW1
/IufNW0CX8eBoYlYOYTQcyGrQ/5DlUDSeMIZRGlPsBj1QM+ujGrYYzhhYUO2aiJd3ijY7WIxxubb
9ha6YSAFv2H3kvPJYCLZ23P9HIgRdTD+50QqjKmnes+jjuDDrf7S11SWW03N+Mn/JC2DkXEBb7oP
dKiabDrD35Qk8+LRoZp4UiY0pheNcrFWb3AfuCSiJdTe3ewhm3ILjJMWNcceLbSobmhnXYCgFEue
e0lglFhsDaKL2AYkfLnePdWhfU1o6ElEAMw0nNV8tEuPqRHeM5tTsJCLn3AdI6RhMbaT5WQ0Z/HA
/WVg6rRFpFhs+cT2P8DQk1YCu5UK33VAVXf5bN7vURKGmeV2b1/BhExybH5jo9aQSbU+dz+jEshC
gOlEJcGIkSYvFLvnyS1jUztQJaKqFZiZZQoabDVnAQcTegNbzcILAySKJ/wOYdcf/7klPh7Rz4+7
k3HxG1rlXaH29Rbr5FNRpvbMLDGXsFtZa4r/kgtvDJ392nCqA5ApX6qYnbJTWshGLavgjnZcbQYk
G0ryqJtbpduTN2Qr7GCrS8sH8a7Cdq6tPp3lNoh2N1iIIXj9sRT6X8B6Tto23jsZv0rKwMfk68Ow
xhH7K6BP2/DW/R8xKXTqXqce/kxVjF/CT4inc+hvp/9sHLztgXXl9TgZ4MOjJME1gaebxG/af2uH
hKVrJ7aorN6L0YAnq2ppU9FF9EgBs+m6SmqDj4NO/j120Oq5QgF9LF2kJaKMUSTyuHj45Q3ykwEu
jsJ07p1F86sHaG/0oHUdKqIDEcw0QYByLb11BnyLsL9UFKfUDXSgqSjNZND47gSgkyTh2mE5Ja9i
S689CDuxXPrD/pmtYCb4vGjdzXo+3EywuaYQLNZdOL61WxQtX/QmC86hK7+oOwfgEyV6tc61zgJy
DvNwhFRn1n5SFcJYcAgY/o1vDNQUpfdVaLiQ0Wzg4aoSbIcB3OrnjjPgCIBUK+1i+CEqSfk7rUqJ
DcF1k+fv8lThKBCN5/coX2gPmJOfyx0K969yaWX1aBo309fodwERD/MuM3ADqX6v5HBzYZf9VHMX
UFkqw7V2Rkw/Aeqo40fxl2psGJkoRUr/BtGIioWLpjBC9iLfTaO1KOehangs6sVYjDF/ExltMlb6
EdpcsWjtBezQD3m/f/4UAqfbeDy9goxIaeIi715lriMppFkKDnCog4f/l5Qlfrh1KCQimNZZ2p/G
0SBzmxszCbFk8MfG0qhwHd1navXyPzwNYYP1y8UrC0SHz4i4SmcInko1WkL38OWAojwazV4GC8Fx
WArs7ONnfSyQDpVbxnror+iCB3EiCix4JtyoccHTrgohQ6qCWxRQGfZ+/bFMLvG7fLsxaIU32usi
19mogYMr1xLPBnlF5+Vt5+5ccPPmouF5WgdHUH3boO0WkvX17AZDaByp2bJNMOMQqc7NfrTE4g/T
llJxLDadR6XMN3WV+xcP2Pi74rov0SJLtRhcZage/wLMDBcJvu7yAghB+QPw4xFdUzeiUj2CUIWe
4beXsd0IvJc09kLGv1F4d8FI67HCn+mFoTmkeifGXNRCFqETQpubtFRzjYo7mX+6HU7/i+rJGfcj
BMVYrU9rumRY9Wi1JiCgnYcMFTVA4OYdiUWWAKBtS1iF6gPPz/1fqlQykHeSCo3uJen5N5n3WQTU
CMq6jd+kMjHhGJiQ54lc02DB6ZUKrzrq1lJfASkwtG0cBp7hDxjRpClk00XaWqK1aNJ35QTVxok/
vlJo6KsPNY3G+qjJlASfqaJiPaZ6FPvDym7ADwKokEm6EY7byjcVAgUpM3FwU6HwxvOAtrznvTJb
bFVItAgGWKM8uErNt0rhv4s+9LPQtspX7E/tQJAxGcGZXnv57Qcb2Gn5a7JrbkYB9hEb8I3l9trq
fqzv40gVGaJXAn81rG1meRjuFZp7wvOeG/mHMtRGTpWKhZ7aU1RLbpSSRpI0s1FJj0/RVM1EYmmx
yY3xNcPAOskcTLJrxTLv/nwHhVNRZUZXnbc5B+YkSqnnndpyKPxrIRhH+Kt9NzUzBBrVyXKXOLD1
PK5Wm/awxWXrJfNwYCFSdDJlCmwkuy4JLvBDjxg4xPeXMeDnvLympJpt2ESTfCC8lCdB9qRNI7dt
l6MtVzUn9c53DBeVsAipRgdWfDqjPGUxB0DgIUs0l+bRxLg93RpPxeIUnI6MNX3chH6VMk7pVh8d
esDNwYO8E53M7a18tQr7gnzllvArs6yLdFANFEz5+SuPJCwzS6PVW7dtVKEmcAVP9s/AohjKkZjX
M1X8A5GSquiXX+GEmfICFuj4D8ac57Z7AGRhvE2WMfDdijuj8tWTevge4xZw3DKCKN/pMYMkN0qZ
1vQ0qG7e9qMU6y8dpHhug52kfy1/aVPY2hnhYTLAwaaG8JUU0OAWJS7VYxiw9mtRjZRG3wPImsBZ
xlGAOftQ9SCEAejrtGUM33pJu4IfkuVUZyf8+ENLhpIJQv37xtsTRrJAEGrhdacpRWe4PzsaPExA
EhuD84pZbQQ0jrEGHNS64oHzqSiMkciOMz9XCOBv4rRmVX3UXDz1xlXGLA3shPKOnV/YyizeJxuM
h0mWXAhrmm32EkIeQWITbuRKf8KLWg6mhB4naUuhAesQPAgQg5oBqRob0SogRr0LaZNbRqiQaJ5d
rOQzEx3fYnQYgiXFrrt+lzQohfGenHqX1uX4U7f/ClZaZBeYKj/CaIsYieSMaTPgRrjFNq6ZqLjM
ToZHUCIJj+w0fgjyEFukqdhuMQTAX4Ei6tRbAXRP8vKHzfLcu1VtWwiGzT0mxFzpNrmhHnBicK7n
7hCEgvXoLQUaE1TwdqOjbOnweOsWX/wv9xluNYxoj/iSBlEOLKlA2i0KeqVOkv93bwU2NzTnedh5
IHQDe+TGV+P2xtvkI/vzfqfL595rTdNFEaLA2bWa42rmiljVgz/KhtxbnJOHtMq2AcTFBiMeDJjj
j8iufoZ2RywxrWBB+mk26avIXgIZgCNV+/7Q7NC8ijUrk+kAxFZz+o48hMWmLh2pm0AgKH4LLq8+
+VD3arCGnbHZznq7jioze3kjGqzr5jM0KPrZXaZtnky9YtzMjk0Yw9QQ7Z6SqK7vTwHKpMD3LSWL
pxSV8ngXBgpB9b4os2moy7jSCPWwLIcdFLJJ5MPx/CyZ5YPRw00kyTsUQOD0cDw9Lq1cKYFBJtpU
oXkDBjKr5xIEW4ThB1k0wh1MD9XaDs2LpEoZc+kmDbDejGxkiwBLVEYNfWi82PTvhCFYhQPlpF2d
q5TcVeIZ9IsI1zcf7GU45O3gHEVu+WmwE2uR16oWhTCxa5YFCCC2Tqzb25BLQca192f0kUXMDjdL
g7Gj+kWAljsXTIpLSfoa1TbE4nqQM42kfs3DdH4vF/ic5gQ3muEW1wify4WOqcFewQfjWFRELaYL
g91FR92HJv1qUh0NtAN6twdHvl8rvXmE9ymU+sgkHjSuf6xikCIaCsRlDTUYyz7RKftnmLw7qftb
qbG/pFiGhYHOBeY78TsH0NKqrJHqd5Ljao5v8/pieV4n2zuOBP8GRvIQZgq47edR+9LoUFu8vmYy
mo+te1CmtZShCrDhVifgx88JfFMMbwsO0boLpYnQU3nf60tL4eMSStpLucXNhLzGMCoLEP+NSru/
HMMM2h4bWriQVIZNutyEyz3G3tUe4IHjRlIPmYbilcWviTJamEsjJLiTESchh+rtutai9Zp6ax6o
DuF8yz6T68b4vEA7YVAsALcsh2mv01y4jCxw/0ugbLuH0KzjGRJrtJaGZVr49nXu3dj5ZnwBke4h
ZAJE/HuoSRhwTKLSgNcIqk6GqOdbVgT2UrLwEvDBHU/hBH0dNNQGN0wQcXjnpFYTjfKUNr5NjqQN
QK0aGdQo+IEv487fj/VteIoHKcZ3eJFn1eM+2etbruPQFq90w9VIqaVpzcZ8xk3S8d8cqwhVEYCi
LFCCFrtJXdy0YzGAE8LIf/JJaN8+OhPmLxauOjEScYHPUpghVqu+wG4jcd/TGbcyT6N/jZ1YP/Hh
XwVy+d5z75cKJExLL4C2m99/ZmSfnDMfYDtKOFtdCAmDuQi+a2r0yZwSkGRnMmkWB8TNWrSWhhva
jFFnubhI12innesJAWCNPaLVlzVQrhcBD9kmLEb/taikVeLwmb9cwh9oIhcnoKt+p/cV/+3kkab0
MYUmN3myTVMWLCUswx5naXaESSFATHJsFlrUkmqR452+gKLU0yvXkQK8I3lUzPlV02lELVm3hKM3
IPWWaMNIj+O+qn1po8q8ANKA4rkxuLRIQwoJ1hwNU1pJWrsa7efBffwkEkbvN3RriBMsp27rK3it
G46PtAnEwhCwFDXn/AVdSlP+zU8IMTKST09cxGoqcLLjfm7ToSz4e+XAId3/yZNh/9QkBJQDquU9
kAErJto4f3iGXu2b938gToWHmdl0VEG127jfgLYnsn4WtdZJt7khafHZfHm1nXu32Dk2erTjry29
Xmr9cGPt9xHIdrgmHjz6IZGtoFEQp48uwO+xCEOUtAxwgk6LoKTIdUv27L9GwuR+gkmWdlfFmqgS
MZKmHzgnIieY9rKcU9anHgJKqllVNGkpNYMCcKQvfwm9C/jjTXkb+r/ntDJdPuUcX/y4vtkmFGGM
6ABk6DpPWScblW2sXWkAvWHwjz1uQohuKykO+zGB+I5J+LZAVOcZ9SXFrUUBa8U003mCT9S7sDMm
LufDEoPQ4630PY7BrUjT9F8FCgrWQfqgkJA94dzaHNqUNXxWuUpL9000cnEBWqeUu9ZAyhrKXr+B
oDBuXoVBbb1gbvos7VTBIST3lbqN/Jhz1Z46izIa9yN02N0+mpG1wKyXcDfxZ2l0ZAlNwdBDw3tz
q1U4BOXrXSM4Cz6anAcq0gK3NlCpDO+Cz32DUTzBNormDSBwcQLW9UEY7DiJibbhRPrjjHdhi3d8
wmhp8CNZv/1B3Lo4Ze4X0oc31DWI0XGyanylwsUvulxkcAFY6kD0hq+9B9len+aOWtQcjkMU2mh8
rVv8s/ajISWZvuDb13fAfBG/kwHLncv2HH02N5cGSuUAlw13KH1lbREJ+J8VGgbA6ytSCXFbN7We
Jz8DYVIapkgtz6KNkyl6IBzHKZjFo8/ZXTEYvEmkdL9S3/UBuUM4OaggkOxvl7JDRf6UdpxKpYEY
/MU6IrtUjSoDWOzijwM+HO/N50MJaznso/GHEdjsxC7L8J/lCzD2OkyBYRDHIVBoHoJczXggNc0q
eaXiYGq4tsfc8JsvSazk/R3lHKk2N01PtMz4fEs7m1XYcxiR6836ukPKY4j2sPedPkU+JJmNJt07
7cF9ZscAWEjdVsGeZYbvMehtnPoGEIR4oazaldvH1bmIK/E3oeo5m0hg3E60Y0VCJTFW7uUinam8
mlbbsRo2PAvHL38KbMrUsixWBucFStfzHSSgWpuAFGQ/PXa26WiFSx5Fd/bXgSLj0S89meiN8WLs
CC97bQk5HRqpBkM9XhTvMVv2hu7IofFQEmJOT2WKeokY2iuVs1q0IR18a2qRglTBmqBXxGLtY5D9
9MOZTuk5+7CtkCyKBrYg1wzXsRMSiV+fMaMJ2AXKpa2XdnsL7uOVwXDDAczgTKxzuWOllHfBnfXH
c2Yxr7+xQMhCwLkC5gi6L6GWDn0hdUO9KSyQjIZ/CxMy1qTcV3KGFC8WqNr6l8zyLIPmr+GKqYv4
y71Qjd4zIvL7hk2q2lxqrnUk2G1UeMPTfboLYM4pT1RaRkbWxoEZfByMvnWpvaiA/H9sLB1TWp7Z
UDiZUQ+l7Q79hdkz86p7RCRIXkRZ6Do8pPJqI++2baLnMgaAetcMzpS2GjkGwqIvsVE/3H/9LHo/
01yBD8/GKYvGs/EIQX3xDziyI6ywjkaA09N8EwG/Z35HWL8yAFZP4jOblQS8KgA/noRRNJu0qrFE
LUAIvwDODuZsa6H5fODk8u3NgYO02+LFY60db0wcugHjVfgPZr+c9YYAEkaNNJdX6+rUF9Z6DapF
tMnP+PRpkttOv7ngDaw1cq/h+06eI0XwCLBtzduFu1ecjsbHUwsACnSOGerLE2xly+/0z9r65mJ7
JRpcRfyMEPiZwvMeN5APYafedUdXZs7gn2RM6SHoEiVUdRoo6UfYuxK1pve7JtjgdSXcBN3HnFiQ
7xIybkRGJk89YzrEvVgUsWO5Ae2aWgx9YbaelhwsMfXmWPTIJlKDKCAmjnnEV5Bq10Zv0fDsoDQr
OKZ300ApIBpXKL4kWyULJjccSoi2DhWxXPK6C17jLRHfZyHAYA7fe7BlwzxBOW94IP87Ucibb7r2
Ntj6EL+ZaDRHaFVIDxdSpWv2+ZoWqDT7+Lm9RJGmgwcecRvFIRE1bmRcsQ3Xss5YK24tafIc+1Qn
mzFRGfMEKmYgVQHnvlhtVxm9AwqgFVBYhy//KsR7MdERNkl08dVHpAQjyTidUmWLLUkhVq+B7LBB
La4zdP67qvUReFZDTZcfC/LxnNg7WLEsusZ19ZCvZYrUFi0YJQlMjqJkJaqnZP3Y5j/oV1rZyCMU
Q6PtTRrabfKlRvJBS4dJTjFsxj1S/TLLCsPtIUtM+ukMhuXWaC63B7J+xiw7HcCdJ5j4mRLgGNcv
tSa5glsH0WkTQl2n24x2zerjEzV2pikG4Bh51bUDTd27Pn/OCU+mufUo+5Q93+0pOO1ZanUKKLNa
9LB3emxmBq2rQVCwLCOc861W9BwPzGQMrdmcT0UajUjZZ/fG3fs2+HxYvrocS9fDH/hOeEMq32p2
OImL65DDcEJvabFseyVdJCvb/aRduDH455jX4vIO+SGgaqc5+1DsIB785EEIFGvmALZIbVcShuv9
+U6YQzujjed7kny7AprQ7xR2K5DmiqUzDv31IWgC5uCAZvlZLZ6WjWaWFFhd3NocwTaDrfoeLsEE
QVRn5RRtQE4dLjOf8C93qs93yfvmJclUylGhSJezZlhS9kEhArsSDIX3+jlKXuKZVlHtYjqCI7CU
WTdE9xC1RPDTP4jIbN0H6rJRpUxrnsfktEnyIhDXlIV4eX9pUnXv5TS5SaHOd3acLnZuBy1hTLwc
Zuo5+yx6/7R38MFPPQB/3XO5QOqbe/JUUi8GUjZ/A/7BJQ7wvAKU87X2aRbSLT+pIOn1WtdWtAl3
Q/0WvKBLX+IFY7mGHhX6VmTmTb4/uVJhoD4sH7UlqgnCElJZO9E0EWP5kQMWCLcwgLT5qcE7tJqz
scmaQa/ZC7k0HFFoMO/oq7YiAek0+IDkLSmRtGBeygA8T8EUuNmFaglYyP4wZql3X/DhnsA/bgQ+
NeuOMnqBGh299EBY1UvAusfkHVSQTI1h8mV3IvnBocYwbKjznVq4qe/AUVm0PKeAsIiwCim82Cdz
9u32+gOB5KVVWuUozH3x9lqgHYe1lc4lbK8/Uh4qJrYCwkBax1AIFa+vIahLhQJUxGAMBqGF7iww
hS3Te5/4teE794HHQczSArCvh3sjkxcwQ/M7Zw2gqH16Ksq+OG9+HBqFBhRThzeJ/wYblnlgz3pM
7T0hGkCUyfAV7us3E5skbSVuOpgXs6LgnJe6k0LSrnW2N7GxfsIGku5Xwk5yA1Td3kjY3ThGab5y
srfZTTdrgb4pQnR+sP8zDatgK0rIf3WqPEqlCjz3kPBFo1qUfKHXpZdKb7oXeKKy9zbFz58ihfae
FMbIc+7xD/iazBTeiRs0EMZ1BAW1uLkHG9BmdoLwIs0x8vV70K/hP4KcmwjuQW9uwB+mDnn/ofJ9
tkY4zccgY2XL/6022rE7dtx1OxN4L9/4m5fwiXvAfi6Z4x5ZES2j1rRy0/ywek3+PMni5bTWd3yO
9S/ZSKzAYH1/vQ9XR8FD+YdGj9EZlD/GPsvJXVgDH3a0ph8ynjzrjTHNIKtTFoXOjn6nfCzJBM5R
7dV7BUDL92JN/ujfkeaqy+dcmiMMNuZZ2dRJtiF8a35VDx8PEaS1QC+jDmTggtXmx0qagchwtrhg
geEsVFzuzcmJKL7eE0/7qcIJZegYeMOzpyHG7nXfHMnFxyPNaRfLEgjRRE9dZ4ZF8c3HWp3weWfa
j4hulp7ObsZZvohlDuoqXI2bK4dmAgoQLEZq0nLSLAEENUkKsrR3blYgT1AyobLfk25rsunGnOEv
/3hoX3nm4tB6RDCeOPB+zNWGs7OoH8alP4PdYmkuFH9rdtHxGl99Ir2nRxagcFA8l1erIRMytZE8
zokN3508Y4IACXs/aOlH6D2isTupwzbkeo+NWEb2jyBgx4RMGp0SM4zNr04DWJWIoKNj4+YbYs0I
oX61TI9973E9ISctjOX2kQMWzjGDgBFD6IVhbzdLzlJx6G6PIo8OzD4yBTzugERC7KeiyEr6NmBA
AIBUwXcMCNrVNBqyou542XZhJDzz3UGR/ZNws9d503XvhjmWd2Qs25P6cSFPCTNrqTyyf4PtaooE
rJbZ0zFI/INHvP1OEwT18/hcYFo043SKeYEMLGeH5aUr6pyX122q0zPObV86Dj+fLXXY0RfZ67bJ
+58e253d417RNWXjPuQIVKrjhIC3Tvd47fcSSs02HGJnNDzbm40IVcegbKySa7dHEdWZT3VVM74B
zxfKn6p8JSzbBJ86uXGoRPLKs8MFW0vbb6N3hFpBnojwkIRF8XHUmYV3hPwRdkYk1V0fBoroPgWG
SvmBKWwT5DAZjsUK3k3BcaC/fokugv1y7ZV9lofz6zm8V/mq8XuuVqgpjLvCyC139b16jPxbcHwu
jHhWStNIR+61eKkchDRyIqyFLOE1lm6PCaCuL12A6fHtmi3YY2THQ8TWJoDEpHTTa5SXoOMzUjoe
EhrFB+vihnuZqunox8qPvSFwzzrS+2ZeYvPp62DGzjJk4NmrXa7e/PiisBam60E7p8ggFSYmb1uM
0zgicqowNIap2XIn7nhGyI5+g5o9tK4kfqEnlppQhPcoN57R4JQgdrL00g6GN74xXgnCKFKwpKak
JHTUfeyE91oM2VfEUAyZvU7+eT9dFzuYzYW0XZsQfdIF2gNfexZOEuOFbLIqXrzDARtDtWJd86Q6
ChBtJxjAY2LirBcbAQPmStNRK4rclCTpqJUPuipCNw8NizimQMOdwJGxmem7FrrJDIjbWPkmfqfp
zdEckc5cGwIm/BjccFN1NwGam17t+JTV0v2Ehg0jNEWYMQ8CYScGP+UmSeC+LwZgvHXYtUvjYmvD
zr2k++RufrYha90M1687TSephHKNhFxCFSEZ5kOAxsv4acs6Qc4Ud4du93yE9KOTcQ3Mn6NWLCQZ
YwMlKlpH9rNRV7qU1CWL0+vEqkXEAy1Ti0lf6L4rIkqC2U+x4r5ochklaGDbPJyhOwNrR5Ls0Gt/
dPAwtKbzjNX/O9ZVidzj4LagLM5Ituk7wHulBNPBVFK3xv/JKuPkzXfXaQ+VjDnQqY5lwW0Jz7E/
PUZiZq0Xkon0LFjP3LogjtHrlaCdu9/fhOA9FxqLawQtX2b0+5+S0L3TsfwQY188xRRDfoA5nWMq
ImJqSmrCnJGSBX8xLhaujJqWj9xnqwp0wvx0y0wJbfOtD9aHZMdbShBkS/6CxlamG6z488cQdZAW
nqWe3eH48LC+31YHl41nMkcTLvoENFKqHAXJzUZOsvp9EuGm+/RUkgWoEgXbY22VW/hcaZyaoYPU
iAHamGESpPNnEg3siM3wHfXs7wZTf7yGNoX038pLgEm5xiCsODj1VjmmhHcfq9LjR3MvHKV+LwSP
LWtrqFD33EYoEQTfXzLVTYQAJDlB1VAL1R5vHqaFOz+/tUovix1EGdr8qao+d+A83ICMr8E/BCHF
Gtub8AyQ3mEnH7zxBesGOuyrE9MxMt6/zTupDE0a49zC64e4XcH7o8IBoTODxV9GypjeYmw8Llbm
0UZubLB0TsIHTqljk7roDdjMlcjBrqAXxhaf37db7cIDSw7KrltmfjKjbZvJav1jgVZOm/JRg8bg
XtCgw1L7qlAvGm9jj4oe/z7QeHhJdzDqpLXVOM3TTpo1CM92F772ILDRVsmDj9H4i7uZND1Ie1dX
Qriw4bGxTOO1rwpXvF3vrGRQiX3CzQIplTHlYVa5qpJkkq7OMq7yN6y9SUH+r95sp4QUuhcLQQy3
cGRrpSL54z5DiqHYhA3x1n2hPS2bFsKQjmQLi4n5KZDFyKPM4HJ9S1arq9cGPbckEukuv1sFhy7o
KI0XvEONKsXFvWO6OVYT4rQaiT3lnMopRytnAUzfXCzPXFm/aKs8NG85dOUX7nujLYqiIg7MEBHo
1Y9KomQsUC5Jdhq1fi2wnWjDfDW52sZAAp+/B/fSjqwzQugEU4ndJOi5sPhnC2pcKX6HMS1t67aJ
4adkL/n6It9//xWxjzdiQ5bbQCCwYRnU60TW8jE5RFYrthXtVCdmPahSC+wps27caRLOGrPeDFOk
ZZt6lEEBL7cd1rvxUD6L5XYezd36jlUu/ZgcPDbo5UL1hJRu932/+yrqUlrHJ/uweE6lon2izyq6
6frRca8YW/Senu5gRhsn2dXfHw+cRfast7+AZSPRavLj2VDv1Aeszn6pAEfZT9Il5yw0+ik0IL/8
nYf++lx9jJE0mCBEROdCsorox2DF4V6bzDU1Yx3212BMGAjx2zUESSSVWUkNpFMk42ITheiY5Ffa
H7LaQeYiH2WJlc3TRJLmZtVISVOtBqbCjkwrY/QvAWocnuRHQwPslXq8KcwXg1NQHszdtX/nzhgB
Zk1nBKeuomY1YscksMiPcOrBAVSyiLEQbHIZ49nreEqP8Xx4/Vjf7vBCvRstV8yod0eO/5P97mA7
VQAlxXvG0JOOO4CL+3DLgdf0ZFnBJzpOgtPSg3JXKgvM8IhXnWBnjy8RFo3O1crNKJfT48zmOz02
Js9NIWR/HAx9yd2C/EtyIbaAFeINMj0+vda8u65xqSbha8O20mC9hhJ2kvwsxJvMOeAVDQrPgilB
uq31pRtYCLFodkroAnqAvzgCo3CKgGPeU2J1lQxu2vyM8JKBhQC4EAJif9IusN6RRptY+fZm7d9v
fxhzJzpwNWdtwm8txbaAxkNVKZw+YQyV0MNicyliRmX9yah7IZU8bA+0eUiQZ0wfc/Po7IV1WOvv
Tdi+4iPh0hI6pFNxmMMmf8VdUScREjdW3M3vIcWjoz3czRKQCh5TrplLLpD2Lf3eFO0z7Pyd1+WZ
55oa+njFXWNABkkRrf1AuVdNMtaTsu5FOjtW59WXuJ78lGYmObnamuSb5f0l4smqk+hgoNjjRgVL
KTAoP7VQoWp6Vl3knQ5Eq/HobXUTvU9A94tbha1DGguKRZZTVegnep2jUvgJl+AhA52h11kTDu1o
YMXBt8ACYP6wX4m2FxaFVgO+LNDYT1jPoz3NPwK6y96HZ8AhhhV65Xd+TG41jEfXogxndM/8uAjk
iDpzLWzOFFeO3DLWvQs6bryOo57JPQaZPFYoPBsRknEk833q6dRdV3iY36BntIvajfmCYeVsIGw9
HzWHUNwWGzixuCNGM+tagVHf8RfPihJmgAJNK+Qcx88dxXYjZ3a/AmBKVhEN5xeLBuD/kxYiCBok
NwEO84ElVN2vTZaawYipYkcw5QX2lb/IHJj/sPwW+jnbM+8Lr83CBgv4WnDfY+AKn9c6JGTH0HgF
m5dMHi566JSXqhN2kamso82deXi5GIZwBmT5Y/g4PF4cVuiQbMnHimdS8Qua1yTTN2pYElNubKLb
c9CLqHIh0xIXhh/IXp2Oh4KhZR0pyKhgehyU7ZSUWMi+SOD+PQxU94fwOHfj809YQKXzjTl7kBfU
YD2/8Js/LeE3YqFjf4yOmsV7G7F8WXCxG7Njjl/Y59H+fkr4WRtwZMMGsJRIRoCQMwSofzq9P/C6
Awqrdi4rKj88qwqOOyygSOGbO8AClmMBOhoJPYJag2srIg4bqvSottxNjJL7809yXFNiXkADlYXC
HNBlpeU8z1xHC32nBEzSqZn17Ei41I1pvJh30IpTkNnNktg0wwifhVPIpCuD1qD9NDxhPtDYV+mA
V6tGfXoknKOy7TNmewE2a7eU4RZKQhIrrHC5lpmysyqQVGmGs/DIGrz7S7BRZWBAWxDPNSgGEeow
30+xvjaUQVJNSzaEDjJbNLzOI/zu1as6TmaXmoDPRv8dL+gpFqxaxMZUGUE4XHlqBTjPr1oHkzR+
9aews5pSU0grEcD/evwN1kiih4jTdNy4qS8+QWwylOClmVUPpmL8NNHcn5EpYGPUZDtpuMXypVLI
xAz7Rkozsgg0wH0APPvr5ygsI8CZoJrqLZA53UlWWtfLhmOdF8UiWh+4y8BAu/u/ly21rVYNZm8L
yT8XnCDmIejQ+nbY3msGIzDJSh7lnZluKPf8x+p2l117duqCTb0ekegUK/n1dv9s5oyvAjTkzzvI
/X+T9bewxNEIV5KLsYYOQ6nLEbk+NZNXL2S+U8fn27HL03nQHOWkoDsKvFSObBMllz7LcrOl4Ceu
0Eh49/AYtqlmqHcyR0C9iw5v8wq7Gfb/jRASWmUt4ABCR4nVWuVUYnjYEqhI3LMmZ7xyRzJWF7tp
Ogu13o8Kv6LojQdORr0so/UzKKTnPWR8bTExKi7mUTpAgo0EObxmqupYYpcJ6LXMbi5+IU6LqVJ+
B2g0D5DBbUorFtmsajuw/tVstDioHcEeJ1erS/A2GRt+nlBovMnEOgQn0x8QC8OgiunkqWnepiVF
apjB42HxbDtVsGISGMCbrOs0TSjYxG0tKnaAFIstX7RD1KM9jjZZxR+GafGK2CUsNC9M/3CHBBlV
yeyF5AFeLBFZl7+++9ZS4pGz++kA2kpVUVbOichMWW51E7zdy7oscnD55jPfpXxVQNEY10HwhrZf
s1otHDpiM+GYUxUcKy3LkyJhPuO0xqZEBvuERfNrTlG4CNsvkJ732x+NQ22DVF7LU22+wRiIAOsk
21VlH5RSusImgeKuNxz9ef9dMUGtcTdRSi1+oLOCmLvkM78ZvPvmbu+9APxaoAXsrqkV62GD6aEU
GpoJX9LsbrLZrtamDEBoQYo1xnwq1A25A4Y4+uKOJDVEXsjAiio47+p3bgqN/P+GxPkk6ppeyno8
egYoSboH8ewfP6WXP8qcCsIOOi57BEOhcCMyvEilIa0Qtk2FuXfr8qpd+FE0TGdDhEj2BdksDXa6
xq/pk3Dm+uXEAGeNd8jHzSnQZP00V+P9YCM5Goe75zDXF83DqwPAZXPOEBD3i5t9Q+USxHDE7wDh
Iv5eaYYnL9YYRM/nwd9OqmvwzXo8w+9OS3DHdfF2CtszPeYNXeH6uqt5PV7dYbMnkA/AuuKKs2J6
MG1etgdWaRSAyMTI9JK8ZxWbSMWRuyg32x94cbZi0IksVBvQz4t8SIyzY5SS9Dpu0qJeNJun85yl
4Rjq722E21pMIrmzOSeo3nCcvtsBu8YxcQLppvgrU+2qjyPf31BTi/8x+w5rmdi6cFinnhz+UepS
ZrJlVBS3KNb+UISm/doAKLdUXFzIKZgCxl9/XYPWVrtqlG9EBAz7u55r+6vdeRbkRHjMmE1sL292
9AtYCMvSDgL450vbiJkm/UYKjqQynjWiJ7+9lTaaCc0pNqGebUi05FStO4tZ+RdTG+dS7df4KpaH
YRklBy4sER6nosjX9FUgxCa/As7n5ATUHgPLX5hqlopS0DncL8OA/N1sthacIm8GZgKWVuUs2asO
AzklkC2h8QxuxdDHItO+a1xcAlW9ntyvTtUM0zyc4Q+atvFcbdvtaAECCLL0vqZr1tN0vcFmhbfj
O3SI1mvFkw4tFQzpGGS12VvlSJ5Xh2wFeStniB5tNbVphFw6diBxrl1IEXrDW/u48Lh0e9AcQK8R
HuypZlJPdEWSh4p0y5KDL36E2xr34VJCgURXqcjjBfnqMyKQ9V9UT+ptIlJsABR66WkP4aN0ufwU
e8rpTBjHRSVIAJ1FSVE5i62qT6Q17KiFQSgn8QlMfp3fEBdGK6E/dL31wIgcaK9zqWuavYmpNq87
xkArfFGNKPVhXK+kOlE3M5WzPf4IyCMDPRhDeMdxpOu1e0JxdUjn0oGxGTLXaaJFfhRrGHCY+A1L
1F03T+cKl46KgDnWHj4gscz1xzIsjSiCM76DxFujpAgoS1GbbPyfJdrD7GCUXaCdk0mXn7wwyulv
cCnkQbdnw7VwhGFUa0GsFM1C++IAuzwp0kD+bDzDApNxc/hPgD5uV0fMnU3bwwJPquaMfg03igH1
coMPX/a5DwlryyRSu9H02tf0H2balZIn4AbU4xsovrIngax8ZGBWyfT5Tq7XDhb983/RitidAmpf
dxC9OnZChtmjkxDkQ/yt4Z/fGf2gjeMEDk2UAB7v+q+fr51OcgNULwxhg3kqJvSD7b11hFKX8NYV
35FTH/1pr0NhWit3tK9QM6qcplw+FaMntybmLLjKwjJXLAwc4QjTk2LMKUxKlES5rLIVmfGT2T/2
hb/7xdaBmEtQxTUbi91o770u/SUKJoGqQLukGF/uj7UMSduR0enB0GTQmeh9xtwl+fMWcwRQIL2r
CcP1KJlZI3mDawnzSEOCV1VEkGfw+r4SlWRZ8CWLS4o8uGGq0+gtNrlGmUqlateMkQ1EkvppH41D
UK5Qs87w82dsLzt5jD9iPAIcfeQPFmdvgi8pzIOSnVogwc4bVNkQaNLYY5m9lqBRHlYp844yRUWR
+sOTB2yKEi6zyqLNOgyeExNzOyPxhAuERQeq9YynO//TfNBI+XZIm/ZHBflmIBuEpnXZn9G7buEY
bNEBpS5qJgdJSQjTKMrHvzUyR27dnjqgH8SUH6q4F6JugMJKpf/yQ3tCXF575HdqckOby/L4wJcs
0KV5VvtSa+pl5mxFVGrw2LCnjLE+kd9t0hHD+JkKaDfrrituk6W7GKe4acmGWqdPvt1b9A+JepMb
cBKr9InKOiBdXvPXN9hq9pcmxHkQiqt6iw8acP5ZKADKEV0gi7eUgFSdGAug84kYMP2vKclzQQK+
MKzNIUar2qBNTPbGCeTO+hdlNEleUS7a+fzpP1eGCtopuvlpFT20X47xuFRiRMpR8doKmfVxEmTX
aOEwcpDPelkBwbwE4Zu/EQlmIxS4Z+jbccA3LcwFCFenyvnn5kO51wS1VU0W06EXQQcsPmwCcNVX
PeEjb5WNRoKzYBj8+OvyckJVIcUYpJdoNCmmsHe2y3v/lP7LTzAxTJhkzMSrbXk1E8JXwZZvwEc/
PnFgFiu3XiKL+ESXBPfRWWpPKr8ViX4amWmt3ftbQOUhihAksnx+BuuFncfpMZ9SuBmhvqK9C1/5
SYFWPJmaICGHqcuCX9vmTSBLs+d+ZiXrt0lx7mxE+vfaCKSlZlE842BTR6ZBaMIFWO6X3wog/Gam
guvpmuWPNizHYb72GRPt9mxuUp+a2WBEut7V1CIN2GmhWpw26wiL/Q6MnYP3uf6ymUWtEb2IXKli
m96NWy3QqMOQz2ovwvUsg19bBXD08EubLlAPi111IFxN4LDL84dzV/7+eSdIeJGGPUmnsja1iejv
q1TtLwC4PgQGmNTEpqLEiyQLpJQwTvxqjHsElzKD7uMV5du9aWNEzBiKETI90qXDZMHMhrLh8Fe0
b0+WSfzj+KSv1SADuuKIBwi0z28MUfG+hK5t6f8c0Z9ORk9LZFPCkEmQGL/QD1S24JclJMQfcs5Z
xUc6Cv0ICb8KvokwOQ54UA1MNSKxad6EoPlF67wHJj3/6mUYCdBLiUha2ZmbE50EBXmbY2egvFRo
m/Di2QAVb/Pczic2CQ2nSG9TtprhgFFLh69JWXqoY/no90lVQ8PjNK0TJIpO9r3FrsLGbre0k2wb
XWD9ea21AdinWMpPQh4i0EESMijvcsiiz9g2kHvmeuu+NbVSHrpBZjcS851BIJ/U6QZarfwsRU44
uRVmLas+kS9DfVMe/0+uM2q7kwfqeWh3Ok11gzAGDngEn8QS0beMvYELiK4CniPJ4+tT3fU3tdZU
bvXuBxXEN7L0+ux8+bC/yxAibC0npLcHzhfcDd9gTUHAJ6JoTvnx3DjTOM7XWudB13Ar2QBAmHLf
RHXMipZbcWATr0TVmbpyH1JPsYt9gx7s/eR0c92YNCAHDaHIGry+jAfYhy3VpL8Olnbw5oPGbq/A
nQe7bPUJaJYDUILVM9c/lrSQcinuYpDO2JAZoeShG/eaqziQfj4F3NzX9FgXYmjpFDaPs2A9uzPR
fzNdzLoS9mDhqyZJvWksugGw4O0aenh0J6ANHOyfu+Ndq2OWyJuwxge3Lb7QcC0W+pBvK20W8RrW
9sHfhXazvHV6AD9iOnN2fgP6sN7/62lydxuH3HkXIQd5lJf/0/umSE6Daz00NIrr/yLoQKUcgcJL
JRxiGZz+MZYzCdl96ECwO17cX6/dKJSTzc5jgBLdfIjUgdOzDpwAuRFxnEUsyqbcXol2swrK1tUq
0hggyhMcAS6o2cVybT6yY4BxpSKtrUE41U+2wQhIbtMha1TTcIRBNKW4aAW+WDA6BiAKC+kDGuX0
fHCcONi82cCGeM39vayoM3rqbn97UdVaIXxGQdjBhq74yPkffB9BzSa/cDGvB0oFIU2f+hIC+Kfw
1+HknHC4KhwhgsyxixDcjZ5B2MVk708mxiUC250TDtfIz0ZOsRYMoCYz+pgXXa2jk5aWmtkU3Q6y
6ufsV5zXuhC+6xWLiybDTXoyzVCO8xCQLo8UVbt9r2OeghJyh83Lm/MSZkqdSRS/3MCVoXRFAvk0
wJMbS7uNjJwKEOMrtejOKbLYGVS2Is/iY33ddd/EtaYgBKOww9Ble/DmnCPix0N5e0zVbyoLU3/o
4FsSCvE3Xfht58W7xJSV+mBnJYwhRGoP/wqhS5nIXh1qb7QaMsYUDdyfyBHubzYx0eY1UXxpHKwn
9BL72imLpAECdSd43Qe6EISvuFWESTwDdhKcI1R+ZVmIp2BpD7q4HD22BaULdiJ6t6E26bSqRfIK
Gk0cAhcZO8f1RDHVU370w/W0ef3My0dCQTyBTnx2dyvCa39eqY/YG0APNQfjoGxGGvbGMlk0G4Ea
CcGffz49pjw3RC1GdTqpBBtEyHh0TDzW3VQ7oroCIfitV5/TKXL34PIVu0jzJ0jpLn838/rCKlnD
DQJf0P60W5ar1Pelb9k3Thi9GilUvjd+xpR6muT1lLHR5Rcpegufg1mUFfJ3K8ZryhbQpHzA9MB9
QXEEPjzWjnkKxs43WQaaPEK6KM7DaRjROYi5J3WNS9qyBl8/pOnAsqEVIeKrROkX0hV7focbeH0y
Cj9HhxPGHuIxYA8bXiLYK2sD6jVorMdiMk+R5Ux5e7ws6v1SzOPYqHawPICtbdIsqS3GnprGVVaO
Is5Cpou1t5iSDkP+UMnR1j7G+JKVVrZb089QLkQKavCtFyGuc9TybSyAytJmF792fTXtRE5YnehU
FAJSLvDxCtR7mrUBoF9lHbbmyqqr1hbKBlWbq/NIMYrofP3j9WGOBiSRLEiw80jkyGSv5j8lcBAa
CK4y2sHgNfjJVxhXmjAuBAvfM8a7Vzxv9yxm4XlDtE3lWVphOEd29fNlFaGyTlm2bgCrei+CfqbE
uRjvYx+xP9QgSHmmEVU14nmi9zkxMXnTfbpnxicf9x7U7Be0P/98xMK7Mo3iXoptWWBTRE/l30Vq
jC5+39gDbMvSr+liy8SE58nzJcD2RV3+Oh/p3eQXiXtK4juCmlLYpNiew00tWR/o8K102Ur4XA4e
6qU0svgs9xMec4ynHKUGJg4JT7TmHbV2yt5rgFXqjwfQ3kHTCf57XRDFpJWSmZ1K+CMjs+YxJFae
waJ+9uTBBvs4oSmMwoUq1rFlOW2zcgI3DqwDuwykg3NfL4nHYMvXRMeGQzQQa13gOXTIjLJetfNJ
g0Oo63Kclh1mgejQwg7oyty0DCgKBvIsklIwd/Ubntvcep7F4fxHMFjR8kScfOBNwSQVf3JxWvWp
PG4tSffO9iPmxZVTzM1Q7VQEOjN+GPSeE97aHyfHuJvh5Z/1pZHS2B0JNUei5g8ascM6tuxowHxo
xpN4ORlKovGpYgg0PXzNjCJO82KFwumSkfIFIH4F5JfWnava24nBB4RNkne+1yXrNp3Jmk1wEKr5
Zklk4otCSO3RCK41yhiLf1eQnzi+tcJgozHrtffQtCS9TwktdI4EbxE1HhEYDduP3q1AoS3Y1qGo
CaH2ZDC6XJjuSg0NfTr2jF4KCL5KVeOQC//j0fEfRrgyvnBPe0OuxKM0k35koqtVqRYYTiAlRfcZ
etj0s1mocPWqDXynxKvVf6DzPmJhSKA1KUSwpQkJz5HRYK5O/kZOhTeWgV4133ZcZfVCoqPKJbpN
bSBcOUSAKtWinPQ7UqrPQNuze0FpU8EhJLM/PhhKNKENvgF0SRyRjpJaFwy6mIBlYYDWqSSDnlK2
Km/3hTUdcHyimv79smRv45XjlGCOJZLfMe8zttm7cAnGN3FSVTcDbkxpFmn1wHYV98shrZyLoMXS
FP4NKK0Ngd3mUPxoaNmjWVgUsoIx/1Y/RXUsiaKtT3c0I69SDPYHlhnuiBvirGbCHZWNpwPf1VhL
LQtv9p7jxupViYCdxWI74Pxv0jnPP+fwzR87AqK6AhGoE6Uqvpvyb8SkyQlfC1J7SZLMxvtLkBV4
73m4W3KUtxlTVyYrwmiI2JhnJd6MIWW4BU+63gUxYdP23ASfLqwFYUUijaatjdCtbhk7SA6HLSqu
8xYN1VjQhwyQOfAC5yhmkuaLM4+qadz73U7MlkDSuKk825wsQu82tblFtfP82BCRtRwsgg4sbCo1
avIlPYuJBDbd2oyx5Y1RztRkk3hB7JofdsrmMZzSMlBrPTsyuRW7aROgxaW6+fz5/7qQhpx6NrZu
/P+52j6V5FzVunvfvpZboZmw2OE2X12JpwMhImH0aFJUZUj43InkQZlzHSZKMoN7mRSAvZbWiiCg
0I4afts8wKvl71q0UKi0ip8PbVPrCNgFcBiUoNXUm70qx/du/Kas/aclsfj6almj1Jv+ty7BG6rE
Hv70peYe4OoWAyc/J9FF4YrFUps/ql2kKxKlJU/peHOmXe2IKDvcFYgSzHURNAZBgEU2kvzixa/c
41WfI6T5P+QWCMu2uBNjnGxbXdsn6qsi/GmLcSiZ2c2HZeyUNzFZaTfVwS7djhBB5YPRADchVf3U
xhGbQA1EZmf4tptPhn+ug3qkwBhmFBKztOH4LgKuZuWVsbcYvCHo77t5VaqNaNFcCzm+E3dW6ipu
j8/2hAxUhMMMeBKsctFI6TFbzpic1ZewLpq7dC/6r5lsGqsr8eVyA2Soco+BY37yoa5X+Bf7mqNp
lMpYbPGgDgVTYexCWTO6btl9ueUmmCe7yxeKjmLqz/vjzqtYHWQ2r7jr76Qzt63wW4Df4RoVrnqi
OD9hi46XVmfuiKUUOqim6u+nlkdZnGYbsL70erNq+K+9pOKZZWhrNTV+YghW7ZbTasLdFZ8GKpRH
J1RrF6Nj64+AVvL9FBhkqmyJOtSSMCFiOuz8D45uGvBYYztqR9f3piHfgfszfgjNxElzDZCfETbr
1ukupP3hXEqtonKuqEME/kBL7AL4Dj0K5AegT9ADMDkjRbP6y3bDZ37nxCGHR6h9JRVKx7IzH76e
JbOCjIOwVagNYg2i/3r12wH2wueb+6rjuP+c05HQxyhfnMywcIgIhgpWxpDIsLAfOuSXRTxE85td
7OQko0FmBsfkl0ip4isTofldmZNHIe6+Z/m4h1pTUQNt6WV5ECp7BPRIKrmhTbggks8r2Qv5cSzp
GdtQdrDYUflPuBkKMBjJ+CZxRy+E4Nx38MTYxHgTKU+fY6jVbWNdervbBjFYKE0XTQqy4hy3bzce
LLyVpX8ZA859+U9o6J0xcC7nxpNtVPFR/ze5cvAbrVsEh1s4dWBlGP0tmXNT2opsfoCj7yuSBxsu
Z4MJbJio+ywE5VO3b8zEHW3ROw3LuysR/HY1f7WlXtjvZU7imvDeW9L2J2NLGtCUvnWr+r3e4+MC
XYHdkwRh5V4wb+yqCfaeaQw0+1Evaas04Kp2bWu6YyG39NiqCEcIeSP26zF/hNwkL3lg7Fb8p27N
UTET05gmvd8NKJ7xGYxvReH70VwxzfmNcXPEgp+7vuos3k9+RhATv2hMjVh87Cvdqb3AKRKnRowi
4Z1caYl2Zxv2uzB+mAlzZnSK12e/jBG05GGJ1esGo8WSD9jXlLOCR2eKKK+fjuUHPtl5z/jfeiEI
ewV2OaPIzSjR9Ja9bZCSbXGSqhHWFbbWJEqVYtfsrQgP2n2iTF5DySm+mxFU5sJxlgJ3jkre+CvZ
7PlSuXoPGT87R6ZKaeoiLpknZhxOiLLSNgTfePlrN18Vd2uk0pUVVWGASVxuCliNN6fTMcTVtUfJ
zLpWbHlWI6D4AVhwkkszRGOet61kBFOtDO4lP47AHfr1/lbYvXSHJ8WRSkyPRRndzNBWGZjDbJfN
ADl2FJO+bWNRlf9EMKut3lGXK/4XqZAmtuj/MNZKs1L7y6ULsA2JHRtjplMtYmJDwwEPWLcNUv1O
JwVKUNXLZyBC/U4e91koF54B1FZbP8LCQz2r2eJE+NI5P1OsvXWzGkRPPRt6ExTjSynBNg49EQyh
Gr2Sk7sjv6aucla/EtGpbJtYaERmZkytXopCP1g4Km1lvm816MVHaf5YvwlPD7YY3Z2k33lwqpXI
gu6CjHm0W9xYELhECOR9yE8JBeX1vGbfopZBNi1AxB0HOnJ7jI0DbwVStHhGxJDWZ7m2m61byCgK
0L2d0Wn+ugi6u+UXBpq2cVF27YTPIsvA00lThacuRwAtOV38IdpiZmHM+OCtcOKHtr8vd7I6Ygjl
HbT8Lf3dLUSbcN0v3SWtDVF1/PuuLNhme2uRh92XvQfMPqQjuBvXLlQ46GEWJCkXmV/tzDws8yjy
Xkj+2MeY4PexC9PhORweDb2N/kMTG1Eh0WWmlem4I+vGih8mqTTYrbtcKPbwUpqT2BH9L7DzC2ju
J8QgCzlI6hPlWTd+ohlDC4f9RH9z+4vZI/EyIAXmukwXxd238/s8EAHOA4Jgh1DZvTI9+9o0pqvy
21HNezVXZJptdDACpTAE9wZL4oSByOLLYwUigowaIlStE95uUt4PYsgLaU1xaTYH8PriZO3xbSBB
296rDkC97+gCQTnly+K9UTF1/xFOvMmHx3GNuIKj/VVu7DZ6OJvOsv2dzeNdMgRE9guM6cg59bkv
5N5Eh6As85ceQrWIXPXYdhOXxMSVCEgXoDuYjmMCwaaic80fjPae0FEbcq46jMfV4EcddvZRzivc
hC9hHY2bMXmLORiOMAlWBk1xBquDFYm6phb559lzq3uCtfEKD9WPz3ySAkpaYMxGvEfVlfoMKali
Uw+pHDuktLtqby2O1OOrzq+FRv+kQqWgp2h6kNehXW7r5vTHG+0wVoBvFrF+VdtyHUPcXUB/wuQK
KSUUMbZBK/ksSxHL+y6CCkglYd5zncK9jPdx5mi8yR7Zat7I/tlIpEbg5F6hbMpYFh5uQoI4dgwF
E5yGPfo9sKjYlehLkDdl640Dzv/hw0VHZC1qZnMTHmf4rGNsXHzuS/GQNrMrprDomzml1HL0mFhB
iD/i3GiGt+U3PH+8gqiWDj5LdDRi9ZUF/Zh89W2ytotXZlWYrIZo5ACe4+h9LIk/esLhosH3dRfb
dqkNn5rEXGJWAFoCdkI7EuxxQhtIFcnKATLfk2CVaTQA5TV3eSq7+9nkxPYAEz/NeMi7+4wPlemn
0kOQPvd2RjooWT3pmmbFbj2SLDa/XLP0FlD62mY2c4VZxvGPiWoWAW8YKw6mx60WPrLeTwueiz29
bpPjSmAvdX4CQaFejXA+f5Zsq0LKrXjL5p/s/cQ8jsQssGyEPYHkvX7T1tDcaPdY/lNwvmBT0Y1K
bAHajIx5NRkQvVF/Ixpozid98j6/trgjjxJDTxOZ2948YuFzvDnzGXALrYz+icNnH4HVrgl/qM10
/jR1gNh+pZvVzSJQH1jVZcSSUmn7+nLzF/NHBfcK33ewMy/LL/GcjQ6CL1f2Mt8Yc43zNAMUrFm+
3T4FC/vWThSGaYK0ifnbARS5JCjcOgtOCYNStcWFgvgO6HRsiTuySBkRfcK492x5m3x+e9V95iRX
wP6opJSwPRIZr7WzcyQ9ahsKl+KpPCVXH+tPRD3Oy/OsBGNaLtoM04CIHWGgavlOUDlAk9lf99xe
1Og2usy2qKQAE98QI0T6ugPjnxKJldty/nujHJv7zLOXqHKo1MawFj0zLTIU/KVaYnrHMzeADjFH
TAaiHstANZYdar7tGxd6SYY5gaId7FL9AAC3UQ/dQBCVbW1trneMbG83gKBoZO+tIS9mkq5QtmRZ
XIql3lita5YCoy0giQh7/bsNfTQp8o1c1GS4oFL0Q5+W0pNZU8rd80Ke7tAmRg+7MyliNbWJERqt
OuLDVeo1vd+Tv1IYTvUwKWt7rkV0SAu1ThGLJ/y4T2AO8cF3sJErjbwceEakcYLIzKWKUXWb2kml
32/5s5jkPpH+riX+dg/Juub+Pg2ZzP/F2RzhvqNoKAqBWtrzzvM3+sZTJXlXdW7pYwiHx7boLDZJ
NgFM1VWfI/LNd1vuaVh1P1iSXaijuZnCr6xes5/wWg+/Ov7H8wT6NOr6W+XQ7hUsAlHAjiwzHqoX
TpJbuUIyQydGDrUGLHLbM0bXPAOviVA3xWG+sjOtfXEn/peE48V6E7RBPjKXdVHuX4p6m+CbzSAl
uRt2ozst24wv0uWFnT8Gp15OMJFDaNLJSqTN3KYj6+iJAMdSJOlAzjEtVXlMYRAgD8Uz/bz+7wRi
pITp6wJn7nabxUELCuBiRovLLkBoBmkYwyrwznJ7fnWNB5Lf+CV4isxlQWaGaV5VZKzL1Sh2YsOp
UsDpmNpW3msIgzh1bUc16VEERXtgagvcadlitxq90kkSBtSB0uKgHAXloC2aT73oiVqZJNrLpXS5
IDPnSG3a8KIhA4lrQPeseL2fRG8D3/Wy/2YxN9qh7TQSkJLRvcW6Yd2EzX8gSFXklvcrV3n1CrHS
deng87J3ceJZkerMGnGibiIoNyJQASxIsn6iPa/TM1vuX9uRy816ZCh3IUi7EPN3chh+F1Q72McZ
WkBTEkEKXRH8Z1GWBflMbESEb8y9MGp+rfgEkAlPd/g8YESBuGm8qzMAh73Bs9I98D7YP7l/XpUM
GKGGyhY4dZR3yv6Yab3xdSROHn/D4POlCjbNRUTVJqtQZUkh4aiPLA2Az7kxs5tAt6ZAesaLQg7q
oxyU3RczuwGHQ168oAcLAjMqLw+kpy1rPjfPl9xRC0mp6Z/mtiFh2LCEQHvN1BPMD1TmVSiZ+wH6
smHqO92rZ4iYRfgUzXf2bYcl3mTRxWAEnzHUQaji9CmGKp15RRpbv76UdWtjC4wZ2gNd3cg6XWf4
YfAn2Bz5GVfh7a0JlHqiFmMQLZqacDhsowRe6JLNdZi+3rFdwH+ICslgJ0HalOnbjFvAXLn3tbyb
62F82Q1BnnlHnj2qajXs33sBMErT4QPH32ofYc+lNxuOMG16MGzX14qfGt45RL5cuWV0Sq1Qc2FB
YXz7Z9bQ+D+60d45HyqjEbg/fBX5wMGNqhdWdcqmWAEmq5haMs5hiji/vmYGkWvGeCmfp7fr60/H
R18/uiqvxO8ejMDE6KMP1e1ve+L4A/OAhSQyhC/5ARTIwWU1mp3R3AvBdHrGp9MkuCxvC0x2vkYH
7n+y3X1YYLGVkb08nGa72CEy9YuIq3vLXKaoX/ONANu5eB02/WWmj9668YKg+/LRCDj+IRgXLFSo
WUerpy4tqkriuCilg3GArWyFwISyl30y7fTGSMlnB47SgCv6JrMUYZQQE6rN3XhYMbSYqqhcXPge
R9nPeKuXxNGhJdYm781PvxtsjUnZ9WJKUieW8oqs7NdcURjqZkfC/o6YUj4bx730lHqm71k+q+9v
ez3tLLPvxTICkZFsfp/ySPXqDxzENx75PAOsaY1sEhRxSegoamb/P0gAlDR44fxtDF13ViSV1CQy
WZTotLeaYZoQA1VBLQX9GQQgBS7yV+7VgtGXZu/UWcNMjzppueHOR8XfT2OIwUfdTUyAl31Ecx/X
221h9U84ZAqZj8b9RCwj46wIC2k5QSMTzHs6LfudFaPoSiLVfaTHY/Fs9EwZXOhq9vfBVzrj+vAl
53+1DvmCdXvNyM2DE5s59q+JbgvW9R4LcLseXQZT59IcIV/Pd3I0RjuOWEef1dO5aZaeSwUnXKtv
mncjMG3IyKQ8XkRylBaQMzTyl1DP8DYaAWRuiY4z3jwv+FTBuS1qX8rq74Hf2/py3c0dWh5xT+/x
sc56BWEtr6LEXnFhAF46l47gN/w2DWUU0nMw0fWRNUh4ZG6hzGaIm8coXTiHppQnWl2xTTXJzDut
Bi8tLNMuVPJh74R3O98E4uWKuGZh4/FOAx1MUmOqhl3ZkUneEK955ZoHkoDrKbQ+vxI80S9ocyxn
zlCW6lCarVF2en51XXGQ+5r4HDsmnpFSL9tK8bYjKgGLw5G/zIw4gwSrtDSaxwUd7uoqMox0xQ1U
KpuTZfTLW9TmkH3XqqGTfaNmKs/w3q/tjjm0mSAey5feT5pujzBZziKaCUj/LtBHxaB/0UYzXxhR
ojaQ2EGaWjo6UnDxdSmfRRHuxWbXCge/4SkKw6LDjpg1IDfRRrzVxHtnaXL1a3tUMWdd92hIUMHO
6fOiMoTc/6Exwzlvprs7ZMzgQ06Snl4h2G+sW15Ffp2XbfLiAQGTPjv8eScGGV9YhHrrDDsznCCE
xYLkWwt9TCYyz6c6FHB2eG6V05UujpuGC9vhHVT+gPsZI9alJqdu2Lpuhmhc7a3S/FAixFPvaRGQ
6bPKMfEeIb9Gyu/a4l6W3EZTwYqeTZuY4TytCr5DyVoTDjkaHhOPRp+WQvIO+4h0JYc0T8ymyFYm
P/tJ5sCaLnSL9ZI30+pCgcP/6ZszZ8Jklb0ORWo8PduxxeBElSv/i5YugzkL+l+VeDW2PAIgDam8
ZGzdWNoOp5BUUgMEljSoEp541FIN8SjHjEg4flBEkoGyy4KDf/x6KAfE8wNyFusaflUyDz8/I4W7
5QBxB3GixfNd39XrpXC70gJGt732u2CFmZ2bVEkoadmEW/X4Lc7WOSc9Q/Wg68yd9AtGzicH8JyM
QqF+OTdzqxEafbWKscVNm2zwU9Pqhb93RoEauYg8dsITmn5QeXUja43ufyhC2t4+Nfrta9320Enr
G8wr1UV+GprcdZDQw5nDWYxOc5nQ8F/EvIKbQwVg+aTI+6RkU1FQ0IXgsgg7+T8608YlGo0M4FUx
7VArBsDfEWpXR2nPf3hRbt6b/PctSPcAcDxAVOqvPkgRk3aWYWCqZtM2af2opCb3uFal3Pz8jLaC
3aXoE0drv2Y8oB5MSKY7IqpCrd3Jfk+dXc4K9zPkImKh4gkejkB3AjzLfyclzgnTTjyOvohRxONG
sxYvoDmNMWoElJjxy3KnGgc3E4ej4S0e5iYa6ELuSfWCnL5CS0AV1cWjs3Cdr/GVQfDDdHx7dwfv
EQZtTuCAg1xsomB8lKwQ6yMgzMp93y7tIAntyFWSQo5itnLp3/iSWynfffBGMH31GhoT4BecTcuX
L0PMKqC8UxE2zV/XKJ4Z331LukCbOauVHHZmIPxPTR2W306vsHxUQopT4k/OpefPdyUCD0OXS/eJ
ZF/t74YxeDkTxJHLHlMP/lTajFxcPFB47XVJm+JfCQeglJvyYK7CdyKyNkXZ5fNGqd3Q17KfYyxg
BS803YrsNyZ+9GoXNNr9Y4qXZwdhTtuq/02/sgugJngChwHeEiW8r3eHTJyl4T7Uu2YDmwuVeDqS
ew1CNAX3sqkPqorHHE+G9srWVLd73Yg+c5qG1/3aUP4dRNm5c5rfDFywYEInp9hsx3q077tkdtmF
q1tjS2NPGg4HzIEdtp1C/RXYTOluvk8LL7Pbp2iQQFKABD10iUofMxP4nYXv31FwGT3AMxAciIC4
KtGjwf/d675K3xQTln1SC8FZ9dX7m7z9gKMJyK3a7s7W2e4UieWFvnKDi2RIi9QMkF9yBRsDZ+5L
n09UY5+HTbY86fxzZEPbC0dg8Ve9+JRmqAYG8ueJ3RLbHcVuNVh67KMwrRKavo/koabVGRPbRKwT
LQaT7jyNzHqUPjRtK/7svvA6BrrM/9yLoDVhckq+4SbNNBHHhB1LNTrsxVB9YOFmyAtooJ83oQvC
sCeKENrIAWy2JPm9c6OMfwzglCIqVD+wkLulmajGCjGCCBDXoyz/a9PT8YOhtbnPIpao7UP8Yn6Z
RPOsGnkWaSxuAjtxojTF06BXtr6nx+BNCRuTJeT8IaoWq6lnPA8oa/qOazvyaZScSlpf4bFs+uqP
/u5jQods3OHrG8P8u9L401K/YE9J7rQiXQGKkMVnq99QuBonwiHAbu+xk9HrhqOeoTsFxkVA6bd5
zimtOoQTxBE6kvgXoy6cptOG4LItMRFZMCfesT7iAGkiSZArhA+CWCIkpunbWr5mNLo/LPkiWMgh
+X7nrC6BG3/01aEuUpQkkzw8vBz3b4sjmjNRZKo1UOeENuKq99XAYBFyA4WLm9dNrdbNykolNZFz
vjX8xJNyydC4864KF+EKOPADILu6h6IH2W/9HY3KWkEkRN52RZhnom3aTkpdNc9aXBcQNQtYUGGs
I6NlF15PFfCOww9BrUFndkI3Vrs8HkH2pihHXNBHxMaearSY5scahMd2OPmjj4ufKg0TcqyDuktU
wilGABHi90RVVJUXsQuaN6oM/WmcF2BBNOF1C2wSLPnQgGCl8+U82WLCnaVBNzXeDKQjkWTJKwGQ
OxDrhLc+kjDaNAmZJkRXSOPgyFl0KQbzcVAUmEEUCiy9dV8SMiqprUK0k0LxhelMDtDuIkvsChTK
rLKvwNAHCvYJ9LJLrIsWFNL2qOac4Yc2yBry4pvza0eZ2a9opGXAuolo6ygBvLU3wpue8/iwGWre
20sqSR/CB7SYRTG+kmsqeZATf7Oc88Cry3DhS33vNgnLy4+GRUNpgJY7L1gmmaRMI6b0UCXc7zJK
+x9V4UqUGRfdYqtM61rZeW9qwyF7igQwaDhO9DxjdYj6HPYlUm8q2YKRGcHai0mw8HlejEO9LmUQ
LdvXgQz+gPyxkIDRKga8ILDzWVedi+hiRvyoi6k8pt7Q8d4a6T0HM+h1hRUDRpb60iy3qZUyZInD
4pl+mlrd32T7NV4bZ5+9GNkuMryKdy0FiZZPt5HagJkq1tqni9vsZnvraCNdB2agFNznS5ne7BjJ
zXWDyd94+Vh02iAUkf9lOS0yLlgZfkKnNF5bOOhNBAQVl3RtQyOUCg1aPelowlJzRhZ+vLawe+5I
r6GZeMdCr25NWuMi6ocQCYQT44KM2vJqBCR9sJK5EljHVGb1YzGy+xWLlCESmfO8KZJSyZUmzMaV
cmrFvORgy5QtQrelnfOdurkYjJh3QpnpV/BPuHfhDKpC+zFE96BFeRHyIr0FdJC0PKWwaaselg/+
BACnoBQtmsI7n2vw0rCZmzAN1J9Q9+jGVtkaa3Wdd1XgQsA4AhM+g0NIBDJUhQoMCGys32whRZ5g
6cEnomPNSRRIcW/97JGnx0cXmsH5TIHfvB629RfHl4qJab+y3X3EWTlZPViXzVaixaPAAJ7NXxfh
nauV4Lc9pUPJoi51hGOIb5z+bDf4SHdZX9ys2o20S1IiyE4dt/rYgPB31an8b+xi8OlpKYnJa+tl
DDBtxFlLjXxc5sIGtckNw295/xVGi5NizYk70FXzp7kS+rrrk1yquixi54TXNS8Vop91/W03++4c
otpGnOEuG0FHDT0fmZi1lsF+frXg3K79xA3lvgoGLjbvZ7oa97KB9WZHodhmXHSy/PLNbib1a7iV
4CaJcpcqHhULILRE88fBIDTKalUiDhgdRivpn9JTghj+zEZ8QBurl/AwshxfjXf0J+05LYGvD0+h
kjVoo03h+48DhIJAC83qOhWrrRCjhpMcme98NBK7ynHXfLWYXcvFTtOWkrZvx2Z87xHhVLBrUBzb
gR/uVSIDwOoOLUHqWW099INJY3EEPH+76fGNzKgFJA/3C3IAIJKN14CrfKR5sCXIFZed+aul6+N6
g0YIs4Wvj//TS4uKq9PA985buh5++0r2rY5yhFqKNb2ZSg9LxDPoal3xTww0KF+eDmAnIZ8FMMgI
Zn9uXpQw2UZgqPbQ1Vn91GFl1q0R3VP8+2CPznWldynAbI+g/iqLU5IRjt95XT77ZG/GKh7v/mj4
OJj0rWbv7hEa0Zm0RKcfxphQ2tan9dgNVUkipvHiXe11WDSpoyHKmP9QhhEDDiO9Dv0NcUo4dkxz
Q96sQolNjwtOjr0T54UwOmSP9orf0V0AGET9VNaSiVlAlRTK6wBsxcCogsZrhAXZg8lL3D5f2tV6
XBKiqnIkiCwLyBfWAGvPjkOtObcyc7ZLYbp1g3pH/iCms9JAQv1qEV0pn7RJXwCkjb20Rrf5/PtO
iwxFR71+ZjaUM1zBL2Le4RPkGJGeMh6P+jBxJzUJamTp7WmW25D/AW8C26/trFiuVMj6f90EoBlL
PDBuZhTuDz2BBTLDj5e7XulKgbGO98/E6rzyimscdbCxI2M1hKrmSfx+gxqMUECpG8sHx1lG87yO
I+AVaGZ+Q61qtFHR/wl8qcyHbOTApLhQy1WhUnyz6bIdgrDF+ttvM0/04e5vhtVpYXCm6u066bzu
7GT+xS4vNwQUuGIOQGyJHEXPUaNK6u9hylBAG15iO4ElngwJ3dVMrsBu/20qLBR2isftxRYGSppO
st9Ger1GQDbypxL6aj23eQBayi0iy2lkMEOtnCnMlifekSw76zlkIhwti+KnjOUOMCxm4/wH/TFR
0YEqxuw+DA7MtZ/VxUKRGAnqz3gSsl8f3gxBqXXxEIY/dNtbo3C7m3YeqBL0fcFjkDugUEbC37g0
Ov5WIaupnlNDj3cLEyGqUpqPf23lWdizwUUnq3T2a0+Ze8OEkJVU5neLOyRP2oYW9DtPDxz7TF7s
zgClNgFuqEDHizcYMGCB2Es+9uJ60u8+YfeM6qK/J8BX+qzj5WqWrQjnBBY7ggK8kLT43bvZujPF
hAaM8XclceaPr2XHBCgpB42E71ycAQeYCokODARG0lu2m+NsBHSXofoD2MI7V7vafO1mT3+iFVZd
hGEYDAM4m2oCpkNit/PnryI/sNt3F4CrqZOix73VaDgxHSMksl1KbZT/AUfK/3DHslkio09HCFye
FgfYLUrvH74g/omeiqNfoRxDsyayK7LfYcMuxMDkxczMupbPhpnCaqOVVlnSDUjmnWHLBSMvuuY3
4D/WXmu83PViHybMPlqKtx0oP1lvL576e0o76/qbqUb+soSblxoGTAG2XOw/gHmQ+pzyLo4eaGfN
tlEysMixIrAY2mTqjC5GlcmjkFOJqaCC34tV/zHcFgQzkSy/T6VPqEpdvKwJlyuKercVV5Bw0LlR
a4116JBgVSxN3HLaMqm6Xty+ozqCthUJLgpyOqt1ENPiYKQ3NwzufC/D9a3vZZGcHq2HTCqMMk/8
malPuufzglC+GlZtqtolMmBp1W1fqJ8se+zmLdnjqzIHJL3bXoNYLJfWDr6tFUFDhEGz8m0RC/nk
znJPbFOM+TV/T9PplS9w/FUMn5XD6J9PmkFc1wrkwWWavYKj8s0U9FZiCdCLFP2jgTyqluHyNW07
hwwHnGmKpj9RUJl5vctW8i6AJV0iPmJGCy4mNsBITtf10NWbCDtpGYgA/OGhOGOn5cOc8luKLxX2
uBQLGncbsM4q//fIZZxhHd4oCwkbqCEdg+TlwO16YEC4AYamN/cUQXbkGfHjje/ckYnHcCeZTHOS
9pzBHrNtUro6iruHLwPbEkvrqu1qq0Eim1ba7QH0RuHGbLK7bBj7MzoSDXs2e1OrBizLDq5HAUkK
NxO1YLzfUB8CZ+npro7Irju5/Bc4K9PzM3cKA59KF+ooM7h6RI4RS1q1m+vCyE8MrReTsRE+AC2T
+/xZDivTAX3Wa5hqn1u8S5pp6UeoJWVyuCnpOEGgh9pyHzFpxyzZYv0nN2ukrPw0L50Qgty+03cl
K2WOyz1x+WZiTAwxXUjGQzKC8/OBljVe5K8ALV9mvBSwgGyH+Ak5UTIi0dDlnL+WPNxmERaFe6u/
NUH6+RALl1r8dgE7IMlYPowmJOGXIOA98XOaz7eGZQXABYVrI9L8Ubc0jIrc7Mh8jhgVAKKMutNf
Xm/9ZUL3oS2Q6rGfhEmOfkRWiuOZaHCiQJDqqnzKwcxQzNLNRsrYUTUNkm8S6KyFOWpN2pB9tjJF
8ii1vDUci4Pd6l1WB3ndithutBhRgj+BiEnpsYSYHxav1K/oeDHXY+qnf4oPvkXTrnVkq7L7FyQV
k2UHl1fmiOzOssOuNW8KG1LCjvXRFpAxt8++OmsCfHuL+g0MWokAym/5igcersQlBE6ps5GRq61e
o0XCuSRV9U9+oJG+zIlfzNY+mdqtxY/tWL3VqXj4mRHvwmjjTvK1PoxgmmahItPNYtjQMvVVYlez
y3lhe9U+SDQKpa66J/SZQNyTLb14RsW3ZpqGQ42BVkZ45Y6eIBZwaFOCaiLL3mmGzU6fI8qRDnc5
2C2nqy944LIDJYlz231JiH8simsCPmCMMsV5dS8dJ+Ew5kIoyPvUH8hEe2toNSs3I+m+4dH0KSSx
gtWaPZ8n7/MmNDzfI/WftJ+XAtxky+4XyA6Fc7anoHyIyR/z68ahSfit8br4vS/LvE+LsMRePsWG
Nq5NX3hAKchoFg8ZB+hTUpX/IX+JQO/VgmQ/TyU0YM4X3+kHzUEjA3xKArVYOUzo4W2KAI5NEKyd
dhMR85nUiFKHQvgebiN7Mp33dCLJY7NiVeFnecJzUOcRfo/U/0S5OhPO7XoLu07rsOfrYCSJibLi
oPC3sTE287xWu/3s0ahVwnTqz0yEuXx5lsUuHVF0Dg4lkutcZKoLWOsC0YsnBKRsqFqFwx0J0Fn7
bQCyBwMkIpmBwZS6c6/+w/RtsGoVwTOxgbg3IJ8GQAdzLI2eoZgziBXPJCrmEK5eZAYdfkKsMRqr
+RFfvJ9a3tZpGtDK+IVT68z2DKP5D0Bq3MPFVyWCdCfoAh46qkVkFl7Yi6S0oNcE3iHi79rS46Lw
kUiT1JgrnK87tShoLzADu4izDEyAAsz5gqAIId6kE+MVxnpUb+uSIwPLNkarLZGff4Jxp82jJYtO
0OUtU3dlpWuo9Rm40USS8hSRe/vm1zJqowQu+0zQZqLHBnx4cJfdiwtwCUm9A5qNK+FmyRpJmEYY
w+CDoxFfZjQ83ov4hS9yiDjtzAYmwkoqzGobzOu6K2oi0zNJ+QwSQ/BOHvNYVQ3bDVYk9ZW1K6QP
Povr5kkAVNh+q24Sf80/pFhnhTdMFFPaIsCBT3uWxz4YXK04I4JZspVdRHQxB0IuRneBG5FpHX0O
TjBF8LcKCOpMGq8//eYP2V8Tg6qtOliJGCwCLVw8LRhzydAObVKuv05EPLkADCCzgofsvd2jI+se
2bESBkpDm/csX8KrihN7iLKUW+OGqCUAq/G89KnlKynjLzURfeuZ43Cti+9QJuD/bdxXYtDN2lPC
SGtEIKRrGPIuqbaU7mJa5wIkBVL2SX7EVQ57NBeOULLBtFE4PUgws3+45HiQD3MrFkFyEtnGqRPn
cNovn82xIrcuSyYwXWfnVOXm0maBpedFrU6aO4s+8ByzBk6yUQPBFA9G0Gb3ZGDcVSYQamPkxooS
7kKAc0sRnXyP+W54y5KvS7IHtt9xqom5DtMqD+BZmCCBe2XhV60UBhcSxHw4aeQT2Pc4YeSfLxHt
n7J71WRic8W/B6uy3kUR+U4Z65iio6dciChonE9fvbQfb0D6wzL+pHFZ7LDi11Ba2iNwqgW8/zif
BmX0p24s3xm0jXpYpao5L3XultQPlr0wLWK3qWM/ClMjTuFx3jeQOtkIYtpGQkJhLWGEN5lXhkQq
Zd7G/R68WxISma9vRbcxTY9GjgeY8brMyplIFZ4t2VYD7NCg/ChACPM7kMXvofGU5w4GX+tmBPQc
2jYpWuUB6smen6oJwHfscCB9mt09Hj515UBYfBg9O1ZGQnd6b4f/lEbfYF84PYa9M1z419a2IuOR
gp0cUhxjYDmXSrcGmTY3CSr8tJMWAU8S7YHPy8gBf+uBTIbpJozJbJmoAPjWDoM3dtt5wA7TSMh0
+FlQfQPZtsdMjHj16sZrravoWOBfbVswmeVNr/kfmv/0Vd4fcG259UbF+5ikBX6XVdJf9ZS9SHhz
MBvGV8XMKOpgWBUBgBr8Je0SDvmvgQNTrBtExkkBgHhg2y2iJYE0pgtUCH2Iz1a5itSuQr8scMaW
jjaSxAm04+V/GrFYFrOvIy0skl6EaGi8mjg9ZATu6rMZ0wpkzzq9FY79u+8m8ndpMoJAkwMJVdiR
9BL2geGI32zMZGeaEDVFy+b0S1utw6W7lq2WuOJhrcJ2zTQVb9CZOi4g2EJccOTDSnHAm+cO1d0b
FPBFuGGxO9NNAvcdG/YnEcuLzxw9pO4guvFTM/GG4iOtRbKZOflCvs/C3h8mLwhJlQxxNabLXxP5
XnN4v9R8uDkWw8EsVCyI3mtdJGMHes/cmZQ0Upl1N7BYPTIhHlV97sYQK9/3XWpMU4l/3qrz+RqQ
bWcXz+eKzVjbVvShOMpLrCBMobPLbKjznG1VxpphGLITKaVTRp5gNfuJryrtHHZtlvRantFWxN+X
hVUYYVClhC7o8Mbwi8NdvaqgUJtkAjkHIVI+cQrJ1WWwujPuZMWA8vIfnYORA+e7TnL9yx8v1suP
rml2hYnlCNAXW4FAMQXUullYUfyM5QxrIbGvoLuALW9NqgDD86+qGg22jxeamg2MZTAeb3ByQkR8
9ddUNfuDwmfGdFmFCkJEkyw/No7KLvDJRp9TBX4eQOnIhue7QXGrx9Be8SvANqIRTLfX5dJhqMtj
sufGbBf2i98cDUODq4UUKYUdOAXzBqTG0yKrn6BADLhIDlMeniWgOYt3uXKWlseOkOIA2shspQbF
tg0YK7xqTGfyhZ5thl4VjDa7e/OKb38iFd4orpBN/aXGPhnAUnaJYqz6LsgIEZ+wDR/PDcHmxIlm
XgOyf62jQSlxRhYu8wFq2OSJRcqnBE6M1pl2COhAw0xsWlgSjH/5Hy5wglRsHGzk+eqVcyEZEzvC
5pITb7AejPz1kwzdW/JVGSL4C5lTHUKrGX8D7mGXo8nOr45eIfsgAwgHvpeC3zdIak1doGKTGfJo
xNxWuhSvM1Hn5RL9dfsraF1kWN4AcxRHkfwl0i86q/TcNnPQyX3O+KxmbpS5KmepXue2aDv6har8
SiUO75u5FPyHU2mcW1VeBTv9iPYEX0CuqZaLEfBUA5+TzOQVh1fsqgjupd0pzMxbVlIvVppwwLYN
DN8QYO6nx9o67wThlWqWnTs/zu9I2e9uNZ2XmGNQ52j3mbNs8OMz+FuzJ0j6xbtuxnqLXiZK4yMh
S0v4nTpB5TDj0kIikrA8bxGaKkxrVQKghyyc89as8APJ/8s/let5h1cqyev1ddhtlm5cPri/EWKM
QyYrhWeEaNqqf0g+X8P1JvgIdvQQOQYWVQ67wsPZaPVA+PViiDRVi5Ba1RO6oEEXwoEGoMw4iRUe
75OQ412//vdAEK/E2st1JIxynqn1o8njWcn6fzMJHW4xA+MyrcxOOHrQBEJjAyw/buWqm4gGGm/O
+R/znkI8clZAqrj3NJ5uBlyqwGOY1t53aCgwdEecQlhq1Vaxix/xfrl6kbvE9eohbwdx1vHVjxQk
DPD//vtkckpqfiHSqyoLyNzaLN6t5oAbYuG1loSf2fMICuhWpxr3uotWVNAwJ6POTLWfZcxR5Gzm
Wcx2CqFPEHQZUmxjPpSVQm9a78ZhcTP+O5k/tiqPD81i+WmrMNYi6eEMtgEhVjhfP1B+fastwMU8
ewcIScMA4sO8KYuzlogf0Sfo1iiX+Fi9YnDqbuMrPjPExhX30ZnwxX3iamze4vc/VGyvqsZelJIe
Dgl3ILhHN/oew0Y4dELzf/evRxd+ET3pCaD3ioiHXaggpEU4OMb8IsGQqYwyUHwuvy87NyPkR30k
+4Mrcrrmr+tIF3F8n3tNcPxmguTYzfLTJ15J7K+5Uop2Lzzw4tu9IpaAmNiRYw2Va/Un0FhbvMxU
g9ORn0GgoNTYfdIC/Mf6DHoDen9BQduDExzbAZtQG4LtqCRPdy9B6tSZmXTsGEk7xHTRz7YR3GDH
u2czsKdE/yAL4fLQpRTlgBY+X1np7HrimInrjFih0CQaVwEkTuS52viEX4vt6MmAKyKGq0yDx8c7
eJzz3soUuAQqDDe5egx1QrckHwZTx5ywYH7nl5d7gQAEqgrxqCXQBKz+dV5FiTgp/fqRLRfSAd6s
uyCY3kN+LmXFR28Pb+QvIQCOtew896+Dw3s5nt71P7Okxu2DPVgcRI6JYUxKZhD1dtbiawqXDXF1
xcZP/jv9OSvV8ofHvQNEyCcs1Lnomz+gyQ3uT2fNa6pKljZt8qFB+RmSQEg/sV478+fgadRoBff9
0ajuY46tK1B4LlY2xAQZt15FGjFRhdVUvc8M911hINIwmavb8zWOLCBfD6k9aqQQYuN0WasWj3AU
LTlQRlK8RpDvjEGL2AHxHlN9LkgL2nOxpTyoFzpUkUb4+loGKUjwo+I4kPj/rYWAJ60fcOlUey0k
u0eRRX0SZgQGx2NFy9xPwgj08cfZCBwKRHQ05oZT3iqDzZnv6JxbrMpyDLasEunjCM4MdfFxlydD
N58VJYdyZuu5gppXEswUMPXHjNvwebk1AFTfxT/mcsM1Hv40CIYsV3VVwUTxEUEngeVhWAIYoBvt
tS4BNzKXZU7KwMJ7Ge033xMSwDyw/9gTFd+7J8jDXreGZRiaFc95ytEde4DazYwpDKkPcBLR0g7S
1OiJ0v6jqnPiWoT1zVhR1FtsrajRTQdQygGZ9iNHe5o3wENEufmfNe7/i/Au1GCoWbNs4TP0bsra
gSlSMp70gpyj4wOz0U9VXdzfLCm7uPpKshTIM+QJB8UfLXeJMUJ1arUNbSR9SKu0kE273jXGOxwu
xYJp1P7lq4uMAk6px9r2ygUUSrkg6hD1Fpvj7ChVCG5TbdEeHOGxl9+f76TgPa5ppIH7NwLvkPIa
54LCpNg9cfS8KkZwdhl+B7yxxntYbKrGkvrmUnJcKUzKsRawV3T7LZpW0QaBRbkwElO4IoBLz3FZ
7GNeKHfD1XwgKfqdC9zrr42ykoIx+qTo3TiKsqoGRRvfM6Q1g8WE8K5Tso+fEsV+tmnLrwIGJQjY
gXnjfsjLGEVqUQfBYs8X0x4t1Fj5K1xDIgkZxU+otxk+6JZ6IgNVtsYkJ23z6qYTirr7DlG+KZmD
nfsH8Oest4Lojd7TZDzRA+Pyw404VzEDG5F4VzXh934GDPxQ6cQ49nDbc8s/yLV/dOqLBl4+bwUq
R/92it1w77I0pG8UNe5mFasEmFQZFO7rHChHnOek3tTfvFKSVbtactucSE9NOw59SiWjr28sDbog
mmBZ7/XOv2KRp3LtIS4tUBtDH+p2Fpfw4civGLhCDncZ/7cEjpGYm0dYyBCbBYkNoW+vmE3dMszS
wf00hRxQKzHNro7I8EA3qpM01lIpGIs7Iu8lLU6tmKDkITR1IZOdegLyQRDFQm3eiADhjN+nM1J/
OBmmb8/rUCxHlk1qufJLxgJzc20xwE49Ty355x4P6vJPo8eToWhGqJaL5mmiZkA3O6R2HQ1L6orp
D7cdPyyLKWk9TuX0FZ+n9yCvtT0PLeEsKKmqagc5EV73TzVoSUV3tcaIGlxpt8J/d/ifETQLS5DG
fJ9iQ5Og4sgEKry1WGYlH1KG+QOD5KQEwFZNWT9+TDYWviUGr684lpQ6qC9vKyK/lA3rWw/P+ieO
21DnlxIfhbIACEGG4MkGMtUEkPOEyqUYisScURgPG37BySufZAgCIojZlAbM/m9/asLbWD6xjWDl
VuDo2RYWWx2In1NJ/a2X634gwxL4DUVUh5XeKbtv2djhzkjWypI/dHjmeoETJ3WIUtUWggY2B+eW
KWCiGjpnIPgnVsCM6MTQsf1uwwuV/NNvX51tXbekcLCUr1wYeUtRumUgHOFOSvzO4RmjaZxZOACR
RcnSjBrJFex8Y/9SeGgKmehbUKqbIx487aUMGaksJt3w0OjSaPZGouV3PBQpc1gRq2ql1leif7ll
e3lr1bB3d7WA7GMhgVuJVjRlWZgLjYpPIQhurGN1VnUHrBKoJKZWeRd6mJMmSK61ng6l4CiKwpk7
AKk6BqhNGxM5DtJRo9DaAfsj44v4uG/Tk9uUl5T3o419kh20Tdb5wKST2h54yrHM9wV6bGgxJ+l3
jmZslCLhBssYAoSxK1lXkibA4kvri1CWZUvnnc3VnK7VJpRDaMC+kBFVYkqXLFVjscdlehHEfzPF
Gzg3Z7UvOCT6TaRYW5HsNX6fnUQCJLeiO+MHyo9trZxJjdB+24BuN08/taTN/RWKlj53y1hNGiq9
7KdqHUc2xAp4WDHqnMFc72h1Nq8RLDhZjclnJvSw6wUAv/xn3jkrv4GY0Mz4r8CxC9qEe336d5HE
KirIIKAxu7DB2xZRnI0PnmK50pAgXpU6we6ak+3lqgfxuJgmwB1aLwNc6hMEk5p4paBgkMdccWAA
mc63RxqwlVp2H4LZqJjXZ3+pilpERODHoQ8E6C5MUmSft8PJ/dM+kN1K1laIqFgXIxg74U/T/eph
jTGpuPSJdsKZU9a8dOiWa5kP8wy5zKD1M45ErNXSVzygXKgvn8Oka7ttLO62LuLmRGh3os9iXxG+
FmiXV20fxcgHQ4EVcztiWUTWFk9J1mQsQrGnSaydSvl+FPtpFhdi2jtnwP1aweHSJIR/WRrE0V1D
+B9/kR07HrvZ0TL9gONoF0T6aosusLzG4t4uphj4UOgPYy70x0LPhNsqbzDnlnR8cjaPoS2kG6AJ
xLbzHo4s7kkBr+GhRi08yft2fQJ3QrXIvM7uZMzICMBtJjRK+aIT8HDhaScJGMruoxHDsKAesZNm
/Uvdl3f+OCehg7TMutCySJhr28ddMU3Hh+Fm6iTpNdDILX8wCY/uKgRLhyvqXY+COSYv13WH3deZ
loqpBabqhQUgTpzEmq9dsN9h+typ9B9auc+tdAdVzVu5A1hJize7X6K+kg9EWEydQ29tdZE9uUJG
Q8YAX/twZDVFpF7R1hqO6stIIQzFsl2WISjqmvhqMwuGhwgSrwgtEaf+uWF5bwWAmaCOlLPXrJ0s
jL04TJCnTNN5vXtR/dukTw6EeXCn6TZGryAghWGaPMAfOmd8f0GatO6fwAgAvJVzQuIalHGbmhkz
BJ6x2XvIdFMgxHgH5T7nvLcEIjkgfVk54603x/Wn+THsUEKuWl7lh2zZBeknL4n30XHncdXug94L
nrE5bIxRPjgE10ayhNV+ufW5aQgYSnI3cGaFaDM9pDsZ/fQMGmAoDwj4uzWwUJik+Tdm02jqJiqa
7fDXsPzYQb5mnyJGbrqWsiTv0q1vwlPXfnZPpNqevGM1Aj9NFM2HVg0VgF3bhzsBUFI9FF2kJXWw
fEhDLFK7JY1qeB8th/07dSpXplrPDDkHxq8RAcDFhFrfYlLiJbZXLzAjOOo89LLv8XmBugL1avbw
TuAriqJ7OKvzExYYY7Kck/yOKgZWYnMaeKBedlbOJlQf66BQSPcDuj5W6C9OSYnkN4xa9DuTTzW3
ii6xUMEZmbLX1y6liD6SwQBkJwD1q0pRkn0+BUejQqkEWbjr4nfmR6Doptupw+upCAk9tFHvENZO
CcEGXvd8KGYRlA34ByTALaiaK38xN1LNEkLGcX6DitYlXoso/OlsWz3Qm+91eDXdVvecN9rhBieI
Qjxi7Q0a+TRkoKIxu3akUdZeLZDHWP1/viug3LuFqiEAl9/7aAVm769MOBsyDNfCjGBudiiwLB9/
ovTm66Ua38jHPHaBgh/sT+p/6LIjFQwfJhqs4/uzf1cxTuOnb0RVzfdPTivLgRW2+1vMPvpSe61q
U+VJQ3Z5Zz8jVSWr06P74kzhGf81YqhSFyuXor/Ut4c5qfAFVjH+uS/NEIPUxxRJ05QIfJFfBO7X
XvAE4X1jnUZV2r3DQqOU8hiGz9wOpMDmqsc2HhsQwKlIF5mS63MKZgKeGkJuAUZY2wTCEiPO8YjW
0ZRcjAF5CrhM9ncK37/FZerpzUrl3Kc+D7osHk81vll2D4EpfmhCU4vCTx8MFjRwL8g4Y5YiyqQT
ydOablYxPFRHFM6dD3b7PJR88dHmmeb9e1m0xgFB5aIboDnS+Pc9HB1QDLCFpMwErxp3YAJIy8oe
T/VPWuI6dFQ+9uW7AnzqmptHRLt60FMnTua+vq61s453dC11uYo/tqwftw5804ZA4mmozcI1kKin
tsfd29Tolv6mO+h5RRSjpBLuACWYVIzxgv9OBALsuuqD+Y1G7PKsRddIQ4X6xFmu4VJDqkU5x61u
wJs5buqSkDx7nEvzOeR2K+m7xrr3pIsL+4kZLkGDwc+HHDS8mcAIoUZDCOcDFreV0penxzI2/lEn
pOMwve51Rs3THrlPQmIcQRkIgwxUaNF4FxAIeMPpPZOcpYs7BwRC1rLuA0HfeqayEbWW8v5eiWCy
KqndAfxxVfaCcgfPJcAMnFtSVML1zJUb7ZyBy2cxZzx2GNmCpvkqK8GBgUbvGtZ+wLqexGSIO/FF
+0ehNnkDeRKkWtGu+7TYbWmJGTXiQ44e9xB49UIg01tKDpcdwxkuzp7pwA3j0wOpUjf5SzMXl2f4
6I8B91RAwPpGzR7FOaZUAyBeDVHTtJvOnbopWfZmi8nbRCNabiy07T8lq/RXke0anhrccqwq8XY8
slvK2wCX5KqOx9tOykPMa2GlfxUyN3+zIZTEXJy2wCrjubBR3GIJlhgncW9vZhNpNaI7XQTH+mqx
I37PBe2uV8I1sF7WTGhC7WxxLm7FlwGDmB0gRhOzHKgycCl+hWIi3oAkB/Yapzyc4UviGHxhKE+F
uALgDHTfR0ax/nOMiJhf2T/SBTrRa05P5SwxZHlkgmKlY34R6/T/e6Nfrtli5leFRtHtwaXGzfi5
WQvNWVnP4tHlapsHlRPzJHsPm8Y6B6g6AWGafT5Naz542D4qEEqYrqS6Rtu3Fx2FJ/vNnQNdgC8F
IcU1DzrAHq9dbqQ7iciu3Hjo6k4pAUphebcVI6v1hwCHUloPBXFItwuViY3KNqoKnjxgaV69Z17l
ZATHs6FQ/nZd1OYXOltWoOoRWiHrAbGNeNmwvc8WcK8i1plPAFz5Ccye+DMMHCgPCZBXbUjF3tkk
i1zFR+Y/xBAKlFemAhQ6dWRkobCED5s8XORp77qH+G78Df+k+ZxU0HH47169jG8JvLuANDBMtIx2
zO7q5SymrcetV5bMgVvvIz0lW+L4VCQf+KWwpKaG19zikRGYFM19DDi+SQh77I8IJFuSU5h3P49R
ap7ZGflD74yhyBeWPfTUxNs0we/P0WNxD6kqX8lziAXHj4jhOmTfZtTiC+xQUbCJvUNmF7GhuAY/
kBzUO67Eoiqnfr3WPoYNPEwge8xMf84H+xmncQfCopMP7lNesjuORthXuDQGjz/PhQxBCqwHEDRi
z4WvRnaARNtPPVFqffUzM6OIL0JsmNdSy2iyu7v5HhA31+2dBRVPzedu3j6LUTIZuDf3DQ3Y37xT
cajv33m+ySRVvOx3Dax/hig9VbybHq0SPCVfuYeujLAhCQaLzvnvKlgZK9G6k5RjSD4k1t8lXOXr
Q6VvQ7pu30gYVnX37wHhYkwo7mWtXFaUyD/9blIFY3mCbrCec64AETk4NeY4IbJ2d4rjtWdc7heC
4AaGymML6Ke5YCQpk3n2zupF6UPQF3FVJz3n15ae57SUDbFuK8hZad8rchyzEMMlNWmUD2tdBzrd
9JiXK88w8tbUrggNRq4TtJjXWT8yzuYpK/0KlDmB9le1o5N7ZnCerrtzBYfsAVH4arkrCZW0ebQn
HnGZO30NpZqXqcMUJgrXGyRWpkqvGCkGD6DFlgmntvSSjiEkEpABj7abJZUW2quputXwPyxakOgx
XB9oTNKMYWgkikX+wxJbypT6itbLhY5W61o5dfsTMPfvQ50gHaWd+gAgz1XEjSF08x6rhLGLVW/V
5RKPYLQtQxBCzlMaYyA1NfyN2Evm8Ds5yrl3YEMlgR4BuZJ/eCFzCua/3+GmaTSffUISIprFln2o
fa8MHiI7JNW8trzWyco9d1UN3q1qUPn1fyzWoevuvLUyXvo5dHeN4HeB9dyfvxUxSqkl2sOTD9i3
kxHd3K4fRnvxGoqmhd4/rq59RBOg14OdP9HALai2CY2VUVrDxdCHAmNgFnFIHigmoOrelRB0wO/y
MKjctOjWyshaTXnebAqLmKVCSdjNa/cCiCCRrybqJ6gwyD9xpK+N1EmQb5qxLdo0Lr3sQA+SpMka
dVFToYSHkyyAuWvs7QMB3aRUK4qTzcGR+COfULKt2sst7w8exu91vzJ9BceZPxU0630+x0GiEUN/
w2LUg2TktwH8/uHAxGmgEUEuJHd5qLpmenwJgIea1Ap+pg2ubbFcsjdoqTrkKjnA3K3UWzgGP0Ys
XmIrF7EmEJrjcarq11dRGtXI0kAkbUiX0nkUBn6LbM3RmBEPwKwNFXd0wvDt3RkVTbzH7lABzcrO
6McMoo/XWgPh9jqycANBjd2iTnJuFd913h23C4MX7EOzoyECAVIY6qzx+jIXCxH81hOmpDUCljdv
YoFu4HoN3lI4DoYVIFBkYlhqIPJU0eJCmaRZOKY6CYp4K7XhSfPvoxQQZO8ucHq8zqZYM22Ph3xm
EPEV4qcAHRGbRVhmxGPebp4HJlZlemh4mor5wIO1NNgFz5RVLRhfYHS6P+WN65mL+pt8T/Ib3prA
Xa2iyI7kSsLKe8Ez+eQKVm9blke/L92Z0fa5HhxwXZWcz1QE4c/O//GSWY0f3aC689v45iE3ZQcQ
i5cctqJtvESW1yr8qCGMpLuhSjyyOkE5aPH3kGB5FqDul7PQobwjiV/3w2GnV5VnQRHLdLqE0SEX
PBdugCKoUzIPWtR3dkyg+W0z22M/V80KpepYoLVhInG3YAPu9prL4ZGxa1bHTXOyujKI9Kph/hZE
TQadAuXA8HEelYleX3l4sgPoJefJXM1M1pRa3iDYPwrNimnrMjUL+YX36ljiYwt33+stepe5h5br
Rhtp/v5REc9vioj4hvXMITkFwefDzvfcbl95hb3C+AyVSqKw/x5zt3Z0QV2B7gxnar+Jgbyl69yv
7gzgvOPpb4F2JrZJaepdW3lszk7Ky/iqCi7/YO+S118glQTbIWHy+8afL8Nq+GXu4EgCrWhl1dVf
0LMz+zx/YKRREn7cwzDCei/WAr5denuMkVZKnOLXFrm673VzWmx488A6s/eu5CL4VBvy+gEC5dRf
3/pYhvWyyxA8QuqapFcuIlwWh+ozHGbnlctRmHGuFGPQMlfQuX8iA3iVE9DKHF5EQ7qygjV8w0Yw
VhA7J0asHsUdeV57UJmD4Yar/JGHy43l/I2CHqfNfBTjkOcag4G97NoX5S7oa9vetYEPXeF4fpCa
BjIt7KmaywgCEfKUhwoshHmBbxnhiMdtdzuMv2Lol+ib8ZFznSHhbjVEH7OaK6d0a55yxXIjl3Ak
3i4HFmwBHZMuQCiIFwt3v8STFexxzt5MOi1/m77bsft9UV2Ym+T6P2LVL3gTbvQkKSkx0bZxkACK
uzJWoN2/sCw9UJ0ulzaYGnviZF/YR43riynVuQKELv/0fg+05RWzZE6+4sqhR1SW9gkpZazUSeqt
CLos+Z85nXMGVhDEnvRrteUv8A4kMC1Afes2l91iwxTk8+DKdsoKaEFnIbVN88xkFsK7oMGG/n6W
6t1FEmXC5WGR9Y5xPVU9Rbv3k1YZfANzkKe7/fqzYMY8xVcyyLOv2HUb5nx4TxMzqnLbgrujHUWg
F9IdSeyW4lTi7mlsRTGhHEyItrams3WKAd7wFI1h40ZLj2T0XK4wYzJH0oqCqQSbo8aV4ZxroTVH
ngaNFhAEihDQemH+1/iW+usPuJigKtm0BxdWxC6Q9SVTu0sS4JZimIKaGGEWjDnKpLKew34hXvJP
F04NjQ2u9Q95jEFhkSpaNk5f02jZusoBq8ztdTuVAd/YH6L96raKu+otXKDRpVS2ggQZf+Gnsubh
5CM3NFEQ8GQYJuQQ09p593sSgssqs+r9bHaM5e6WC3dtOM6jPdEaHZNV4I/LRyfVuutseFRFkS12
KhVdpIlSc3sElfpEcv/7LOd59KalgaHZWDBSIBEtx448JMhzpBb/K86xvPmgJrFTaVHg/e3GC0Oh
3BL9jd2KdDzjz62O6eoovnEMiV+qqz6d/qMP3IG/VK5s5Y3F2X2px0GzLkbA66nU91lgcmbdPQh/
MZcNEJF2EyfG2zBX2LA8DkyoLSZnu7GvNXcHX3t+8KPa0Wm2L40fC5xZef+2l+eLz1wjU9BxC3EK
lTxvrje6/92vbL9PBWXvsfrnTZgNKSwYdNij5MW/RRC84bl7CRL48GM9wUIIKg0yZTqjofXdGeIA
RTTgpYDdgrADqx9aoVcMC2dkoc8K0Yoij5m1p16cYM4zabGB8h17Rnh88sBGRE8hoiJaguzP4UXH
iOLP8YXWpSGJzIoiwdBoZgO9fnizIHj/3TqTvcupGbplIzTIxj81QssJrKW6jy0Zkx1rsaJu/BrU
ovqdQ0OJso1prj7PfbFEkjjDwWf0yf/bpR0W+QzkS2uXHfC9LHAzjxTbm8K1fsEPKmUD4E3ld5yM
wpH6nWkzTFRSbo/5+F4SGg3rN1zGFdJQS/Zxska1d+yNU79eNzJ90QiF8MFTH4N2+bN5aMSLjgkE
5BWmNxnPwttqfmEeuz5MdWS6heHnYkuu2+JFGVnMyzY9crvhWg1i1gZTrSoFwrl37mJdIB/LZP8X
R58ZtyHdnIh4gVeW0qgRDT+NpsY+N4n52ZYSGfcJ/kUH5sDOmjT6gUZE0d3u69b9Se1VTwNH9kBm
H8BCp6Xp6xDUl7gJtEPAay5OC8LlkX/vQ5jWzfOhEZwcZ1N3/RELeA/WwBLOzcvsuv9QXq1ts/y0
93b5DGZ5FY95hmB41qWFFT3W5CpIcKga4s3Ti8iZAXf+ymt9u+31jSGOt5xkFfWa3p3OjERygcgt
QIwuv6WuKe3bDoLOTb5g46Fw1j1m9b6lOo8TYg1MNiRHw6uOuYaKRLJxd/MRWjHhZIaUbEEBzAce
QZ5MCxLdYfx+mgfI0lAQ7tqTVhaQB7wDAMfsjg355ysyk0c/6NwHGqgBmBHTKHBGy00qVj7RJR52
holonkSaMZN7qdLV+TtYbmwTripeZX18LtxZ/G7Bg4sFVjQvlGnaLwvStWrNeqDPjUVyj/IYOf+z
JNbRAdUpYDAd5+MX5J6LyHUos5hKf8zR+e9bXkEIbh09OBpF5/YOhpyYOxBFUhLoE7WiU2qvFHAO
g+U7wWv5RLwwxjMvTwkbroDdcnaDGSBcaUJgBKAsqH/XefeRtYSDd+AOlz807IDI/OOtHeXx7O3A
eg7vux9G7Pf1Ce9usEX3ON5CPX00EkwI3McYv3oXkylmli1Y0Dp/ovCOMdKKAeC0m6muVmyRqWCA
SkHgnXslHEpgFgTBuXd92h9E9ItUGBRYrG4fqS4Q463TpAlltqTxWIG33/FswDwzFM0LYZCbWIP4
W2Jb76uoY5tWfSDg15u9cMVbkDid24iicYO4TwUUAX2DwHzk2il/ssqSP4QKMnmmVqw3bGVo1MS9
bRQCaDmc+VBltYg4KyQMHlRTY6RjeKTOjVPGsuDVE4QYEcrcvn++PjnFst8LE28RMdS11x+UFeYh
kiirAsxsHYmoBlctBfCggvhwDX+X9sJOVfzKf0uhutjzw5VyTpjdpVoxgQJ283TROkYhHDQhR5LW
A906OlXnIEXB6p44ke04bTDjlFlRPyqqNn9aE7PH508IJcaVzvtuhcBL/Vde+Hr2KjRQSkTNilRD
g5S+6AnEV0oSJ0SFzhGXAnX9knYp0jlpLH0Rs3Ghkl2h7N0Q4TX56SoXklKD7gdQ41mbjHprLU+Y
qT77mXTXrA2YSsVNcPpRFr9/KOaACz5iTo+I7KJZxELcIlYJ3EwuSC6fZGnCTL0O/GxQTva6wVvv
Hbw4E3Iy4C8qG6D+IwK3p4GHc0ZEzVwKPhxtVSDv8Mc/NDqGnx2aVeRS91N1axhV6pnVFNqjv3O2
fTQYeaGFyeT6czm+Y2LsQaarCOSYZaiO+b1OOo3CFcqgt5EgkcaSxfeSiIPsb1C3AyjtshKLnd81
7qakh2W8omcMwL2BBJTdvZAilyayH8uQ3GIXKLT5I1VO0CJRrXgl66eP8WP/OoqZQ/JvRPfw1eBH
kBwceUyo2A+EXDIL5YgZ26iW4xir58Ib3ZIkkn4LtXhHtjnNd6uqTpv8dxiTa40AlTn+gXEHs+In
ij0lpOo/Z0bYNGRBTqBaX85oPqvz9Cp7MN70XMDPS7jODzz421kn+e4JD+/ckzkllY5ag47Li5Yr
wuWyhG6eTiHXiOK/zngXIgj8X28hYcz9qApoE4fbERqYO0Fy0v6XKfBqRyfJij2bttMzZ2i7M0yZ
uPWEidxC8+voHZqHh2oxAqR7q6JUeMpRiRF754+XqbBcNUb2rZWwc6Uv/fmyQjjKRBCJV1td+KO5
zyHBmS3R38M6YyW4NvfeqUxIpnqzQPjFsnMbAQyNlb8my0UpXLVrOF7tq5x+MllBJ50dAwY9vjN3
CE0Ku0HihDALL6hAZF4fKTGXWL1DSSbN4DkBfPMt0aQyiEX+ECsHgVIJFFvqWAPCWAs6uE3ogNbQ
Qid0RJ/kaqvZtBjg1P2Eh2fhmb3Lc3Dmc3FOiS/98WrlsYsQXqw388l+LYvTB/jLUWRS/AMP5sKP
mOw8klzqtmCclibptKToSO8z1PwcCB+uyiQcJ3VLeUkBtX28B94m0Nh2HpMHmrvIsHKOo9VOOa9z
QTJiAP7j4MZvx4cPiw2nkCS+yFnz26Imo03OBX3U5czmK1oeksmw7FrvGhCNjl/hLBBronXxqGr5
Fy4yO7R0qp0321jpuifK6aEJc8WKne+o6DOoFMs8GqxuooiO2xuxSJcm+PgVoOlMF66XD6VS0dNi
YsiqI1DdgltIiDgmUb1Fn3qFH4R8mPspSjpr0jrpIxtkrl50e5sv1QVii2dYwRX0zdqZL7d93tVl
isaPjt46QFrZRxWQZWNED91/OD3uSxCNe6UKGxbGJvwI1La+y42WyOaPqdGVMPaogRRnx6QGgG3A
YJYjc7rALlL+wJXoCwfordVHQfq1O5KJ98rXHTH6opYHOL1JuUiLaCRJdMx/Hv2S9ipPMYhrOfn/
e/Oovz5YJ6NUZyBoocXcRsSah+3/QNAK9KtnOoi59Yd5vtCKHDJiHTkVkxgZmuXaSTTB3QMrVg4a
o9IRH3rjtUHVC55bpd6KJxM0I4m4iWk+RP5Fn7OeFnjjQI3kcjtbznvju/wue9TDTBFdXlViwXZn
pC0tlExabaA71Q7ixJXO262HLcLHqayMHibQK87clYV7cwqNmMyD6Feq419dswqPjvFz/ECFGdk0
PmxDrlLiSs2DQfZAc3kcE10RRewFLyCtwbrrOP7DdV5CyuWE7kKLgk2InF0iPeSo7HM88ThvNorR
8rde+Ce4gfZ47ziWFtE2wMRqc8UvwXLxdHwBQPUPLJzMkuVS1hUha7JqwFp9mlK/5GHMkWr7vCxF
FUdgRFcD5rp7Oj+uqMdl2sTCb4uY1ES2UnMvrDVisA85Heotq0Npc5qli3O2ID0W3wE92TKRUEe/
gxNRZYbVYERFGbMt7IVNDA5Lq4Q/APzg2S8H+pScT//fikIHk9GupKlYSuYXOGYpu4xw6a9/vKiw
H15wL75Jk9zehNLefkcSidlOJRzPHEsaE6xblq8fdjahWimDtx+wvrkyfWTeBsiT4h/+Y8NO9qnM
jvxv6gbjpCGRiv9hHDENXLQD/mz8vKLQnKnyXorf9buzGikvQkO3TX39Z3MMD1yI9H7mzg7jjVkQ
NNCtvUvPX2Zxym8u5Qa+AV/CDzYvbUGwYzNFr17kOhAFZCwmK4SlClFX4YEBdxCYgy5G9+PAlmmf
1pkK217YQUoOpGA76MvRd7fVNecNvdpc80Lf1tJsN4ogoYcDhwwWYX2bzUzgke0qfGJM47dnNLOY
OfmjXUQyJxcPZqsrD9zIgkhAbQou/gxfESp1VXrp/c6nzM+KF1bo8fMnTbWrDjcH4MOUjZ803Nrs
CBQJZAxf0l6+mMTfVNhTjijX1f8imOKSTqpKKhxchpUipEBaubFQz5GwBEKODkjNeCs05hNs1s64
Wu3u/vXgThYg0ybtsFwY4yengQ9f9ayCfj2NW7g5/pPYV5Q9kBmcJij85N5dUNdcqRDbqlfC51K1
XmXmA0NSvgszD6qMvs+bRso9mZjZlTI9rtAD4OFFuf+QGkZvpAdp9dZpm6pPGJsWH8kCwtcOh7Bk
Z4oA6V8ruRtHteDwCpJITfTjB2M2xzEnGm64ribHPR9vJYLxN5DQuDbsMpLlfpJ2LJtKkwb9VOp/
DBWEN1kLyGy235q9IaNTQc4IpRCRFtLz/tzZoJ6q2ubW1ccPco7QtUm3A4kvSr6l7jIb2fMQfZRo
a/4iQbtWIQGjmU7Fksy57XZEsXQDHfU66T4VnE7dVY+hIyEPa/9MmseFxBg7xwl2ypg6c1X1U1xV
oNscPFU8cvq9FVZZyTiEnBnHMXgMMSH4TIPSOYhdPmiimfbQpyMbwCRdPYm4i2wu3pjSPT0mC0aT
+TXfDDWjPJxjXh/JiRYg6lM4CtNX4tPe+ckfaqCpdiKRT8GDuIVtCZiRtB9mLRftw6STN8ie5WpW
UlP2NiZDs1eF02GQ+Tyoa3vWuYIMLqZROxszvzeaIWmlAalfgEmfcLjavPCCACpJ4FFO08fHhNpj
s/NZAo0P5ka8i9WavaMtjtCwoBneKuBgeh+oqTuAbO0m7AzrfSZsgSoxHGjstEh+lmTYNnVap/3K
NQjjtHCIJgP51KORvX75B3YUxooaZVHIbVIXFnNXUpbU+/wt90PV5x0gDkGXZ5T0BeU82dg+02jF
IndHdk0GN98gciy5kOjTSSEBKUBc6YEQd63pDYvD/IVU9qUdoIJMh7A69xbsYTbvdZr7b8Kur5ld
w7t59OQydJ4O6OrQQEGDGS3TSKyaU6cL6TBrP6hY+rwo4z07+2PgSJolNiP5jWVa9ld5AsoHCIzW
PnN2QtiBUa52rlgycJ7xpd2jo43hQ6vhL99wsaBFc61VbgiKrtsh+satOG7dwPVD1hVJNb1hw2QS
DjJqfK+7cUoyAlICim3ZQNnuAqk7+Txw9Rx5YW6XMSEKyxHDHavgHddqIbu21MXElS44aGzkfTVs
O0ayHnd1XPiF+n2B9REUaQc6McOTC6T3Vh46jVBARRPfA0YsCTV77283DhQ0zSYTuPWRpy2zyCp9
J6awLoQx5iIM1YzpUTrnr0Imyj93HEWqOFiJ5wEOktG+Kg6WeHzTrcnAgu89JwygXE7zW5StWl3D
yGrXaAw20CjqtiYpyg/vlv193XGx3qkHXDy2/G0C4SXVFAcgdAiuiwB2hPA67cN+3erXQpawfYsA
k91f4c7IPQ28Gg/XpscNK3M1wy3SJLk6c22X5aw0Qcnvh64RuSvct1S7eHlKMmNiTcjDhmvOcJ24
iI3vAfmPRC7MueEoY9A2hrLTZtMXuBgM6KQIxr1EKLR0OWhlyLbq+ybgDWTB73h6osc23Q0BaCF9
RwYyqfaNRXIYQkbsXnKiSnYTmq4imKXE9KJF20AV6yLnHg++Jou0ts0HP4HaaanbJES3dasfg6c2
DrwrQHnkvs9uNJ+iuvKj6E3501X5wKe3BX1pYbVYyhi5Mevl3iuY9x+c6FQsiTO8UN3in6N3ZWTO
jqY3Digh8UfeicGUW9bUL8IVyD6zNU6ZkN5QhivwJAwZOQWZm58UqHm5JxbPLTCRM91wThV5jz22
CZULAVwA9icq5Z5GdOPutlw+UryIkIIJzT/4dONoj3jo5oKv9WWSMuWuzoNSk4Rkp518/p8oY8Ry
2hBZqml0nH3bj5rjbLtbw6rLVJ5T3zyxjn0u0tY4aT3tO0JO8+bhwomY9COv4ev7QmCC7m5mwV2j
dSNepo1xCwvhG2bd6DVhF0BkBeY5htDvNKYnYCgvWT5OSpcmK0/aSOgsM9A7glO1aJJHCf9uvlYy
YQsb70prPxsY1FuoLG4ifFaEw8aIWy/pp0toU8s1Tfuu7FTSvoJYkrreSaPFKrObt6VVeTjlQg99
Y6X9mzsyGUsghZle6a33Dg13ikBy8EybU9KBTL3Ux6hJQ7CKxQnoCuLraQn7BYK847fe/mjEjTf4
yMu4JCdS+PTfXH2WZIDDvyhH/71B4XdjjxNZxd17QbBggazqc/bqoym2CeqYCSTS5PF6CwHyLlwr
MIQzZ3Eajkf5G/FQeHt4LLlJ4KIjaoPHk9vGHvX1pL7iNDHcDLy3Uuq1X5IBFHGnqLsBxPiRqtay
Rxk94gYMpjmqpOV45UIzXimgN9JB9XxVoA+oLHvgciNWWxZD+vsq5CFhDqhgguFUFeo25caiwIIK
KFn52O8eu8CwejYK2U01v1RhAE0BpENuWPtYHlRbTThTTZlePPs6GCxGvj6Im1IYX6ef+tYw/6jg
ZqMm7rkEkpxc86lQsLNb3EXAIfnm8KcawVgN42gpH0AcplR74p+NOR/KFVFBslMaU0WJYTqGCgra
fqTbw7RqWGNE46kbfNkB+No34y0u+aYw+4XCA7YzEkiJ1ZAQ/X08uTHfGYCknQYracJL6bgFYGbo
4NpeXRCczPxcCdgAiwzLsrcjPVJhgZpeNiWFkUO++Kk61XQPumb+JgfkiMlQs7udwkuU1A4M19JA
AGckyq214WHzHiy9KygWv+7JuSsYyNwKilfjLIgx817HKvwVQ78XpRiP7ZZQlo7lpBckWpjqO+IJ
T/VhqNsxwZucnbS8ROgTLRfJxW5805tBePKEx0lU6lFKp0HA+1vVmTZeX4C7S+AzJ1s7MSuDrWGF
tUO7XUtcO0W1XI8qQBq6CDjhseakIV5Vlm0A4o7Z6Yi7hf6LwoctgMPI+acmIEwCSs3pRoEXZGXO
E3YV1OWoIuS+np1f1CfRI4HscAZvyWw9+6vwSBNUYJV7jzl3orKwdrAERho+0RdowtNY4xWwst+9
wqMoRlo0td9FBXyXQMVSQ5binY+NGi7TM4C7cY7CDnRD0MwqvLp0j46YTrdlmsWgrjceaRlguDPu
2FaC1ziV05S8LdTAHoR5h5NgeVaLs8g5tTrIt5DzNfh0VJpr/mo/+w8w4o+4L0qNx61gQniuKlh3
Hss+cr46YRHLxFvQT98g10zJz9y5yltfSRhNM1brxojeSUKWOxQGC5iKax+Zv5TSGiMt2hS2vlld
JD9hH/ZbSglRVlv3SvO1FWffT6DZ6EE55PtK5A4wYWltZJ4G/lWoGQaAXWbNAxbuGvB5vRA2vppk
1PhhdI3ylNwNACoq+asdM6ztG5JkCfSbaODZYeUL76EDIajgVKA3gE/vSuiTys0hNCrR7xihqzUW
rjEgq1RcPFYecrXPmiy8koL855I/Otp1kg9dhA+LZur1+vNBGYFM4+ydnwS2RPn5a0qOJDnbYG0q
dfTiqsLzWl5Kds7MeLNq1S9ICB2wnD03E+v/ks7tui8bDHX/iAE1abdRrQWlrVr4UovuyyX9wuV+
VtXwIF8EKPMEauewWw8L+AiIa1Vhpjqr+EumD7l/rGHeD778ajkRHhZ7eWL6r/zDlLGsz/bKz3N2
63U/6F/KEWBW2hFimSL7F/CQZF+xcOhxcTa7gnqBwkXcI7eYhmT5w9zT1MYudwQ0KDDQdCy+Dgw3
k4Uj4jnbzdEqnS/FzshfMQGhKXEzBe54QvSkn10oCfCDOnCT5ZqfSvdib34PzJ5fk8DxobMUCT3N
Pkk2NYTXw/RcsyrWhmkSvgo3wh/7uyw/ZwedkoHXt8o7U+fG6/mq/Gyj2HSRkqmA1mXkIcnZ2iI8
PyUwof+b2ogr4oa0bxt12zw0JnBwb+LKqrIQ1kCPguoA4pcI6AyH/uXekcz8GVnzcvCRZPhwGS4x
4RvG+Q7KDtKOwcDTJNCvW6m0MeuiyU57NnkaDGxPrTcOyvfgezrK4hGl/Y4KUu08t8U71qLnl2w0
VjTz7TpGyC/QrkdrT2hLfog+b5qlEI6hyX5W/6X049HYew0WKRtXPQzY8labHf8kyMB14/AG6+d7
o3kq1wvbaVVUADKeBrxZstKKtF2tkeEFpBHJL1mi8dOGYoszstM+iVNg/KDYIkjDhTfbyxgRoznW
ETKXCGwvSdnbxB3nQP1s4A7lErY8g9qLDz5LuHYT4r/mUtJxhHOLQUc/xLVTF26o682wGS1DkNGD
Mul2qxU1UuT69fmiIQ3EvQ1StG6Vho/57TJZs5CAXUPI+onUqdIxU7DpPm5JGtS2BEhl6hcznOx/
Uwl2yR+KwK1byNi9LFmdqwIZ9ViN124V7fZKwBBKG02GvFjvNm9l/jLhKATkmyImFAO4BqWBBJuk
BRfSZpylzn4JVl6KBGCu3JJEQLHQrkX5Ls9cBBMQY0jTwJERb/MoMEukY3LfWzlihJv76SsAR0rq
VwopqqSaAtzJSStTqWufWjw7EhbFqOLLvEhnnU87hASXwVuUf/zLOo/52raI9eWzoSfuxXoJbp19
vHkhDuucCyky11c4EQb8fa86CqF2/N3NoYld6lbu9NrfULOSC59DfJ4J+zfjrfAHvBAFyI5n5LJJ
0gnh6UEKAnWs8B/n+tq0WnWUHmg2EqTsbGAMkDX4e/CYyLP1P47KiXNaGdJjVU+wdWewkIs4Vh2A
9AxA/lSqLHshWdviwKKILVGZkRYrD1jEhtlsc+Ryp2TSJ1bZjWcEk0jPuZ/21j0/auJP7pMJIEkh
C1rBXF3OJRU9irN10EIwF2prNKWlEugfkVaD251pqLGURr0l3MSUZTwD6zUh+afdR8GXgI8HuFj9
SPvwBtYYR++9wSv1a35odAeoL84KEY3vivtxg4NDwWzrckXle77I2oq2AzLGaKxWFuQ26zuX78b3
GDk1fGkPKtcTSOkNsiImQDhAlsYDsbzeOLEka3yaRoAnpeUTNxt5qVokWgGRLGTsLi6TIvCnRseN
Ip/TFpamgxSw3IGwqrmeyIh5N6hG4Pdr2Y24vwtCBFhZxFwwcQ8wWgUwBzGzVO43bM9GmG/tiT9E
liCKWUddBJmiAO50k8kutCmpHbY+kfZoF8mTmV+aNOLSCkrtnBZw8I/4IGo2nn1wssfV8Bl/u7zv
NQEORcaf/V880oxYa8wvZJ77HeTPyhiTEHNVZhJo4TI/vwAGeh1hxKi+cTZMLQJrOEPU/cFbLX01
ZTN870wcJr6iUlI/mfyKOxp8Li2mBY5gepIzDm7afLIt5Ti+kf+68ggOe/5O7pY1R7jD7zXhzfxR
U/V/Vdu6nWtSKVBtUBGeDo7c8+KUj2S9CfVcrResboLhXXRXPsN0R/REsVYmrufwISRfA6VHyVC0
9OLK9qdmxuWRTYazinyT935iWDNebCiQ5mWsMK3nMp0fRs1cqSLfInWcc5LX4t/+ntpL3tox+RlC
r0DC4SCtYgnNbjjsyyJtaIAiOtA0o7Ma51VvL1mcmQRN/ijdJutJtVqEyuJmrfgUDz0jAYtDmPSG
lZ5/FFKTqkE2qalVFjGYVcglQbwPV9i+DbaTCU+zuWXbc2oB+RSZSeNGn0D22JzzHsxfJYq7Rf2E
V0uAQyXHUf0btIedxyPnrCaB9bbQP2Cj4l6geumNHfe4mPlRIPxcNBjNDG++8p9rzPyBTIU1WEVP
KOq+WbFI5pyj4E/+ST2cBhGfTgN/yv3BRHc2zwnBKU5HkEFaNJKGaviBj5BXfAgRpvrtrNxC7lPh
5EkRcGzeEVjOjWF6+2hKuvMfyd5iyczVDj+tdTh4PMMFXRfhlVHOulPniOSTw0ZX+8uUryUvwWqS
0amxcYNgrounhyxm8SHKjsEayQP9eQIw1une8HVzdPd2L3Kp8BkM6/YqBIpo72WDe0yAtJXYmY2V
keQmdcSw+KfbpGQ0Pt9h2LiJs5VsSSL8gQKmbp6up39+LXgzJmYcxrqxn0N+CWilLhd8Zhcv2Uuu
LtD0mRbcwbdKVnDHEhaV2H217dTYv4E/JGC/rWjspXpP0KS26aiFX4lnI6bZ6jOit/co+9hJUE9Z
NaffMWJM90+yhb2rxSE/BIF79XMRo/Pkzy1+nXmZqh+vpvnalRov7xdv1rcyPRwadrR+rGE75Zmo
a6cNdlbZ6kLmY810g0n84LAUJ/KCku+CN0Qq22A1ilJERBYrqowVn6Guf5e0yUYDrfSQmCDlJ+Pg
6QwRp2QYZSdJj04N51vjhutxMZxnUuJMdCrIRsz5aMfHYsuZZ9jtuu6TTlPS+qz6Yfym7usvn10k
V9Z5n6M5MS15rCDRNwsrxapbe7epxFSxKSyRN9kF18gQM+rCuAbSWiNKQtckMtzhSm1rV0dWF2E6
40Q+kbdLWXYbJM6wi3ED9FbllNXG59Xub/o6w9/7jTf4u6xK2R8JnIeNMuEkjrKCxNDqxB0kSOvJ
v1DroV8DJv3U8w+s3q/ckDN0JHMZMN0Ee4l8Y8bJdFL5MH3UekcKzsseJeRgFZQfjPFK14TYMu1n
DgQlIkUXSHsBVfzGMBGFO2pcvledoCt1ZH2NZgBXZxVLqxKn6CsZZG0mHGJupsT9kP9AkZndQ9Mn
z6CvuRudAMjsk4hlmtCzoO61g4N1sPicU8vVA/evsQDn21fCsGcEBxg13FSPSiXk9F5pEQJwOJEy
oIY72HIU65bRuaPjAwXup+riizYX+zTG1jh7rEBQPdghgFxnju0IP8E7dOlL5v3oju5SbfdrVP1V
XUqZl/GvIAZHcTf37jQP5TEP9KK4OZSVPK6Q96hsQDDjBzPYa6PyNVgACnDL7H+mS/jT5IkngtBr
xa8XnVh1q7H77xQfSFMYWAQ3fYBNGJo9D1O3r3k4affuHQacWvTEl9AGFyLq072JpQLBnSXvz7XV
VEhstdPHKKb6J5nscrXNjcZugC/pVLe9TdIn2VAWYRidWKg0eJbGk8m2e7Zmg2VBjMyT/KTk+M9r
tmp/38zmWCH1vgPapVsskbU4HM+Wi4JAobhHQHnCcdEOLEdyR9UF+OezbLqA6z5MnA0NYVjhC1F6
G81dejMSZRonEqrjjkw6Nfu9sDbn0sxoWeob6ujnhtyqhpe2wcepK8L8Te4Np/sU1IVgoZvaLxSo
mAYZkcYOt7iYj6FaOp61dQNeG+Z9Zj+oGiLhBUYjW9KiC6XYnAN8ALnXtE2r4XKhxHjeFvygH//2
kek71qODBL6aQtMjmEbFfVNuZeE5EX/TZeCFEG+jgMt5DHzzWMnKUJ+VLkVnXY+FXkTVEEHVBdan
oS1DeQT2sdp7tpxqVecaXirrT6tW5PCyU6tngKpDCHExDHfT6UqEFA+80oY9UTl6tVv3O6KVuUwI
K4tOBtLHfiOyE/QFCT4brHxFp2fm3AlSmFfB6oiClJKt97pZ+QYjPtcaBW6QSCM+KNUfgvuGCAU/
JdHXl97b4rf9Jg31rQINUg4Kw3nPldKp0bAhru6bjyWoONx42NjaODWWNpiF/F/QAakLJjXaPWoz
TRLP1txgnQsurhVOXxbWtLfuida3AryLyfsZXzJ+O3Phdc5rP6ChjA1kqlvgsg/h9a8M/MbH7/oj
KLHGah2/kWibnhMPqwW5+cbZ9eHHc3o7op+kTo9BrTFtEdbA5YWa0VQ/dKX5Qp1vffIyLTsyC4B/
XPrdk39cOO9ypEUEPAv8BBlwnrpSFZkUP170agIfaHL4B1ydjZhXJ6EVj/kv981A3iGvaFt2OTCJ
Z2kMmb4B/LvHxvOd+fCxGMnj+AgaYVJHXk8YHMw3iSMuEUhgSUm7t3uAKRL9pyMzQ0a7RLmBUhv1
41jYifIvMri/ADrc+zkC2G+L5znbEcfXNumzHpTPOWlO6wLFwstjN+gCpv1+YrqwE1otTF+w7HWg
ADwxx7U/28Lj4iDi4VO+qAaPUyI0E0v6a/zpQiqowKi8yU20VVqAVK8UuFsI1hnoG9B3jKiEkyPH
Lr2tK9upSj0qDN36Zh38WJ/67onguAVKkZcHUzjUX8dwc0FK99TS3yIkXhcrbeAPfMUbsoHIn0fj
lLx31ltohDicgkosUzf/jmsjekWFmujVxxWkOyLZLy94XKDg1wcoqhguJbHxbUPRVcvGq8Otpgyg
Re1GJ1pQlPOzkH4RAIJfx1DJwkmiVP9ddGScENLNVIkIl6qz/m3SQgy7/k/WN15RzDFKQOugcyvk
SNSNpyEedk5sLtA1Fu1Kk5BfSBLt4EW1A1daIr22DzSGh1XE6mxaSgFtP1Y/g96jFGM2MGl+6T4h
VWiZbTUqfs2rV9HEdzzMDEAwK0scR0VT2CGU+mYhWe+qPhFa5KIjNvFULxoGGGRgXSi5aMEBVT2C
/V9Mjp8qHiO4z9KB8QWyXnDEjSXqitqNo/On9TgZ+GchB4D7s4wUJitcnSCdAbFK+D/pUDsn1371
4YLzU4QYHM6QPq+ge6yuglx6DV38yZm7AvLlAT1Zi0oC427iEx0iINCJsZ1kLerwqMh6LWrCVx4G
IXJXXyeFTtXMPnTmXYURYkeYeMJvI70r+y/LXY4xu1PkI/5yB836i40GVQkUE9ju+eQz6/E9el3c
zrg9gpZv/AS52spydgJiHtCvk88Tbul7d+HsAgQwJoP01Yz97RyPvNoUOPk5AvcJJJeXGmWPY++z
/oWhHCGTsClbSDJ1dIYLCpMyO691e7as2JkHgJ7PGtx2nDYI6rjxB5LqqTpDUpM+1QBVM/A98OZz
xWGQZyoJHL783HMzNlLOL9xMglQqc55tl8dkj6tsFteZ6gV/janbGByJ2h6KLkvRyNUpX94JAPM8
6ksSxjUvBHIMFfyjJa69L8iJ/FGgQeymFOD0BPRRnh4fTLQg47IOqrTDdchhrPmE8jXo7gq1KI1r
3ZSGpviRpK78ZzLAmRdqzkgAMSUGDZbFh13SNbF6pqGZwrGRZXCyJapwnrfBjB4pEV/raN0SDJy+
oY2rlzXh5jmO23/wNMCndM6/aSnkYkW45YD2/bcb4gJdbzk1KfKPxdHd0yF5FH+vBWRFiNXBLe4T
rWwJTTCdEKlaqk8X5YEwzGAD7Gjsa//1YSHpRyVFvky2bwL/bFu3KZqQKvLvf6rHuZknJ4V+gNYW
Oixv22nM/FDGmzle9t1OHgeJhSTsK0EqnzkVnlk84YTSIYTVp2yBIJvV/7IyCs0uPOZBMV3KszjM
1tzmYtXxjpye7vvSoc7AnZNr9BAtA20zzxZ+51UwBlI2bDinh0l5+XZaJWrSL8iwFxDvxDG/3do2
Kt64Js29qwP1ANgE72LEMqECvjICF3OJ0dFkRZWwSuEzbRfCinRGuIIe1C+jFYhe8uDelPbUvMTv
fjXgLmTBPdQlsCyFYzDTQ4WAkHUrAJsOgePvvI1Q8bUzJg6hVPFMOQsOPgRRGyewZ2+CndVFfE31
5/KRgYwD8sDdJLYbTaOg3AFKIDf+4UCWHAdZKQD0ev38p/0dixoKAbd1qA6C7AQBBC50zUr0YceA
3xzLiBSuyug3Egatpi8D/7MWLltbz0fFIOB2N2h7bKItJnOjuPVkR8vLEN1MuVFf54YUIFuLCWZb
HUaW5eQ1nVmJ52w3Ah+YjZM1HSt2RbhN43S1mfjx6ucZKspNJDFpqmMB4u7kJ3Qm7JNBWc+A6diD
/3hvMPoWtRFvt6us278NfExDDRDUS9YZm/75Y9fpMaC2YVTNrduniVs8Vz2r1OiC1reMEPLVMsYK
k7+Kuiw+nhmJeDgWK3FjMQe+WOoKCJli4vPREq9kPkanK3oKIrzWtgD3m6vP0SwsMUfLrrFKnZiM
hwHpnK5iXtWFtb/6f78BQTSbMbFo5jdcn5jWyUoeEeC0uCb8WvNpKuCwgchNFDNdI6od9WsPglEs
u16ZHR3a1NuQvOHAogf7rBs8ia/2rZaJJOUoP2s7zo/U2bRQMiIRK7iqtCQacgTvl+0UXk5dB4OI
rmCQsxsqDJoseaRdyZ/lGwbHya0DzBv6ztV9RhTWYyM5SyrroaNvZpBA8uw7SVRmClrXQZMQU8Px
p0gY+lGqrTCp5SPqCCbuHO5ft+g8TZJS+lOlz0iwfyZ94yY8uEfDvapk94v3bYrtmc/xVwNRurLg
zLHG9DFU/OoMB5J83utSak+7hqBElaHtUQ/YBS/W8k3V2EilREdz6zdTufDdP+YSX5Q0EE81i4nj
xgIaynL84y6p4hmX6G/6bRI0Y87+tuGSMqaqjhObqhcFlaHw/QM1unazHomsTK+2fXXWf5uA9kq+
cx0R8FMIqm32C4XDQ55XYv/tE2azFG6VAP9LD6aZiAgwGOQFbaWHAyv4kk0FBu6yNUiXn/ISP4fK
X00ei+osghiNnxYIdxmz6jfxHkQ1GwgaU48eHxHM/c0djZu8NNlFHwdNfrh6F+zXmxhOuVG0XJZJ
iMDTurQkC8iN+1iYiAcw01S6OQPZcwpfNq6BYRaz7dekg3TEuk+3LDc+JTJ6bNgOFVhBim7KlxxT
cMcq4uUyABhyhad3fohvvLQhRfmp5+HwcbBCoHm9NEXyZF/5fX6eTEV+Xyw784yetv7QRfJZhgMO
Ti9kv3JX2Cg74WDVVQHIgLuGueR92DNw9HNOCWmKonVKgsiFOgyK2Jtt+rQkBtlmCx2bZu9hdawK
w0ISMfulbfqNryUXIyE1REmndTFDMkWFsViZEnxSwrMnRlg4DUSOUj5Lw/AHwzbSt07OVcXZUWc7
CZSxJPSXo4CxNRQXtZeOrfzuxFU14/Q5M2UfnYBIzFohAc0x6Vwy//tzNCiLErn2pPhhePvleZfN
Sjk3zbxRwKnaEFrGHR6IhMIFvWBhLXWjepj+rQYNRvg+PPTttuoHpAan0Ptwx8mGy3cTVBGeqUPu
FWUEx6YyCLGZLGOToIlGCkln9HueVPaORgZKI+JFpCzDDMLET3g5jHPrLWna4POF4vAKY1FVcIL4
y5mcUsn13cuSGXZZHB8XQhLgzqxMN/Z385s43KVMz4u3SvyGxiEIr7I8orJkOYyZu5IoYT7KVV1z
HjE19zZnsqFuqnVvuh7+gEQKegDBUgYE9q89CLjYhET89MidlkLUAeJk+8OGMascroNq692sAdvg
vph7lVseapXuKBVCOfxBI4TshZTffgoGMFqEJ1/9viVxMgUIpxG6rJKeXAuAAesDbJcdQQigqCMT
6mT4ncbX7teVYI7UFzPToN5banmeGEKEyS/NkcsH1oPPEmwovT6OY8EnqaNk65rN2QdUl43aZ0na
R9ughRqdlti/P36hGPMSACLI0U3MijGtS3qt83WcIstEGgXE2m6j6HPf4S9ZHuxvaZyk14rKvc8y
YJYR9i/QZeAlFV73nVIeJl57hzw1blowhi9meP+vcjKtEHovUxCm2ZNDdOqXvtr5AwB/Oy0ojtTd
J0grtodSpTc9Or7DoZvxwFwnMJauCG7Nu8hLgISGHm1Ghllaf1cPZGjDiCOe57iXAmGu+haMMKy5
XyCApAkXtO/zGu40aZtvbzW4QHHSLdBzK4hgL0YCKxN20kXxrtv16b8lWPk+ptlHFwkE7dZOrL9G
bJukIVOQS9oymkdZofUS3VRPMPZjwhd20mpMv5dk+iqsq1+iahw9btIsqG0uB64adbsV8vMmKwwx
bHbdBAozj6TJY5zrWdm1VKLTTf+vWU3NC6jMcHWsNcEc3CyQDvj8GbRE5GSLxtj5rNSICwwNHjOl
XT3AdQ5mT3LIpqTyqlRo+nK8skWq9zIpuh74va+m/j5E9+S5bmAHXsJsfFThK832qgfWeybS8Krc
zdn5utShR9PwDPd9rQ9+VoCsxhAs9DCPOPatZLjZjSskCXuFao2Q25r7Yq885sMA4S4FaXWVNBA8
goPcBlqGnDmv6731B3LopqGgCK2JjyAJ2e46YvcjdXhqUH7k+DxobSjNJ6+0aTgJFQ09btzvYoRN
IqNcIdjyYvuqtIQD41XdMv+H51zrwZuqP9BAmJ+TGxtGhWpDIV7FRprJBFP9u3x/rIsoZ8uhgX/y
8f8wtk0+Ck7z/DM4mgiLzrP9Ip9RX7TpbdlZSXGhebFu3CDJhd5yHwhkwjkW2y0/YTG9jNI7AZWl
avjjGRwdhBqAUvAcKafFXow/Q2gaGwEWDn/82QqI2J99qEhRTaMtHDJkEl5v/YTThNQAT6Pz1SgZ
O2T8Gv10hO8o+vNbhrSimbBU8A+OjhM2N/71iTkJhZuGRNf4ATUVFhhBWlpL9rM6d9aJLhW7GqP+
wO2YFQta+7QwbMCkgPEpAhmegKzvInctPmNJTj2yWPGCcrbq46mWhM2R2qGiSRBs9tZKP4a78X/p
UrgcInpAybGBvm3/mdTWG1R/GCM8tukVLlXH4J4GmS6hPNfQhjta29I56r5M3SVKqG372QZ28D1w
qZsszKQbBlE1ES6rvkjEu1DjfCR9H5/1l6l8T+mk/AcT/jGRh+W4VHdEoWkhlHvIX34DxfakSAMl
Rj9DO7lnwMe3smYNX2IKehlCHQe6GIGeXDFg+M/IJ7G6Z6mooewQZNwtsUZaZjD5+T5D1w6iMFCA
9MYmcKWLW5zOw/T32Scmp0ZbzhncaRmC3VJ7HBzRjKVJTytXRwqcjxuCWqyKooO0hj8k3bIwruWR
lFj8L1qfefNAInyDf/7xt51YJ7htvpXdyMxIgAv/7ggkMpjCqK6Rqoid6Z17eGcn8m0Udai/0Rk1
7D3ASQWwRYSJF1qon5n9YkDCI1oLFrvBeWxLjiwcGApkbBx0z87VUWt+bG/otTihLq3WSYZ+W8n2
gcitC9AeBDlSfinbgjzqKOK68+scQIZbXbNhkqzo0tVUGOsY5OzasnOJeQrG46Nab3MrK/dHAtU+
+ebgDS8ZslbXw3iPm8C0FsAJYCEuy80QOo+ezva28qoYjnZTovpm+4Nuxf8IB3uC/HUDmQFOHW75
VdUjYxICej0J0OkD4p4oj24LXeBHxxMBG1IsRRo/E7abBWbo016Q3icC8VRaHv1uWGf7CdHdKH7G
fCy+ew+kVsw811uxtqmW9WmrcLgRusMfM8jPGiOrXWrly+4NKUwIV5lh7OFXMnAf86uGgw/Sd5gq
Gs8tn6UJ8GVMi8f2lx/1O+YuzoPcBVdHeoeUst0Qa/mCGZXn738UKVjYhTNLVyOgVZ58W8V8oJq8
Nf0MxMvRFej5je+0QcuTd/yuiSlzBKNknjPQBih2sqWl0Mx3E5/S0slVvxaYJmPp9IhYtB7Teu5Q
52Gk2Vz8DNhx9cbp0Hfiy5BivWDYWz7WpVXdEp66CFChGX4IvH6QsRCfLOPhAr5EkK2SVgjtRVqt
mae7dmxUFVDHARIV9LP+3yVJFbyar4YLhjjoTPbzbpqwwWrvz+Qrj7yldHRffqybVcIt2s03VwWH
VHvQ5l7Fo/zTmotkvRfh/Pi9ETBmldGZOv8huJY1c8ODvkMqNEMNGiaJ8nobNlN3L1cp1HB5JELg
OdVjeo8hF9x4ggrQl3z89PDqQ2sSg+ci2qwar7xr1CfKqSSwg6i5UCLPpGIhs7QLQT552k19SN3z
V5c01f+QfVUKlPcc9BsMUiRCfXxO0K1y5ii1OcWcJtCYpwFx7aWWAaLLhH2FjhOive7y3lMkq6t8
nKFLIcdxW2vaEqCIKXWCSARyqclmttmdcCUyi5BEo+s+jj5oraL3/+Hkm/OeSLRj/gkJ2Q7RFHKI
cCg8zBI2+hhnr3qsLMg8b8Cjcs/OLx8/CaOHaI0qccalqoJxoeY9o0YvDjd54/V4gq83FOpAr3rY
KuEiFLk8j72iQp2MyqDxAh11v1/x35DP5VYNY0BLNCz8tHyY2rCWSEqSjR/abtQyJyE+Q5uWVqNq
2J9TtnTtsOFR64Y9tc6sIhyQjtfs0eTv10VTRD1vnOnfWVaoXqdY7OfGSISRInP6gwvc9dmXHiHw
ajRGo1cKYPOoGyOON6zGHCz0/1tUGh3sUSZ+uf/aCrnAeLc+cEBSinUQL0Jh73APH7+a5EhY+1qb
KRwvJQBdRKJJ6oBxcO4J2LOZJrBqz8al/aqcczkZZDKF9sCTnC4GHQdPG+nwGYRacnKgGwAKomI0
Set21lla/EeEw9WGhGXLr8w9B5XWDlJ+r87WhaHbtSmB8/yj7nVcFbLcubqj/hMhJhzOCq3HhhiK
kXXgg48DaEcq4nzp0qInQxYAULrkM4bj4liB/GF/buiOw/pJoy3S74FZKog4Bj2DHQdR2ub/XHpc
XDwzAbszuwyo+gGdIEzG/PINUCvwIGCR9zXYSeV3PPrl5KPy5B1veHcGDaSQTksFgoJHGBeRwxJF
QOW4AhVQKY/Kgh5KeQ+hOYFxhMhIWBaHVBUeh/V2JIfQ8iPUz6TnwPgWHfIuapFFFDv+gj+aNzP1
9wYpRe1Xmk1PiqlMkuwmDq//zhYIP35JH2APJQJsa3ghDm8k00m5xY2sJOoDJTS0yLXaaEbAtkAp
NyW9W1pWa5XKVqnHa7mWD7ltgDJ7ClHM+EPXf4MCEdg+w1qbG3J6WxcHOyHjQHhj2aXM81M9+UVF
6vEkMOPwvhSBPCjHLnYAzS3aJ1dhBUbNEhHspYfDsKTvlJoRWaeIV8CIxY/BNC09+nkIMgIeHBub
FmsXLYVIsEW27xT3HiEVnQKBSVCqkP9eL/1TKMkmCoR7fvJtYL1fU+cKl0FzRlkvD5Nwgu9YyFS3
mq4ZPr0KHzPbqgXs6ZSibRd0EFIyzfBuCJ1eWUiOY1XjGu86fByPdslPvZGFijkP/+IKJwaZaTzB
Dvtw1L9WKttm2/kIIRWArL9NiBQZMf9IBW34JwgciHzJnXbS6uKUbLeY9XGw0UMLNqXEMlN0AIbv
SJ0NrzPt7nqgTKtxpnQ4vR0acDFeF/RwhXpl+f/6rDzXIBf0kcMlgEMvcLDyE9B9ruTryQRK14CA
jveRH3oXld1cwd1kJ7k5J3utXLHKN5br8gUPdDPIDuwTfWLtFeU06ceEvAdUrDHxMNJE0t7C1Hzv
lWSnsxPi8AxRWp0KDIXNd4RCkBsMeAv0fC5fRNDZT8EArJH8PMtEEpMhZfDA5gVWaNEtPq5VUHPX
1VsXdJqiAF3f2Zj+G4cYHBv3U+2I8PgFjJXr56K43rZx4SI5PnffUwnpuWqeIViTienzd9gjNbSJ
i2EHRbn4vTvyvZ1enOmVFT0gpEE7SU6/EgacYRAJy7zMJWTMqpwIdQa/MV4Z92LRgQ/7yf1WUqJF
cGh9itii6BfLxDIUoNs+4F817NpZ66jKM9N/7ubrcsosvRCDmg8elwzR6l+45fsvJibj39hW0K4c
NXvZelHPotw1wrjaALcJ85rZfuClbv+PP3xugh7bYBQ0VGVKD1lP7qm/YM80pAOcXEfS1iD7MKgZ
f/DMhPN+cMfVZlKaUUiI6siKHDZRYq5tjJ9HrdQz/xAnuH5oVtRmQaEYaJrI+E5I2DsOfaUCVql4
dZCqbuX45NMME9lh29oqYn7wFeCPXL+fiUGCOCeeJ9fNiE8rJFV23p6O2bB4aSjtWTk9jiJJ2RrL
yU83NhaAsrnHHS/WGOltDqn4unVOyBex5GZV6uaQx5tZciIIVwa3U9HQYyBWxXhChQNcfJmmlyHF
n7/ufmRutFUIeiOhzcsSm9fAcr6nSAsY3I+SryrhGQPBTRNbWA8sEmisgU8ZQL56nKq/6SQnfIIS
KHZLwPANtzHMK6Sb1+r5Z7uEEK1zf0BbzMV4a823ARpz0Vn8ST6ZDG3o5gUjqIlNmFKr4FaSfBFa
JOUtLHh5DaVKnOAJAAJ//xTb8yho4VdkB2gdmoEgua6zR54oIJ+ncbqoZZeHm+nqo+gBLxwI37EM
uJ/6wUCRDlMpgycwhQyWeiSEwvUl8G3vAEp2g+m8jflx6C+T88dap5Ru/V+uBjJISxQV4TeUBx0z
TaUf8ExRfM/sEPU+11hrjs1VZOTF/zGy02LFCqbbWrwEQSYfaXLJ7bJ1NRXtaFSl06Aub7trO9Os
8V93aGzgxvu2VkQ9ztY/fgMaei99WFm6paUIT6jkdvm7UY70oLh7h0ToL3/22ZosCXydWIpuWhZt
PJaEoeuK1BxhmPr9/zWkD0ERPTyxt9yliJe3tl1jFB7ydBwe6qOt+Wu8EFB6QFTql1n7Wi8Uzfs2
/vcTV0STwre/cjQqUXrSHyB7Oh5HL7Ot6UFPibk6jRGGc9vWjnVkH6wQfq2C90VCaZjZRbQyepiD
XS9Uy+kbpXq2B/WwQ50tOmf/QiKhXskLU/kCLwM8gjCNQcWuuUwpzn9PNnFalCvIlnodfC+99D4G
Ws267372NFaSTyQyKG2cVO/TeNpPi4xvHx4VCZU5r+1WQDsd4Dvc3VhWJc/MqsCKNrWV8+XrC7Z+
Zz+1T8cHAD47Kve5WyQgzEgDyzevAKf7K6gQ72hTvCdKIFjkQVVwTucUW+D0oiJHKuqauS4qIXtE
jNGNbJz65RPjQrLSxbquBTRkC41B0QVnTQM+JqVRH1apLOyogNtKMLKR214wDzZikc7ApI2yPlUR
o73Q6gwMVY8lh2m9HvGPMgzF5zABqTK3HYt6agBdgL9b1LOAJ3CcHas9jlF9I/+/aQWF5rtkoq03
Q3r+vWHYUCHMNbH5M1qByno8gbbKVWLYGQ92G1N7hMWx1HdeoWFiGoDpKsfEQt1fDztiz8Oo0T4A
HvZRXiwVe3I5FM576Dh/4/AwHuP2+uwQG7T6zM0dyvIxKFDgu+oUdvYK00DDqWzR8HsSigddomCL
gwdVaVza4mdQ1xzoyKi/TxWjiZG6KUMn5WD4NKi7Npah/m+sPZPRxGDf+WywspNClwEYui6vL5iU
YCG7i9Zw88yLNbjYpL0kHYIrmwhnuD+t/mJoyCrZ7yXz1iY1nWB7YktjB2XL9hBRL91sN0xlq4l4
RfWZl0ZrnuGR9PKyyDazQZZ6L2mefgxUykgsvJtgR3fL/zEjcZxdLVVKiQiXVx9SeauhYxoS5b+8
4GgmzVPRVwk6h6i+0eg2NVNHin6j2Hwk4V66b+Y0Htbh+3+ZSUKcAgwMihoDVpX3WK+nzeJ//yz9
FnX/+kM6S0lgVczQTYKr0Dj1cn2kmXBxvRq9JPw7pBNI4bBkRXAsoqLMGQg44X0TxgwdiPv6g2Ir
irZ3sDzdBmdruFjkUB45q7LWlzx3ARJaOnp1/Rr8XwrLslREdLnYd2YVBjhbpevXYP6s5/+HpOQ8
tJYFV9rBK9cMV/uQpFx/DjU3+0ug/J6QhoCnxEMo2gdSZEZPYpWufxPH0GjZmdL8samm0o9Wc1oj
hsMl52kCtPyU/lB2heGQcEiX1pH8nj5dgvFffl2EIm/Csh1Q11nFv/8GWJx/DQbrCHG+n7Q441AS
Fn6AyB+C6phTcTbzVvVZnllT+CaItbr36P4wJWiloVlj87N46SEk13EmKKM+HGx5d63Zgw3IbI29
gRWrfckbk2j8JZS8FlHvL/0oP4R36DSATR2tTh65ATlfHLVBdlinLdtjcA66cLozhpE8WPxRD2D/
ErVLrykyTWBsLISJFPgPSgdSF49JLPxyZ8RuSoYsBq+kMqMNZvrp5/SHEcrHSB9AkGpjdwif9kCK
jKl1uhaLWjuxAni1GFPVBgANtzA5hdNF7O0J1p0AbCaL7pkfxsbSIRBSRYTuSLsk0h0yO4Z+Fe73
szcPfmHWHvi+7tuq9VmCaBHfICG/JMnwXCG3vw87hRzsIz8s6HrhL41Srqwx74Cyct6/qAuVF0dH
2eaIzHUFA8JxHVI5cVGVUhCas6MPxpdAMlgDP3E4m0Wmpx0SVhIZGq5XNKoOGvvce/s38SLZ//FD
26byYczuYuamCmLfrJ58iBfsjQ4xQG313ylA+zolamWDzkIk7tOepf83SPiqXWPlGhxfuMAFjs+g
0iG8E/1teYJyRVwZrxYYaTRQVRWmBwRo1zAX1LvS4AnwKdTCi0Q1waayURUuqk+SSOjIxXyLxlfH
LrHrSx1YIu2U/Wp3GLPhGtzR777hFpwukPYFr5D7Xaem5DJT3Z21ODmQaQFAHd3SgR4OzcqoSke9
DP8OsqTu/0/28B0duzo0fZZfM4LDQxtdx0PK9jOggkbfCcKAjIUYWTMl9z6Hcwi+4giUyqHIdojR
VFoDYAtOhwBC229vMgLMIJewKqBfROgSRnJn9X1Y1IJSNEMKuCxpBZUIN3IJvBhqhNeuZmJQjuVH
mAnZ8d4i4Rx0fS+Bg+HMkDQARZCBCAh5fQPo8fj0ymoUZMrHxFNGkd6ypSI0JOD1AImE1anBZYcc
qNHAqioPYO1m/MonqtNEoOyRFYXkZaSfQkwpq2XAldO6T5VEVFqCwUEjQesOY00l3qprhVhsUNQF
RtucZ9QpCiZGKITMcgt1ht41455i6g3jhN7YncnFCrlmIBPzP/y66p0ghKuW7Tg8KAiw+MoULQ4S
48ggOjazepuWprweb1PPfO88xNJ8KkOAEslr9UBKxhsi+UXReDlR9c//Ggdra3hE3piZDYy1EImC
ISaWR1nZ/hGXaQX7DUyOSKuXMd9d7OoQlUldpjtElCO2ya9HUZ23oozeKKG4e5EcTEKemCYjUrCd
ZOljBvG7S4F++PWhmyTFnnmfPakS6yCFsCaRbR6RJA6VnyoBpju7u7tdwRHoikVWqU7seOaVPt6V
HJ9Hj+n0EYtsU4T/CZzXGWNuzXrvq5xvvsT37J1w06CboO3a1ZUgLS4a/VmtSj+XPR8IatQxiTs4
v8tRSJT4M3ryPbg4yUjRdMksbIZ8PXU+RMvDVMkTnkXrcDki31PnKSwZbeF4kOb8Q4KHiXtnbrE9
9naGFfP/xKCccdntlIHSICh743RnMQmQcnfqhvGpp2NJ0hC9dUA5gGiMqDt8EkdvQWnJ1zutGFg0
CjLcANiDHPi44KuPk0MFmAmSg+BYnaRcqQG36mJ9qa9LLYrI7TsHWRTSrvK9OMrzypxvZ472ioSQ
lirDPMyMLjHBKLhvSrNJduP/lbE3YTE1ww3IyElQl/nK9cdnevRVDHlx6Kw0N1xNxqfmM8SvZ1yB
4c3yMH7BOSWuL2Ccl1JZoRHBwbvGoC/b5J//eAtxjb+SKZS/U72OjklXNuD7oFzxtQj5vsizb+vC
rPgAL0pY8T6AOxCkrHG9E0Mo5HU6/GbnwIS9AeIVLg/dSxjZEDSUao5zJd1fzMIumMiKX1lxGkgP
ExGIhSCB0zyb8RmeXH2fhHuWI7JR/dFV7AFOINXBJiBz3EbBgthEdMYtEEEyvV2q7ewdma6j03Pw
Vs/9p9cgDc0wFWRug7JLAeJRUpOGWkUipxt4H74QmwI1f8+j4ApUXhYJqcgNiX0mBpZ7hHE3h6E7
sqGQtwhxYRI4HaXO5dR0ztvmFC9tuHed8hckCQQgQFVpvP8kXYO/lq+QPZ6v1EaxdsGgTPpIemep
B8bErExer2H5wtT1TUZDtBQ8x/ZX8dyiDjQuy9gZoNpWfuilXD/4yu+rSXk1/3PStZEqGAjOPwTW
90KvxFibU0Fk/hEYBKDPiVqdbDtaHXVW3LwcLRtTVpX5yrM1W3QU/Vu0OTGqltaHY1CfsD5ByOAZ
yK+2hHZemCorY6ikOsKnjTA32ArYlS7pt1lfFREsTcDzbU6rtv24Clkp0RZqdpjGItDO2/1ruyH1
bMB2rze2WlYDiDiofBc6bURau6U7ApeBIZcmT6FDN2dDqqt8nKc+7f1rzpQMdmzkjk0xOqdTD+cK
rkPhsNAvYtGEs0qvAwdTmnCP+d8olzTF4tfJLVwTjmc9QxQsnHLn6G+Zpn0nOK4PYAm6QYBTW2hn
7jeI4igCaRK19mwoSIp/HccmKsxcVz+Kw9fW4hOVXjQ2P2xINRH3BCtuDnWOX02zgVg78F5ZIzDx
15ODq1IQ6JEu+Z6r0HNjgQgoJsTaAsrg0lp4zw8Pq2Z2ja7hiO54/1Snk2gqlON9hvt2zqKvcYhx
Uh6yR8X/Etdg7YTMDX6l2XBUqm6q9jc9hcfysQBaPnDHrR+3xg5OZ32My/mh5yRQ3+x/GJeD0Z6U
Hu/ZGNvfnYtu2cIppA4A1zA3UGWCL++5Wo8NeLRlgakKqR0+GUIlpRKopFm9mtxHqAARlnZnubtI
ogYHSPRfrx1Nw8F7I1xBLJN4nUBQR/qgQfctVYBBXB0PjiNIM9ZsSUW71S3xOc0o6OzOI4cwHM9Q
r+WL+eYjQ3eZYfUY2dkaukGCoUNYHPb/jPT/7ySBfTbqOkmIWhqHTyezQnE9jJIoXtY8eODNRp0k
fnDAlVFNjPGJELDuK1xkI2b2e/tbw6PvnxDJ/Ts4ssTWjjA0YRLJRJ2wHz+nIylNntiD/oLpLHiy
aEqixl03TwZwn06UnPxJhsqcaGLlyHKfRHNQAiKl3y/icnrY0E5Jgqaqtb6F+sjHUe+DczxKk9o+
a8Ex/aM1itVW2omgetCD9uxCTBcgwuYqDTyFJLq4rmi66cXmNYySioc4kdxHy64NrXQNFtEOQFjp
5KdX+0TTcRDB5iQR2Z4TGCCRSsXWlqV9vwyrXxbAqdOGC/dppCXiIgCB+vSCyjOAmtjgASYbusXb
bw0zID5HxRfsdS/RkJpau2GD0tUJ97CFKNnGqeEJKMos+xo7m3Iq+pzBF09Qrlv1kofEtZ3Oj7Bl
VvfabPcJGqx2Nbs/66kccZ3T7Zf5QfSHOAtChYOAteHBk+NxZ2WBG/lt1krYOb0EyRJSM8PUd8zV
t3eEMTQtIbSMhUxUbcI9xxYsyH0Ey+XXLxwVOwt91IsBxLslUS3nfX2vcwQTseWLmRhx9KGL4Ctl
a4WmN1F58wyaGTCt2SFnrdEmPLVOyDxPeCGc7vEWnM7lCJCRHWonn5Am8GjmVWTzzgztUfSVO6CJ
YCliVXl9IxEx/XanStNz4TsJ1SZ6o9zrpxuOMWHwPO2A6e+feD8VMMT+e3713qr9KOSHxzR5tSe0
ucdz1yDqNdMYx6nbnb1l/a5zh6p5+O4d5dpTtoefK9UXMru9lUCET7ebyujpPYr89EQPT+R4yAtL
+OAeZ+2p3oSUcTgGfH6qdfRBtoDoUhmmekYXFOAwlcbjiBjI89wbhkq8Pf6P1C7miqlXj3U9ds7a
CsM5KWUxjhJeCjLO2SlcuqDIxUpX9sPee0yhBLvTqDVq2+o86CcDmHQIl5HZHGgIp8KJtAsSBVdL
TZ00Sr2FDx6W7w0KHnAjZZpONO6Vv76oEoXWm10cqoaT/Acp/AoTx7uVk1YdtUMi+pCpNft6Q42c
CPSo3beKhyiQD47qbjk1yInj6oCL9l9Au2XrXW917vuflb1ivLnv/QxWGG8aLEGFLwRj9KtrZ5Yj
knqUPa6hh2YJ12Plo+qMEyAAWOL505Gwn6/WAnwjVG30A7r9RS3PWRTgXFfQgO5Cy1xgHgM1Tfxh
zkTo3CMW3z0hn2LxFlgCCcnEnADZbz/ugeCV7ZWyvDrurbgtjDlUetB5ZMykXGSOsTe4sgYRL5hY
aGpQXh6jOAP0qJcVtVOT5fUhAQ9PP/6FG4H8NRTHfO5eGP9+L9lqok3t1mV7XAJzyYWlE8pncyXa
h8maPjZCb7f2omyiZEAZH4twDPw3hYwXDsLbrZVlqQe9dj36lOHNU3dyw6ba0A5CJFSrG8qejz9z
qMlbv7bre4PTetMgg91rIsCxbfwHPhtoCgLShvyJ2NGA0Lq2WDMXnEhVBUDzH8c3Kydk+xAMNI2i
w3QIaQJ9J/Y89nywxOxTIsvX4q7tfUegnhB6yIplXUCO+7qj9dFY9RXsAqg7R4NtpynzRezhqV7N
C+EIhpaOZbR4bzFSfa7CdzLBLfVwmQUCEINBx47ErkuVksK0ub+PKblYtFc9+td3VgfS5A52i26G
FiYL0OWDWK0LiVf1D9Fbpcnq7cAwj5MZwrf0T9FzIzuoTa7/l9gJWKm6YHpWmOUNyP+M/m+m8nVn
hc5tQXGYJAb+N/k1dEWrNTbEDm2xtjG+5hMvNyQqhpNUIJv5VYrewKtgx4hv4toLeWsL77yrLuGt
CGR2ddhArZE064YRBpny9DFFsa2w2vNsBNWHb/mOfTHRdsgCZochzkmRLlWWa8Nt59a4VrYrJ2eL
AKoK/16EWvex5D33PO56wap4Ynv573uV48grqShXzOILxzJhsz6zKRoQK+0pPmiZ2mAZz74WN2HQ
iin04IaSPoPnYzu5BIOz5kH7fXGFLHf9EnMlw6A1RirQS71qCkfqqc4BLafVqxUeOztqaD+CQ0+F
LCGpIsdCyCXFbjw+F0Tz6GGhdCeEtv+D0igaEA5tVHOIJkUZVT6ZTY495w0wi2+0zRrYU71S1yPe
GdP3aoGjV09dfbs6VtPLVx6DVzKqkVVgWAYai6C82eDBaHnUnYDOqmTFyGfKCXEneKRJNqNLt1Sx
xFJ1FsUulHpZTzZRQAfGk3MyBT8zVnHru/VqVFWBEZX6Eniy4JojhJaYZEYAy+fs9EnNk2/+a4ca
iNvEgCCIXjBFhH8KjRYtW+kpDcns8PzSxlApZqj4XMeXOEMY8ihu8SD/IsUxx5hkDjZcWMR52k6w
WDtE7EU4fScB3sxUZ+YSqCDOqLS033xs8pOu3zTEVug/sMHjT7iwsANdJdp+f5Fz0MHXy2tEWG88
iIwxjh3BOkGcGcjNlBPyVWKSMiDbncC5vWd0gdQb3GCzzjLZP/OIcCQPSgGX8ipRbXjlwliFK4eS
KeGgMjfdBbTxNfkIremkd2KYEtLjDPpjaPvr3bkIIOiFWMCPFOzjvuTobxzk/4QUTq8GzAyJWm/u
sa7sfbJ0SFa0RC6Hz9p8kYnsHo1OFH1YCPJknN42/t5IsaARLGpiuDh5T5lg/TOoK1pEwENHtVbP
ccKc+x0d2Zbad4uqJC6B9f2Fszvl58wWUnKUr1Bl1ObLc9WORmq8fhGQ7h5GNp2ntj63q6byAgEm
7clNnNAXYRih/TEB4ajrscMXDbUMkNu9NwiFb+SVOTEm2GpDLJ3v1I1+3fnocbTXF/QtN6Y9yPZf
KMUsFnqMdLYZg+fZTRaVl0oUV6fH0g9+JiNekUy1PAXKx2oJk/1+h/JTZpX35kmGgqiWZGtDrdtW
BQwsjnxWiG0idUWlimogzsg9z5Xpo2QudYsZGtGVPQLFRybdV/+MrTsdaeBPQ4fhe5Dvp9Lii9v3
w7WbCvrbVdz+SfpZUWXQXnSq/hYVy8okPi6i87212pTaeaRm0ImcDPy1RsAqZba1tuxXTZcq9N2q
I70c18hl6zCRf39RQ7yOi8m71VS0mekJ0lC/73KPHUAs5SvxrETinoVaz1HbUS03yuphTszuPDLU
JtdWRGctpPfQ7hqzon93q9ec0NzeVlcr5pZfKagNSpJ2B/c1gwHHVrCFoVzNX3VHlUljDK8cm4Jm
dVJDFHN/fCbcOZ/JaZrNdxGoplog7/SugDYiRg+/gdxyGgpz2lvSpSAmoU8p7Cqp/FsyL9kEA/hh
2cLqN0XJugpn2FgOQ3j6P4J8xqTZ/gWYFuZJPVRiV7YpGseTd9XcoOAp77+ERrskcazaKWwH3PNn
Qy349o3UTdPu4d8xD7j45puWqdUao6wJGtbU497I0pM0IDnWjChvNh/ko1QA5yt6coOGP1MdHDrN
/rvtwX3ImR91gP78JK8LUtdPgKljcQwn8eFkwslyd4vdaNKZfCS0iMQLEGgRp6JPY5JXET8a/o0d
caj8rzx9SM0oFdJYMBbQccRY7l5vU84zzDKZ5hvNr94JQ0o6isXVA9IxkZ1WlJEWMUKOeD+wJSuo
kBAG19YAhXStQm46r0V5PiBAXyRVlQ/HUHt9Q0uO2b3eKHw59Gpf7o/O9DGh3xeG/hiDjfxfDqGZ
HrweD+7DwXiwfka0FpofzCGccHhuZyiEGOIvzOOWqH0aWyq5QDrdDOe3wELSjyG8bVqyETVQ48Ow
4Wrq1SjY1Hsm6VYdkZUSrxMMenojDjhWsQMUnkUORYaGPID+r03Djtbom/0uvLpWwWD1/sXrrmwc
UccWO0BbPc/PklQ0imgp+Jc1G3+flO43fQ9cSDL3gPIO7fYG1ODBAJwh7rUlLGjXVOoQxjhrY1U/
KVUJUXKdislNXAf4qL6velPkq0lheixi/oOr3yo1tGKI96J0reC0VV+XI4upJlCuYRyan12PxF9H
wSd5NUWJGtEw4XX8SCzWTdBgMDvXWa7CJFwW1U2KeEsHmzSAVzZj8w5BT0qCFnXlzQe8VgQBIRxt
svlNyk+erjuhLnd2UUsljRwLVEYjxf2FKtpGR2Q2XGuVpovPn4boJzIh25w5vF7bIa7uXzij2vvQ
hRWCG20yPKFxQxLdKou07+Jc/GPaoDXNARzC05LJjXHC+vcEXD5Qz5fwCiGRwSbPmHnz84Qf/PFs
Tvl05CwVL65o+hrqcsPIqd3dQLeNhtHW36BOCtvUy1JTCOpbMHGxR3qz/LTmdYn3E39yrKGpnyiT
FLRL5j82q321HuQWjkTyRo4KuZzXFgDqq03QoFJEU4woCjiFXADi3u7CpBMSUNK03OFeUgKPfkRf
YrNuBQyvG4qdAZ1JUeBMkMgo8vbHyGU6oBJs4RLhuWg4K1RzxJAVbDJBg91zWSAtji+qaFB3j2/b
KqBL78fw380FHshCovvCEcQechYXZFwXxIqtJehi4yb+K4pLLuWf7tVZmRoEThAm4wepGTMJz7M4
FNvHy4rzODPbWCbkIMntcQ7EmWCG5WclfJ5K08FKNdOAd2AYjiyxavP/i/CraQ0tpzS1gptLktTr
paGPAc+lSzQo549BIqb7si3YqxsW74dtLbLdo6jSobt+P9HMu3Nonmon0tVDcvTSQFfFxEzJeGrc
6mH0TqYAyr+wDIlcv2YYQFA56q1xSfVbn/8pqaQCOQ85p/hrEHGuUMSBtUkLAenkMxxwDrYaA8wl
qlOnk9iyvt9cPMVsBz9EYzS/xpWO+thWYUimp+TTbYdw0R1ypI/IC7wO0BOl8jmyP+Bh1fEAjVPp
3b3cBp/H8DP10ZnmL28l3NbfhHA7gWZ0rHFqBgRa2sWPQQ0ou/yDrAaW1BUiM8mrHXVjO49VHl7w
c75SKauWabv3VS9iPUPdKZkZ5FU+JZ5VMKbSZfYCbLoD+v6VLZQDZ28izG1zHkoJxjGaybp34mdG
t8rAN4S2QKxpJ2G/e4JFXUI6/V16M7OnCHJgPtwnESlprLxRz6IuiIJy4F4Jy6F9GZ4O1IUW/8R3
5sh2wKwY7Yq46vZFBn5HXXeKHHiA98R6t3zX/hubECGnVIp54l5hIV6pZJOb7oG7VMyluMbA+n7/
1sf7mREYKBicGDkjepCK45gsSz3EhNhHnVUHlrmb9zJMb+gwB+IIcee2uHzkddTtLu9+6ZtlDP+u
YaaBL15S8g/Du2lSoJPlWHerjTWG8dPDiRI59yjVhl+ixe7i0y/laDk4ZADK+yYtZCBcTTGgiva1
5/V4rhCbS1vm4lXO6tMZnUq7JBIuHWnnJt7wfA6eV+BfyL1W9K8S7DeZFseBN8XdZiCdB4ZCjQ+m
kQr3ohhfXUMoLmPElpilebXn4rcWFu3TweiZCL0rNgArfML35bkEDyLfb/X9aTTOiwqCDky+wDjO
lanbXoVIej9FcJjzq08H03K+wKZpqEVsMtKVfeKCFsNgnk7whqKsnA4ikJvoXvzzmKkJ8cRPwpdu
uMHTUYLJLbFK/iDYUFFYxGorlke1SO8aeHxy7rEloqXZmSRYsw9vauL8LfL9LvZWsXAUBdinunlw
R2d/+GdQRxEIAgjLWMUW2kycAKFKChMHvMjaCp7DEqgrDI6Ej3j8t3NGMsDzFnmJoUkToX3v06UA
c8fMkNLs9Bx5p48gyxy5X78p1ENqvBEku8aBxU+agkDrfv2YfYd2brnPQbKSS/Hwva/Tx+eEH8Gy
PxgCAjt552BxodzNaotidW7DbKk69je5RRM3DuOJ4iDaGvYAhPnKwQZEZsKzLzpwq8WFQZCqChFe
6cneKsnmBrtj4d8m2BikJ8GhTovgfbRSGNCTAYGIFLUDxK8jNXsrqje/u3YU0t1+kfgA9LaYOmpH
cr3xHy3FRx1qzva/6t2B0CApGxxzplAcmoCoCadMhWITLIffUzGwcRLfmOTykLn9DH9AuhwLPbOr
Qa4IYL4geIUyQFXAqvbHPYzM9j3ncLEBSoml1yr2NYGxNOpoda1vZYigjGOayIxzei2hsp4hF1Xn
jdQwC/HGrhbsSMJkfH8Av78Gcivid/MvRX/M/prtSPh+g2+DELncjcKXygYnCJIMLvIfRD7AFJ0N
pPC9AX7Yr1hptGOSZTSY7mdTlx1nAZpNdx7LdoJIuiO+Xr64iEer/4rrBkdvWSrSuzY6eCRxow/q
NjgxHLwk5CpR+j0qXIbnEbqCPBGf8wy8BHPgxIQfTxm6OCpbjEnPj7qTYVDAXfh256GbjsdEGXBL
QDqASY8bimrWfApE6HcVaVQ/6ktiAaEIrU5Fb7NyN46nrH5NW2fs1RaHkVALOyM7vpedDEFIJA1r
GvIosndpSmlfuUcGP06iKCHB48LSsvldIm6msddLa+dZeXlxlTmR/UOSnzLd7FMsZw03217H/9cm
MXTf2USK4H61/j6BHPidBncf+ON832MNfvpGU/TdOYwz9DMdLjUjcYh+ItV/uwzj1P/p41T7V0Mv
l2RtkywHwhqgaz6IhtVh1Ey0mgptp2HcRI8GWIwBZutC4Pi+YI/+IClXFhDe8QbB7d+dJTrR2spC
TQP3QGVC84NXfPtIGYWkjoLCVHaiqv3+tl292ifEKsKu9VnRjnErB06uObBbwNOiy5ITHyAAlPIh
qvRI6T0DqFeqCxS9VAevsZsNy8v0ApzLN6nJwaGlRZ6/dsTllT/3QCMYlVnAX/sieghzpeQ70T4c
kqHG20ZkyN5nObK1vxrKcG7xC5qzoNPb7G4J1BWMnuDPbXylQGIDCbUSHPe9bbdNF0SfniABydy3
qTavR1RGzbU/VE03Yq3i82LPIVt6MIVbAXukWjGiTYQbiuKoSoKqaEeWTwBPYd/GZlW4R7MVFdU3
UT1KiGG3Pd6AMjJZTw1xlvsrP6cTsbjKv7h8mtTSSHk1xs0M21ZCiGuicVjV+MhOYwugFDZGHpCV
6FL9EpX3OmPeAl4/nsx6zcvToFF5HqGrWMv0gNe0Jw58MvxWIJxQU7m6a/aYO5UH1n757u84wu3D
jaf/UHZVbb7qqoIIKJiyKxncl1z3JUpkj6dEk0V+CiCQCXZJJ9YXo5qGUnoT7M7tMjaZErprLZJh
Ku6c1e2dmLI23efQ1/5CRbx74Wfo5ldztaTLlnc2lyfbtrIOIHS5IEqu25jOF+uh2w7C0Aflx3fz
5/Wvae09XpFvxEyshdkTfkHBDCMbtRNvGcN9B8eePqs6PDQErSvVpxCwhJ+DNfskD5+zgZAry+im
TFWGDYYeAAKVXejUijidnxddGbeOzasaUNQLWbTaMgX4VeSDf/Y+bjMrMOPGzXfL4XSdli1NOsb6
CyCDpm6gLRlakeGw8/azhCX4iWmsW/+/TYqc7/fn7L9c3RpVYD5Vr+rfbMnAtMb+vkihlKmNxbZU
eXQLKyS9oXKU3dJl9rAZdXkAJaLzve3NB3Aeb1caLCZPxm9ku3TfXkxH9QU4eVQrgwiSkP21QWNc
srl0+CvwWLaKWHFjTUhIFlBBWG53pUqREbuHHuxuPzkhHj+XCPBYVA9S+eemgX9XUsdfYVGtGsyR
KbWxMLEv/BBvXQEp/e35UWUfwg1asgf/s+IUOcctXyQc1Tdu30kj5L0M/zVCV2KZYqlrOxzPyzZZ
mUcfZq3oDn5s5tj1Pf1PPrQ5Q/Ux+owMXdo3PZFQTj62zO4gNRFthoYB9kVgDOsZF9pdCWXROI/3
eTdmCdTUXEVXd76anG9dLJxp6eC3/r3NgGWgYQkLm40lTbBTZ/5pRTwwMHJ1bpgHbUxeXyZDLtDT
bleI+YjR3pj9eRjsnDWraAz6nkJt2veqhpaQ8l3oXLxJuF7COdOOkDR0QTEidlUm8JPkA4hw8mQi
q+xPRpgd9fDs5xxfKeH392uA5gNtxkJf4vRZecQaNH5hhBM65ubJwkSIV1HYWzudo4YpAFOMN4cv
Q8pAbW7V0j5OK59HLrRjt/TT94iCvZQCCDCJebQS4T3j7eqoy07DhamjW9imhfZSsi23Ab/QOzV5
4IeDwTYfCLVciKFtCGUcQiWCqzBTIvNcywt4bzB8aS1L0DNMekCvFgPl+blQoCUx1WVdWQYjz94v
WPEjkrSERBj7U6UmWL9rlTtRPb0n2eA60TOoQ7dwKYpfcUBn+KxESl1vd7YBgecYqOScaaj5ZjwO
6HHanJTboac7Laqv+E/6hzwOI5jKVyVxUWdBPn2XNF0DsAbQLqk+AgplayXy1dAC4I+mhbhuYxl4
cH5NWlN1dSFr7El3To1WhiqPptot1sl4Q4X7hJ2ptSF2gPipfg4BgSwk2lyYhXxZVMRSQ5t7TLyv
agyswk84XXdvzCljfuxoudRXo3kSd2BSxjNSo0G9dJXCELxvVwWBROFHHb1kWx5DZBhLSZ2NBClP
utFT8/zkYE4EENV3jxYSojiqIAYEmREQQvED+HQ1eE6kLww4Mkjq+Ohdw2xlaE0FhyBCU9BcDk3k
BINj9+H22+YFtSnQeO9r3qGPUX3h5o02mrAiZO+EAIJRGIEDxHpkcdI0mddpUdDkNGw8qN3xrTJm
E2nWv97leF0+CkcYH45FzyFs7QR/MSodyGKu164GbHhjDoT1BQEI0TlGLJpTcvggrBaMXeo6v4iR
g9vqDL5lErGpDvvg7C4RPCigXxgzRL1tNq7Sjy3wxYAmlB5J1M5K3/4MGhm+uqUzUGkOT0FfD8Tc
JVOqXSnj8OVkTRgMgqRG/Y4RDKBpdlnL8xDqjc/DO6I3Q9gKIRvdSDZxHQKZVfF/T+W0qa6PPnrt
XKLra+Y65q5SPZGjhg4x3h01yTflnvGPManWjuuNtQ4JEF8Wweu5GQ9Hq3uEDVUf6iXsta4LxQFZ
a304+DAKa75QL9gLAYxoaZbVOwucB+TMF0OJe4O9PLLpl7WyQOL1t4vQrv4P5FXEwRuCGjGf6oEJ
7dt/+JSoAH1OR+FIk61bZUWa5t7x9GI9JY2pOcCIOyRAMFv7ftPG5/jp/igTx1SUCYgNl8lKFWtY
P+HLWXPAbVfhX79V/CXhuuPGYhYS3wmDtlWbgOhnCYZJzAJewJLqufbka6B3eW5P8sZO6kMkvfMu
4U3kq11PJtWbFb1SLov/3snyhKj8sMB0Zxc3njwZnMRv1gvFK7G69INi6FUsSMOfcZtsSM6B6/wS
vYYQqqM1f1bjhgv2AQ0xg6BS7ZlujJutzCWaHdqQdovUotXs6O0K9/nAZ9lUc2L7nvQJQPIwparl
ymHMRgSm+uNnm2QrSX004hsXBJkHNeRyW5HXNu821heDwo+NGCW+HHZ7msJcTR95sfz7CQy2JpGb
6hT+mOOY1FgPHMjLnJrr107/DfnNxuGOOgDULn1Z8XCdGgrc4QTOgVtBkBIQ3hKeb2xpphrqXTbn
lpke8eZbLzI1WYxi/Eis9Ozn78bEWVgUrTTKtnzidHr6CSXCJcYGpc5EYNSe9FHs8cU9Xm2jvZ9l
CA7o7HpiwDkH8POXndk8AhZT8337/k3ovqkMg4dKyqY3ZoNmVR2T/9bVBhNekyTcv+N6B5KaU+SO
qTyxn8g34xkt5XeS2H+MTI5QPfl1/3UI1IVwK0DCrH8aUzqrVfBRDBZmE4Lnlna+YPa/rlT9lhP9
KtKm9GhQ8IJBBM/KBfqepGKjKkQkhqPA5zTOxF3hAFV4Tch+pKpRCgfmBt8D9DWCJeCAdftN7P9O
Fqqft+59/ek7DEcj11ll80TQp/scwVMbSKYI2W17uXoQhTEny7dNGRS8hio4/M6c4JdWv98UTm2c
9mksjuVpO1eczp5CipFMvGKOz7amtKqHC8/vufM3+V182kFGhNZhYJfQ+6US+zDwkaGaa3KT8Tqf
qn0AB1G1zTsF3GO2WrTUTZrwQyTmen4hf0Be5rP1pNwFIElo8bNBjDDPx6MXgnYvct/t0ANvH/aK
ywpQs0butpa5z0dLxJMzRDvbxn1kb+DIJmU/P+cQWe+SlFyLB/soTYqjjA/iDU2TxEV5JuzMvdJY
FESm77WoJ0z+cXDfwCPMFTAHIXNksA8X7T/hx5X8PpTs7sEHV5/zAEiWD4dXoUal4I+HdVjRGAj6
EYUPBb8/75Gn1KWmCPtCou0FNYt1cTXPL9FIP0hRXBOCuycqj1qiboMzcVrsbH51wIuoc2Bkp5Os
07Ojh6EO2JU4zJjSIF5JX2gyMjHO1X318S2yubn23bQI5djhHnIoh3myBXSsKxga4xn3q7Mzg3Vq
JrXqD+E6snAGaUjhugRs9+EtiCBHNYp3ENV6W1EBqhHGpu25ALtW1F1cX6NWgVGCDExfodCFSkZC
+CPqdabXwkCJQ9diBvq+SLLYk0ssenObO+NokpLx1lKoIlePYFMxZxRJhvBd6KvAlgIQjBGQPZCy
VXr9U1fFBCRJKv1ZB5vjlddDD2LbzNytsgLKKfF3J/QpVyMgza0Z79dZjjCOWUeK8+vjZAGaNjSB
wsNi1uHmwT2TzvRt+JtY4J+XrWFpv3/Q7vHtb03+9815eZjIHFq7n4HfhQ9mvJjkEtYH26JiYe6E
ABy7xv8QrFJGee6MSKETZDFJUcZ19EM/TSJB32iO3OTx6PFQXpiuKSb57I+1REZQqUksUGiz7UZu
MCXBMg8KuzEZgBH9k5znjehK4/vvfqvirMYnFWi/LCvTd4+GSDbWr41BB2MoJHewbseoQXCAAOo7
biK6sSGwmQzClKA2ePb2f3s/xli4sg+stRF6nMUBfJXXJ/DKdNyE+GBZXL29LzwtwfVQ3bDAyhzO
ugZPznKN+v7i+LmAyhEkX/+jWodkCVkE6V7F1XJGtaz5HjTlw5qWv9LONR6/+vloGprdyQPm4vXi
orhIGRX1wJn8yDJFjxKUDjsYkQITf+1QwsHGBfUuLD0mPFiwYrS2b/hL5rYkw9QAwI/N1ZTCWjz2
oTUoBRKk1tBRDajjq0o64z8x2JOOxGvVgHu6XNRENUB+rhDL3x8ysvGHIcxPQKz8+/VyqFpM/nRn
W1VR5mlkwho6x5hZ4DDXvZyd1GUMW0YO6ycdQ84c1Uo4ttB0Ig7JtnusrM+HPj8E9zRlHSJyke7E
g57w0gIqZISrWM1tP5WPEH06rovZJNLpiGoorj07FEoo2utcuUN6/ytj9lTl98a3FaAWuKORWjmI
YnyBAXjgdJV9k5scdRy3o1h9hd1Gp7K2qLVlZCjvpA+DO6x0CJhdhxY+nNdMR62hhLAh3kMN4D50
bjmvP7nz8Zwn+p8rnyJ/bydNN8RhXkDaeCXEMo2GLg2bDVgxs7tiYqO+fFoXwyvHnmfMtZHFl77y
d+W5LwLCM+K8IdQTW39/sMCgDm44jP3bcUWbQ67ih4BV8oggsxnL8CfJaurpYjqB71frXA3rKnFl
22nfJzxgXwbLDr+sOqaMrb3FWXZLUFZKbM1XMoTW2ba9hqewCG2Oo3j3tw4DLjVsLOBsNASWjPvw
PTPDTra0dRiqf6ciAmU1vIXZnQ+d/dMwq4N/UiYcbAjx4+J/y7S+RqXHU4tbrzweOV3b6LUz2/Sv
7KviJWNmtkVLIp1bQj/SWOfyU7lIaDIJqbWTAFgveRr426WhmvT7Vk+X0m8fwn+3JlHe5Ugkx9BU
K4KBQDJwfmXgzQGi1mDMS8KmezJM7QNPEEvNbfV+QlQS8tp/TM9Ycsi4BVD8Zh0YEZshqst9AJcF
5P4rRZ93HYqhMQQNUnnDT2Q7F8qMgLrWFgmJ5VGDLsBX5czpdNNknLIVPq/odLMnOt7pC2PF1f4j
kfBIMnUBsUjc6Prt0+CCA+kQE+YQHsHFx7mm5xI2ZysksOuLGXQJeTfiKXjz5n2+c9iyy2Ofy6hw
9jmmchs/smOylEWOCXExTyUOodInz+gkAgxbPXva9zVBwgTOkTro6Ub1qtcOPXsly7CNe3BIFOy6
S8nuskR616d/ios0mQGAHVwWVMctN3zE1fStgcqQ+5x9/GHsrs3dsz20Ave7d2RJHZ3jF31kBHCy
FYbjt1v/lzCfuYzuvJujyhUMO3AiGcOlmyy5id+JwdMGdMI4q1gJzCDGOCGCUYr2k7I37g62KAb8
4XRGBfhFLsUIMpJ9kmRc4hEMsXp2VZUBhAEp8iaHnPdPRZZzjXE9HyAdu1uDbAoCz48HDg/+JtFN
GFzn/hyqGuws0am3ngaeNVGDsvcFFoDzcUulHjYK5yTxLyantuy/kmZXO9TPMxjlV6vahi/qDXj6
ET83ak/BzS65HPqr+27fmUew5GHTrjY23L7WpFm9fn0S4r6/ptxlb1cgyMR0YTBC6VSRDGtAtQn4
8EAHJ1Sr9lClFp6Bx4E0X2FXKfcY/ywKkpDo/6HOu+99/3fKSIOmmF2quZy1Kit6FGKv9+4VfpQG
iESj7xt93iuSBleg1dA7QsGlxw6rXIsQKPtPPaHXrrjyB72zvdV/TFfbBme5P+jnd0/4WrwCgeV7
PEVhmi8u5FgfkRPcthMCmiY5qylajQQQ+SEIpqOfhnMDeE4R1PnKJdpRL8HlUpYzCergNol3s5di
B2w+3KL8X0dDtwTUCDtH+wll3dnABVPZRKEJvc0fjGr8ClfwK7/zdDg8YhoCRMiS+JZTctXjwbB9
pB3fcZE7vPUPuiWOUuJBjV8GZQKA9nKThy3nh9dS5KrmSjvHxDTPyAGix0sd5ZXGaVTO/qoqEQFN
A/Chi2+4x9/2PyR1preaPzT1LSqgv2FZxkEJhhm3vFlUNNrFCHUMqBBKUBUbIaPt3XeNkFgxBTGf
/UHr1+3OuJRMWIUyulLSkZUhhAysTsbuRkwRcVKCId9rDKaGLKwk4jm7dNUV79pb4fIvbbGQuM0J
aBpa7GJ7Kp1SouMLuzdjNNivdsT3hGWRKv9tOB2a7Rq2VBz4OyU6qoLL/IqxZ7LBXh3rhetTlUxn
1S0fgooD85ddfhDD040HVrsCpP9T6naGJUQh4JIg87aerWPiG02dOBdd2D0Y+G/XxY11MGyGr2ar
2ZRAp37dRssLU2dMcBdj7xjuwvzbWhnDY63lWg7wosQoN+QCRTJNE5f5F8rRXPnRHOg8FGd1Q13w
9QJrEG6hotaYBw+HDCjqHE+jjYS5m5IFCVDYY7S4o6ktHzOwa05VNHNHR2QSeCWTK1wALMVRRRUF
kkgZs18iF3lgiW9Fu9drZCbsSKpugrBpd5Qlz0J17UIpLUXIwo5u3eCHyH0Zfk1pGSb22eVasOuf
hLwswoisYNEq3zqJWT3Hn2qSBS+lu/2LWvzQpK/a2sEWx3fPVeSThuU1K0BWy12LTs77T0WYWoFI
4EsdsHlyq6oghh6YA8R1MQJBU07l9L6vWlnSR6ibQWP6zwS3QlJQS3+C0sva+kLNLr8MMoH2etDi
CAULj4KnuAhaqZHcK2XpFN+ryVA8zzlCvt6Bx/8f3y9VMEg3SdQyVQD9rpFz7HVQ/rueWMO2MvcI
HRLromJCRG/uI+pwFWanhuOb/2rvVfff7VvageyyIdXaL6xKowetBkKnkU+dOpgLpHpNjorMXIAQ
Mr6gYUYmv6u2lRYzt/OwJYpy8GM/Aj5QK/usHNNO+l1inV+Tl5p9SDwaryIUrrdhJ2bLGzK020Vc
HDHQaMUgWjzOPXsOOIkJsOzAi649GSrVoUUZceHxg/BD1Av/ljkI7ZxZRTQv/usy7dwtipcDqFVK
r1KYHqZ33hSkwfJ9xGdDwKS+a0biI2NhxvqyMOtUDVUUqyuoXHfDwfP0at6Vo02yqxJ5dM3A9X2I
zBK1a2mKWkKz2RX1cAZpJOkmy6iSTVkLwL5sbVzZzqDQrFnO+TcyrJqf/00KN0QpuIC4WzDjlZWk
0L4bHeeoPRQG6Kuppdvgf4avGS5yBXDvVHy1q7L/VF4UzcB2pwA1LdAAKFR/J6ljf1dY0Q1Tlhje
97g7AWMD2PTnTbPptZR8lYe6tdZLQzdPZwQ/uBQMFtxb68bOsUq/LQqPYziHdIre2g0J7XYhn4fJ
pfHba7Ka3sJwJASERwKaqG9dRHKoCCo7x2K/XYfpT2BS8murSiW1LUJfjJ3V34Bmmcj/MxPh5bC+
6R8J5zU/Tt47CWYCse7Ih4hkPqYFf1DfjSff+Eju+ENgoaoAZR9FEJdsqG6xjea1V9rLTVTY5Ddi
NWj9vcYNAFrYvC740JUahbj3/Fp+rzhFlmRrTXBxfiCtBPJqT84G0eCcDQZ4+fXuKsIbltdU/V3x
jPtB9zrN2QqGAXWBq/6+zYUmZMWofS7UNLr0pIjiUI5l30qonMITNSDinn6QthJP4XN/LSea4LzQ
Gx7ktFE+qszezOqZ8fCcPyIvZhgrHJz05bJY3pY1ySXUmI5Sa/A4wRpK+WTRKFfXymchJXxq2T+1
JQxosQwPDQKeY/Owx+XMvWd57n0bhU46l3SiNdVkuzKpTzZhAsMmnlEzcT9j7lNdl+B9+SHr5H/Q
73gc3Lpqcl5oRXqhWSASOMeK5sxumRnRmxx0YPPn13F96LOz/P/AupqFMLqohiJdthnOxy/47MqC
+VqF4EJL5Lctjl1tNnuFj5bdnIUfAncYfftMW2Ld1iRO6uDZ/F7sHm6glE8pRd6NQrC3LMKxDqRU
wmU0tI+t+6ZVsJidosnkKO7/0ukC/uKxod41pAlS+HZDUM94gSunvfi7y3uhU6QueV5/m+3Fpe6Z
S6ra6yljIu8wwVOmiAbuF2lepZ2lI9SR9cDXeZz32POGLDGAJ9viGTNLz1BbFkJkyYhpTNpA8FY4
/CI97Cd++TgRdy0JTrIdhip93whQFyw7JNZgBBZYBP1LfDIAAWiGNawush66kZKX0vPW+2xnno88
2XBr6GhrSaxnxSwZNG9bMae+ZhbOvU031sK47nFdzqDtfHVEXxUC77GcyvpUM/7T/i1xquqpTclX
bXTtfn6uvWGTm/hpIg1hEBImI+3RwucnNSOO1fiqHedKGzOrPLn+QU4HR83HAsVlJzrURxvJraFA
WF8KsaNO+82i9VOBmHnz8M3etHQ0/9KlivDyyS2vEdODRsSx3v28alAd89zs7NMHSiqRXS0PeBLc
p0NoceZ9WgGFGClaPxX1kxm33J4RdA5+HfdtrFPGzl9PiAvCNhOa/PXBEJrLwI8rHquBcHu5tAQi
o/jPEOSMFRoGWGMzxwk0VrEVij9XSZgSVGHMLQxsZCeVHhZ6QMVk/f+rUqO086oLCr/WZUhd5cud
bCfKVF/JN0LtKQaCgT3Km/mTxKhtXu2Rutf7OszxwjxmAt5h8iFCgt8YXP/Fbc1/4wYB6QFrSY+T
WoYzG3A5L1Mvrn8eB0RPDX41iCGI6saIYfw389ihUmE0NwC67GJbmDDiq+y+5ZArNph7tECqMco8
xBzMZ/ykaW2FMCC7xMKRLaa7dhKCPZcedHKbOjxLkRHtrGPqi8CRv4QSaLtdan09EpnX2GObvdyy
o6FFYPvfxP8ReCn85j1XuPFQqHAIiZfc8tkpa3R9500V4Z7cL+It9bL3eEQUJPudQEWz5k9rj++r
Iup6n+q1gtmaTn4qMOdpWuOdkQ56h3yrhBdUox6RUVUUgKCy1YIvVuw7Kv6iDatpGSeULTzp1b7O
70fGsnQpc3XWZNkGm+BPGToNQH8JZS1pN4FoRyZ4gfPEJ9+Mhz3IVrlZ7kQtnjzT077hAuoeonml
uGlE0gRxbTABVsYmO9hdrGoQYu5D2w7SVOeJCz6vAQIyKhlHjgsExB43RWVLdzCspuc1n7D1hesa
dCrRKLrCfSaKIRh/R5i+Xf3K/oBVsqd7KLU45EBR8cwtrQpna7ino4awZqXcyo475G3+Vi3Kl82m
9r2rUYFbPsR+e8ggACQa7KM3mUpJc10uid4hC9B5ET3X+Loxemx6OknG5Pr1tvc39rddsLH8+kz5
EiAx3JYqrJmG+Jm8Twjk/ifSazLURTiYLoUdwVRelVUtkd91/1N3QgwMM8vMy9kHpVvb45le9qLT
zADvkS9sl7SxT4o4gmOKiLkQHYNaBA5jxlCDTgXfmXME7lMmjSj07KJZynZ/nq8XLAzU+BpVP4Lz
dmPLnJMi1nlzqxYY+i5djUes8mElF8fuDo+vB2Tr3020pcEstYDGMTec2u0VD0mkfSrjbLiDq+E5
6eQuvpbzk/343rd0nJdeIiUlKUenZlXCRccM4uqt3ceUPPrMo7dNtJwI3f7vMDjmW3WRGnCMKxh3
fnIDOVuIk6VxbgTAZSxHH4Ye6il6MsLLGqXZX+RILp23KNl+UkrCZ8WyYB+mByi8nfAqvYrj0TWB
eNe22cckE3e+IuAaFF3yCV6XeWkRvuDMxN0a3n7NJjv5Tou41ynrFXIKpxj2+5ZxYmO83OJUOdam
pTwn4+2Pc+MRr7KOOAMsCfFG+VsKRaDxi2JTvAJO8RswtHSznlTb933rcr/itlqJu95YNrBYhlnG
PBU9Mq0E+AujjLeWHGVcdqJYhhjNxUBnriGizFNFTHG70ESRPcnl4wbhLH0NPArk5fQkz039rB9S
TOuVTeH537Sn66UiWT65PzcCkSGgL4mHuObwGVhRVFYzO8S/YxZNyTcqS+lewp/Nhrx0AYzk4Ywy
TNspJKWDts4MHEsvopNXmMAm5t1VDCnFrSITQz8ZsDa8cW1h8jFu4DZLrT+Ia61gePX49P0Whjpu
dureVmUWQN6vjkgDIhY9d+4LkbB4THFSE8MUn564kLfHHlkoD6L08UBLu55rfW6Sg/U/rDP/4MX2
n7CN035+dN2H93+jzhC7HlvJcx8AsNCaDCCKYxdtqL3V9KSLFR3vnTDSFmbp/IFx35U4ZahWX5zJ
drAfycZZLswCVQT5dYDANEcwTDbn29MmxGXPLAFqgkaFz/6Ku8fei9+L7ihg2faHkQ11ruXmNoIj
fkmNubTwi1rzY3HZaUJ2MIrB9dIO/CjEMAVnTajVUSPFi5THdg0Tj6cCVVNklkjrl4KQ3cy3E+ta
MrGwqfAZhh73MQ8BmHHu45xSa41yYoYfE3iUBMbSTCL6b0ba2/hXIhAEGsRWyJ3s/aYfaUQ2bwS7
ZBpl5urWizeQC7FjAc1F+Db3zx0MJU3R4OmdBkoWf39KRGeP6r3C06Lc8vwIdNLPn1SdzTQf3GNl
uYx+ng1ai5kl5O5A5Cf1vhbqMUyngCSTQYo6nT/oAHfLMB3Me5kTYJQYCmH9fUqiOaG3a9Jsyc8Q
E3yOSOZwdAo3KV0m/+Alg3FxG6vMij+l0p9O10J7w7hhXoV9Cg4egLuj/7xNBd//HwKuaEAisLjf
kF23MII4WJIaDmZuXjlaW7pNsOwEK5ChKT26Wkhf5Q686L001L3owuimnSOX5iryo7UZtiaIO1Kh
+TXRsPl8gMCphYVe0bx9MLnJDDbrxLlK470FMYq4ziqg2gbCp99VAWURMJYZcU0JGPkY5C1Xdwra
dU9fzgsthc/J3RJFt3A/gDU9xezdC2PdGyhfZhTjLHJq4r9mMZQorIQns1j0GVDlMh043VybAUMb
qfIJP/6abzlEF/niS8VH9n9fjUFtwkIlNDNEHZz8XbTr6UMfYIy39NHzTjUwiSxvZQCtVZ91aBae
VyzYPhwCN83Urfxd+vWQDNypLjLOtwKNW9tGMXY7Yd2QAUVw2vwxnFecxDa/ZjNiNV4p6yjYihzu
xTjS+qztTFDjzCW8EGulhozWZfHXfuAmqlnl1V+ZXbozGyrXOJzn/N68SB/LvT0MLHtzQXwscV8Y
YWdo5wpmkHc8UEGx+B3NDajW9TWKjTKC4RuVglYDzxygAWGd7aDYt8lzFlHPFeHJOdLkQOqz9cig
+6BNtL5S7WQTVFmFmBBfXec/ZMicTuNWqKW8dY8ZvLgrzIxxN7hFTS5mAkEmQyTQzVkNXL2NSm2r
9t8E8H41N7Mj175KHz3Ps4pXE0K0qFoCLsBtiOfscWpuMCoSllVCmyUVvHzxfwHtmoaL1jrWFqmR
IvJUtHGPvCcOZ9M6bnkQLnLg5L1mUNz/nZMMFiLkCbJcicxjBxtx4xFSCu44nHRt8qAU7Fo4hmaZ
VigzwTsyRpnJqb6mu6nQYZZg0Km4+pGsWjD6ybSYmyE17vOfiq5SaNfE+fCQDGGGL9DimaTCAX7Y
Gjw1Geq+fmvRDqiPiDB7Tw2BQAmk7lXdcyjpadzYpWl4KT/7XAtrpN3cEofvgcFjZqreCo2uVg/b
Qvq9yTjR0hZQZNDrm7rnciOfXLPOFrQWxEqGhRcCjTWjGR7vNuKrfmjJQs9hEeDIDZloGkSUdGXK
Z7BGQ09XaAy5QRqX08lnkPkTtroG2pZ6dAnzZw2R9/WfKjO3kOsQitZgMyoulntkAMZ/j0TPiqCs
KsZsLOR35JJAkMO7LsL0nDMruyd2vpOAd4GgQn4G8VPd87wd72lxdxNn5WYepU7b/LcMWvP5lHRQ
wN7JcW2xYHbf8IARo6DzN27xUzAvahsaDZqAdaizlBbK5Kb0xThckb6Zj9aR5SrPvg3v/82xe2Qh
Wk5Rhl8HTHwV+Q+FNXpqkEJ3BzS4sDhdUzYNXkqCMEzTYqRV5T4lpeMR1ZLdnLKY5QzFEr3MVJIt
m/Tmt6xtR8ndAGE/HGuNUha65kZft+JWfABEWk3tgJkZA6LMfwXIHW5zAaWgUqKTarx51MTwbzqA
NvP/Us/qPJIgHIogX/FXImED5BPzaKSZ0j5TSYgDXB3HBKrmZ+y0gAP9D4m/Tn+h65dhOgjoqd3i
N78fGIr93o+cTNY8dRoi703fXFQZw94gJIDj8r8iO4mxEaPDT8TJoWhhkGobVBQmCzd4ivDnwg/e
TSt7F+MDk+5ST96D9a9QuBo6FrYi8Zgv5SVmg+VpHR3W9zVp6btS/WitoyiJBzCFmJtStjji7awB
UVmE4pTt1HfmiFlQWYlctqcRQvM6CjYkA93udFsTqbY1H1xp6QUZWhEykqRmP3W5k7UCGGVozPEB
LmElf5B0JvwjWlfMrW7xNToCx2V8EYVz01/16o9kPuOHYDM1TY6LusFqPYJKfuFpwKprAq0oozEA
Cq3wDLHWoIAzbq11tcgcEk0mae7joUm+KROOw/0VDSgdfu+1Ixym3HMOgzbX928Uo6TsFKHixxrv
sbpC/33qL3ZKRkoZ6DnXIjN6F7j+1VhMKyjNfzGilTI+G8NxW4thC62wYRv7J1jEVoyjT7eqsS8q
VT/ijVDciC2ZjSYYTUi2tHMds1ZjiRoE1/PwEBsZjFMVBgHWw+iy8evwplcVYURSM0Xu3IXF1fFY
alYH7mQ4wnb5yCEdYezPsfbkgenkf7mAW96dNEtpBXJ4IcwAq2Lct3298rACKpb2ClSqlFTHMUOk
4JeT+tdWP7eN3IPe0QgGJeVe5ihrYUBy3v9jkocK3H5M1jIfBHd1DtmqZq3ufB8rMkf5iQaAdVPt
NQAUlv/U6K+kwOctGXFQdn/Ad6t3IzoSJOHgCw9pQSByfWN1HVH3FMoyAOfgRTDKcFEAoinecR9X
gzyL/Bps5C5v+GY5msz/6YL/DTdJftcyVKDimgRbrNyfw0znuT5uTSwexn+6bB4Qkfp1w746bVA5
EV6Be9Uo7+pL4jEjV9G/IFOg5tRRYkgQn91HFOjmpRkuFBwCtRM3TcoJLxP5U3CvKNOHZoWJ5G6p
mTIwNqe1PUbzkvUDyJD7c20q6XAH1oxmGVAk1EnpRXeG27SkOYpO+ll8yNzX7ZHyW2B2sPHiHs1o
1zqDJl6uXLkWauNk3k7qVkI6HJdHunY61trlZ/T6er/BPiA1CILczeXCOo4TMQ9VCBPAiXYDX0m/
7M1JwWL9BqiHchZg2vWeYKtcM8qXT8emaX2F7cR5k6gdKDQkN2of8QqYxzfKG3z+qwp5XJn6insU
/K1XisMcyFblol+oZUpEzEtw3qAwV3n7pjJXUNMe+YJyK8iplz9AdZrV55WTmqEk8yehlw7rvxzS
cTRg/scU9TtvUt+lb1f1p/F2jmvjo1RHasqFlQx/H0gtGT6t6mbuKBHfcbl5ZsGCqlwmdJWwQLul
AhfuwGoxqacotItEj8LjyVZMMkCRmdqsLtBenheYfW0vm6qi/4tjT4SJhVlieW6YO5WrEy9W1NDe
bXa8+KvHUB2yh8UchlTcOqzpGOx1SYvpdZIXjKQyyGyZ32A768mI+6GJT19qBQy/3mbZWMbsXmDo
vpUHS1joSwEaHIIeqzuvrlh0T9NFiVM1z5Hahcz7b5/i+c/FGNvnvWqN/gxVNEfj1tMxH7tnaIYX
oPv44A8aa0OUj09x0LKvFqH2m3waBvyk3DgjmrRoqhbKWo6bP5YZ/EMQap0d2e0M4TA7bixWRa2v
h5HNft0/dqK8ck/t9DXiSgbQN7g6oyyM/adLreZQ3BuiT4IuV6qxeVcp3x9s2B1D86totL3c2h1v
Nh2HEcbyckxITenRxjDDYn4Z1r7KKF1TZRHCyGkfBHLJN0FLqE+PbdTlNUbZ7Ra+KGlG4yeeVyi8
sa2glP2vskF4zGfh87LJJqkm0v3X860trZgwPWuKSZIlzlXSLdU3J81uw6ne6b6lFEptbMwz5yKg
2degt9xHXqCpz7LqmzQh2fX/dV4AwqeTPd23YXSAH+i9ECOmwzszsKn7UtEHL4m6t6sKAGGOjdIJ
nOae35L63p8W/F7eKaws47Bzlc+6CZXZGwrg4sPLsOx2tO3o2+ySYupA5bLwCQlu9gNqTieH8Ojk
AcycjyDHp5ceC9pSHc6DS8zr0/Xb4AVIVVFVeOiaAuvZEX453pCYrL9KzEmdKb2C0mHInw3StXoT
od/m+gbb1Akk2EEjT2keQ/UM9/PMaylHi+9H0cD8pI9xUue8DH0d3PRem2/qOjraIFEJoY8KrC/R
4C31lGOTwO/F8mCcjVy9mk0TttFhINfr2wIcPsTMzVVq0iAzfxxT2qs2ATkCWA0QW2bJu0q7YwNm
GV4CjoGujKN6QSDkc1tbkjAyRwNU3rUTMU1jZJtogRyhURB92fWARtcblkTTsrKLXIH6V0/wQ8T8
JohHjESkmHizsZ4C44ybqmudwQUIFr3A8tqyH0/iBd5lJyB2dnYzy/2GyCLf4Il/oMKJzPw3wpzo
v2Ws7QxHNUL7V2XWxJK0Dr57McKmPSpxnQIYlbE05KIKa1OWdNlTuVb8R5vFv8L+h2PzL7RKqyup
+UAYDf2BwCTTnHTMSPAZNZeigTCWnZHBkc9vLnIqf0GDPbbIxTcB/4BcJdQ5LGR18R8VUBe+EwcH
AugBIrDkR42d4DSguHiKGdG8uDXgR/gnuPus+DwFitr/x58A7kqeCTIH3GUvu+Bla/lqWv5QYboI
DQx1KGKhxjIn/wF9BkGFWhrCaA6fQFmJvliw9ywnc4vbOxoHl0qX65hPqAjGMj1s+ko1R6QvQzJl
71jyjNWJnogjhTAdnMkK616tLOkPNz7RLjlHUHdOr1n5Cg7coyqqkh+TFtLp0GtcA76V7+95qcFZ
G5OzMg+W9dF+lIUPoYB1PqErJY2tOCp3NODBIvz5r8hmo367uXqwHevPFZdV1MbywqAB53lIpm79
MrXCXPSsVVFYMF6qh6V7NisFU+fkOFt4mapiqEPizjXPkEPhQgQkcQQ+vSRIuKKIY0601h/46N+X
0Dy41S8nf8ktjMtjZutdE97/12f4m1UCmCAYMcXFQas0LaLuU6+GAplBKwufw+S6AuQ4S6uskZgv
GTg+owgfK+NCduhaEvdgQCrZX8ZbdNH9WvUlUK8wlrb8C1Y3/JDi44U9GeqxKQ6YYk/49QnSFkba
Bn00WwqKpIYW2JrfhAqgrXdfKoPdMBUEzUEs1RgnSH0Ep7zbQem0VSfEWRFrm+dOM9IcAHU0k0tQ
yyItU8n6IIkOKsDkiGy6J7wOGOtiCLcD7CJjlUsxO2yIYg5wVI+akxgTZyxxZyysGIz7F8yXOYXr
8c6phhrc/fURaD+GME0uvfbk/pCfwEYDHcGa2k9WP2f/dIveO1xxybtK6wCFwnyMisp9ZSSdgHyF
YCE1CBxsIJPcmI2+I1XDwV2oYuewma4V3fDPq03iSNf98lmk8e2GW6reHrE1e9hPE7mTxsMad9ch
q3AndaVXb8Jw2vLEIeS6rzPCPenFcN29u1cxBGaGPC9+db7ecvfB3xhXWn0/V4Of3boTmAj5ps5e
WzXKNEHpNWEdrG3bzmzxrM534utWy2YiI9oj/SfrZzPHZKVpJTVr7xbPdZEvk9PkG7jYk9ewnHZ1
PGb+XGgsovW7UsZVyLE85j1F+fuozXKPGSQWP6gPEIEiXecnZ/thfsXKBNtnzycBxYBanjg6i+NA
cAWpBLpW0rKX31pZluVyuua6ZHvJjWrvMJ7tP/0i/YXcFaiKO45F+3ITHZAsAM9vsQjkOp3jxuGJ
IeHKnK8K74Tp3l8nC8tIjl1ZGA5jwWqhTD+3/g5jwU8q9v2h28eLjH6KC5N4UN6xZ8dWk4S0C2ah
ej0X16oYIgiLK2KSmEbLthb+DyB8AKee5FeBc3rISP82cIg06/N70PJW4rFnrnn6xSj98/qQGKQz
USE8eohtb/vdRMeulP4AHICgmYh3Nd2lfXMKatN+YJ0snXk6Au73YTRfSoypl2902O2ybIehs4xr
uflowu/qz6Geq8Qq+1oaTSj9wC3kJImpa6+/O7bNHLxN1oN+gPgdz14pQQ8Wa3E8fYa/o4rnaUgz
Y6CsqmoojOxxy7wtLiXMwWNsREKm9F7fv+tXkqy6563gLqoqdkVrD75m160rUuB2hwDvoACRyVY/
jVNMuRDDkqg9/mH1o5zgsJ3KEktp+vCovlvJRzZHuNnSjYdk8zE9AZTNeVazhgv93mQgcyA0Sq0M
KHZRjpze481wa7Eo0Rz1qld17Rckgf9S4+WoyTxWo1/9sPa5LstK9WaMlfWGrdT9YeLtTTOSlxy3
63u9dFBlxa4w9QFeENx0h2mtgF9wY3udfZw+9XSPF0KxTvB43IGKMsPPxYrFn8uGHBVg8TjGtciw
Kp6P7aYANsbt7/j4BcfkKGGA+7Hp4BRrcjJsI5koVMeG/kj6qg95uVCeMhscQnMmsJfWtTC5MwqW
3jnEp9NlbS2aUbkWQjl+q9kVYwAk1EUj+nwCOiT5geg1Q/PJNbzblH5jnhzdMcZzS4eLOLEyJnIW
g0dduGNyU6Qnuu2FTmGStpPZ3kJ+inWwxL+p6tADy74FJFsHbT4qdkiEkyeQV9BwA7uNuvPX8ufT
pHSniWbACP9An1qFqt65aFTHAzQ/k8Vo/88Yj6qAC7xkGPYorL7JdWbcBm7eHRnY+eINB123QUND
0v78NN4olXF9HgtDbbeNeqL+nKHPkioPSyBTy/2VS+2HUDnY10s+NNqXfGiXWW8csrF+aa/5nEAl
+CuEuBBW/pnBBhcdnUCHeuyBij++Sd8M5YBtHq7d38U+pUaqnHfp1RWHESejiNrRh8BW5LiXbE1G
loNmnwgTIkA6IOBWE+JQL8QPnzJp0xh54khjbYNLAcPSUmjU6TPWmFkv4dti4VW79x/0huBYRdaG
i8VcSEhH6tAKpPp/D7fJaYp9+c3hDW10N01vt3K5D/y1xztFyHyN1Qb27O9KRSyuoFEGO2UinU4j
O56h2HaTARgXib5eKYOJZWul3xM6hJ7smxSZUPJp5L8k407tpnSS07rCBsFuY3UCswgVQX6FIzZO
r1jBrsQn22aOpw5jRw6rJ7odJl0YfYveywBL4fa86GS46VGXarbhMqua5u9DB1+m+3UzWLUkUfcA
VSgpB0LEYBQLq+2m8V47gVHcLjQYdYVFnNzQNS5CW2N1NtnqDSnAIr0i6++vbEdfaVKucW+LSX2s
Bw5zEDrfrDw+lCb2horTnp5Tzf7HKNIRxS4bfhN71R6gzDs74lT281czyz3J5mmJ5thKNkTUFZ36
r3u+ogzDDSCKpDfuRYGTWkGc4OFKEnndtq/YQJPKkyhmJtJMfBt0p7+ckMIKKapRbRXr2ErG+9Qt
1Nz1X4YuWXyto/vr5QUWkX2V5XbZy8z8OC5d1jt+BX0bYhwN4eFHpXtoUPZzr330ubu/sqQEO/s8
vQyPLEmODm4zQQYgu8btJn2H0/XP0jX1jDFeSVqnbHeKYPnVQPHtZDDwMkOFgfLuXbDLhuXqZ5UU
ayK0FvTn7Nf9dNaBVkOAok429cgDUEvcGwMeUb87MbPfXBqe5G9dT6nIHqkc63Xel4aL1Y0dWBD5
1QAQ6YvMX1EZRU2jNrJx/rSWXbs1HX779RsuIWKarP4MmpY3v/6dvghBa4NXBeoKMqh0sAs0lTXl
HUtaFx49T2i7ebRzXBqmLrU4ZRO726gBe/Gifp6WnuHwYRqAoMyDonVV5qs1QQGUGtM0n9KaPwsH
MyFoybhAlU8fPx2Ps1X0KDSKirba7QKeEYTryJzCxMUxrM9tHsudIZjhItD5Wfw00MGlCxEMkHap
6WxtbQs/LJRh0UN6RAVKymnitghwzaQyfx4LLIvZ69+TgX9Nee+k68D6vzZ/b+N3HSOHUR5Ye2On
ZIBxiZgbHxbd+2zRb9A7S7xPgjRnieZr1YbsCPVdvCzDO5VzdAJvKSVjuUIOhnZ++JyyaHEanCg7
qlCWy/vbvEtd4/Zt2sROiReinp2+nAVRpfZLYVioUHoKUnao+SRqGcIBLTZKl5GcBfqsuZNHO2It
Vo+e+L0nUk9vWFNRd1JM5EBhfhtetgJ6tYkCvxEG17cgqySkHFc0xCpSTOAenNhhiRibC8jPNqLI
zo2iS2AQAZAwkwVNu3nmjNuEObkGIxGTLHcoxRpGD9VpKPr0KjRTSdGHOvdfiJEre35GtGILce4k
YRJq4tKO1F/2YcLx6pJKtpMWxqlBmYFoZsLndv3gPph4opNpEsamdXWC/FDkDB/UzvLCVkxg81MV
ChHcMXKpykufjieGsRe6FHqqEPqp9ZSoB9qh4v6927K+T1SCnFHGUVqJ6iGwI2A2NuHKWuSUIQnw
XSe0OI4MkpaRJ7S/VC+uG0+o6gPcDbklSQRFFudED3bscrun5JaJse9q722zPUIp8JJTVd19CENg
vSzEP9QzsfV0wBH5drPBGj/Sn9rOkkzFo9fmmfGN1w+HUGZs6nQWbIc4OuX3mCeSTr0um5kjmDPw
4zyRITXJgoUyEYt3L1Wl8jGvWd9aK/wOqQP1MswT2FMT3OU5M57+HWp2nE1LDmefE8isTFNsmtwc
MIxBXkYOgN+F95/GwectSp911wtvF8VgPPpMowHSCPRFIqb38zWKGEfgR97i+69tzGP7LpMvlGYz
FthPEajP1l39+YShXzKmeo4xZD5lt4ugr/wTu9IQsAmXAJKljaqIJHG44rgFyw51J7G24dPSmi3Q
V362hvT8sMg22K52t5CLfvj3hLvQdbDssHYT/h/8XFCqs2HiovRIexE1v2aO321SMnmDPp3y4SKv
NkmXb6pkbPC5MY6xjftzN/1Dgi0sxJrFFfccnAc4g5lNq4Jx9QOiT4z1D00LHtIciS75J1vi0D4H
+YoLG5GUGLG1eMT8TSZ6nG2w8oRXUqO17AxN1IWhOztx0ZPHIrVw11856iYAk5Xsx+2vp5aImjIU
Bjqz56FhsIye6SBZ3/JTw7TuY5QAV+CnaAAl6gDQWuOuoS4AT22v2N/R+2YIgm/EhJr+KfYaIL2b
n8GIAccTL8bRO9nTtPkZWtRxJ4Njbincw4crtXD1/uiS7SzQSgr8LiejyXbf0k3MO7urKqHvp2TY
5S2p66zA7T/h5selonPUpQUpofCs4q2Kjvn3NV1Xa1YvrVa49nSkKCXi53uB04YuKBAGnKMJdYCO
1DtS+x6r2fTucKmSOSmY1QOzzBzAwAFGkduSMPGyja5Kvk2fXOCCoPyQc39FF29DrJ2imXrscSGO
B2+XecFp/A3Wpx+GRAUVjZlEGPUr8I8FxxBVj42VmEZB0oP/I2yDHSyVS4pqLxRjqXMfFZK6vLSm
kJY/nbZ8Qhjj2PaFO2WPhsunov154cNibp6+IloUQbaCKw8m9RuxpUCTcrGSeY9AWNjAXT8ZFA/N
imB4Sc+575BJTKTfmUXszBp39PLwxsbfUlnVKSWhQlvS/lZPGO4UlV9ogIoD5gvNxBcd0FqrZauQ
D0kHPaPZDjgmDjWV+i4qYQAZwFngrM0lOJrIEoCqE6+pPkPvX57OPTGgjHe0LkphLc/Slhb1FyXA
x9GlS+yDwj0CD15OmwBBTO+ezF0YMTXbQXAxsyMlR+c0jcEpu4+05Yn4O4hgs+CbezM7fORYcF0S
rOb6q24SxYfrO+r7Z03/n34QR4gfM9urPM6IEhHI8geVooqHo36ASM1iVJcWFehdEA4y0uKIhNgW
PFC07pZFt17il1+JBOtRWQHEVwDiqQiKGU7GLhOIRT4M8g3Im2JsdUTWFEYs2gfpTk3U7M0WjMTx
mtHi2uIBvvRefd7GEFYS5YARz91lzehDp+YqTWAPDbkZIDYkZ1OYKXCJwBmNS30iEg9sJQeH35Sy
abgopx8W19dWwligUV/8p/Dr/YFEnR6wyV7LouKRY4Dt+r0iTrGgUEbgbbavSUXuRrsl7NZ1x+uA
CuRTCT/QW2ioP0WUL6nRmjYqJfmoOVyIGWRVWg6dUoW27NSs2+O5KcqRAMks7ZcON70WhqsGzDl+
CHxo19gIp5IT0uE4KkBDZPZt3Jq4zsKHjMIlCcdvRvst7qjKZJg7GJp3sHT1la9rqAx6YfLqyHk4
zNjfNwU8hUN7e1l2Nxzo3X4SkKTFxuZ/MVoH3skFNjcYXqeSONT5mBkfAwao/sBZyrFZApiUE0la
mb1fqeswwfyrZHmuiN8AYzalhHFwrkwbFVL1ONXKqyeEAf3MOmku/8J1MLi4Cv/ZLwO3EkzyVTe9
ZW+9SR8smx0oDFLreBBOiUv20XEbxpLL03c/U+hIaoz6qm0bUHWXIdES1aODOWJv9Rfx22nC4Go4
Y8XlY5hyCE/NRAmb24qVBbAUv+nNbclcD73q5cpCW210DC5Jsbi5VQkzHJsp5HStZRcfK/Gyc8xb
LIEffPOioTZDst9jVm9Wdvv+KlJiZpRRRmRjeIR2DNBbgCvISzbIVDK7JG6V1GKNAy/mjRDodVWr
4W0sOiRO+h2SziOuhDDJzGp31PnTk7wUxHs1wxZODu8RyfeCeLZUNUavk07ahldFRMpPHzjPq00L
DAKmfUoQRM1a+A9bK04iQEZiDH2awqNkruhtbwECpitmjpXW712MXcGVkSBppgpnCTMzR4oZyHBx
S1o4MKCc37qFr6fh0DfAB6QxD9x0J7Q7++z9Rbbuum93TGWd5iv0b/Encuyw8SAcfA+JAmxXlHjQ
gzmtNiz29HMbbPGbOGjT8ZKbDF9Yw9lCQ/DN+T1PaViQAYqRCseHTOmcpjXeTMjux7LTqpRqk/6p
An5ByRaPvIN9ghbKy3SmtgKqZFsREhcedPgbk2tUkY6rdW55oMbrz/8ynFrjvyY0bVVg6zsCb8Bf
T93P7YGAbQ6wD4D0TP5nAzimON8DPIDk3gakvS6SvVKAxS/wG7ominYAyagftfn4CJ8CQYaeYDmw
Eixy16XBuxuIvnBpoyJOwErlTIghu0QjoSN7cLD+kFmDYHPfRDHoAX+oyZaIiFkzmOggu2OiJjx1
EQ+GB48GX2FxBaXkzboIpAj6fK4r9XO4MHvk/zjvB9FzrGNf9OiOupXfUGIzQxz66+WEpKX+/30p
YKhxVT1+n2w6WX9y1oMgAb/gI03caW8qhGxknPaN01StwubYYIw5NDsQYHFP10jRU2uarAAI1/qY
5ppWI7i1kVU0WB4+Fcj4BcX/69q9QssaovO2v6G+vLM1fW6Dab7myDc9N4cRq+mLiEKePzrFf1Y2
4avKkGbZ+fDtZ5rdZg6YXoLhl6K2eNXum0WBtWt8E/5bnkZd/S1fQKnYKXtjxk5s4ieU5etci5X8
phuAggRPx7YOlOnVfW6M1K5hMGIVVF1VlQIiMwWN4vhGaFjSQK+KKdAlpy+GigRN8lnNbcHM1gKY
dTKhl9FL8du1YcSJR8jjN+5PRvgbFTg0S0LzDZFM0Nq1q6QpPdfkLLEug4km5PclhwT8e+TBH04i
za2hKu/NBNXN8zBIiiqRfOLFjCs8BM4IxrE7Q7TRukP4fIIQv+WDGA2T/LGqbgTM+Q+cQt3ZAFz7
laeWMi7MFpuzx1+64Rd0gqmOLualSXXWjU8cVaNP37xP/htGWcjrNCUgqI+r1B43DD8J6lSg7gL/
5G6z2huO+VbC5hluiLEq/xOi97yEkpu7Q/d5PobXjmsrnZum0VmWAxRc6k1xI5O+ay91m3DW+HVr
ndtNutTO28+g73lV0Z56NBxQ2wRkm0V2Gd3qUR3Hlavk83IL9/rikvrAYggdlT84QP+LgOBSW6o1
GO871uWM5MDhfEfRVDeN2gLmzvdged/A6h/gOU+/LwgwP1fzzWiDqcm76B1Xggjp5rk2rMqo7wZ7
rGImhcq5Mu6BQB292kUuWkVjLQAdQUo2ApoET85ny58Zb9Kacyogq7nGLk17kM9Cy8QjrsaVVJvD
0qhkKoAFGAXpWC9dj7Hluv3W++XySA4hk+UAoqmBCEEhvJU0tOA3TUb6SaX58+xa6Z9s+TMkzwXt
Z8F1EcUSITaDduN/cASu9dnBby3J6sY8agfVe466VsOnFlm1zrioZpKgtzCeYcApq2CCU3NxNBCu
ZWng/vX0ryw2fk7r93uWF0hwUCM3iWJGU5XhNZaWThXaNuqJqp96x8CowojSWqPBc1JdWSlfyt93
jfHnf9EoRF7peOlVm6CHU1qrBLreaLk8oyCMUBukSeIX/8AKEmynexQJZrJiUUVgIzYvy5HWousd
hSbiChoEBjZrq6fYS+dgzzAgMkVHYwzYif63ANTbgjWAFHcod8Gb3w1wUvYOTuqDBaO/plzMLWiQ
YmEX/BBQrh0P73NX6bMqxxo1r1by1IVdQeHf7VsWGndTP4BbVMjvpmk2hOYN++tj8yJE4hOKNrkG
SMENNU83PPBbblWsJsn1VE2XGeGfoB0UYcy3gVhVeNMHLada3G3BmURtLJ2oX5iXIspN74pzjcbG
wwTXwmpOB10C1Yi9YJHJiu2z3nL7w6Y+KGm3ZBLhILYyT4UMWSc44mKFPXEVUlWsmlZnJCQscoVt
EqA56QQfTIBv6UPFW4epv+T+B8VuDPZ32960kQDYsw/+luVooZbWHMdWGLbp0SITYJaqqnWW7j9r
FvhZW3gYXUSjVF6gmVj8hKU+rBCNNLVK5lfima4N1Ekqi2TWm79xce8u/shEvCbco9YnPxilqalF
9kguz0o+bQCaTHoNdwAivt5CNnRCAOekh7VfFa5vLWr4rnKpLIn0UVVhzTdcEN4JJ1Xi3wa7waz8
o+kvexHOQepdJ52BENqjJa3MpIiJHuoFSLpfWaqKhbauuxK9wo7WqlrMeDMhtrZ3s6VyY9YUfifh
2IjcimZdE0cfzrBpA5bnAn7+u11nLU+oxiDUpfH7BgmpH970RW9L4urZYU/89eM8crnOAyxCcTtN
XLMipfBthkd5gMsSeHabcR+itr/zfNCszEnWTQ0UsHPuWB8pp0wW58ScRkF21MRNQifVIRF3Gh9L
BOwyfY2C0h0tMmhG374UCQKZ85j0qTSZ8q8XBJLt4W40MHTa4pZdy+h7MesJ9JeD5tW+BIdch9fJ
YQeNZFYEQdpx152hbrkPWzJdQyMbk601O1NyaLwXCEmA0xWFl2BYsRAZxucBzL2+AyrRqwIHZtPZ
W5+oHiuCucIIxYjfFea6XY5Tj6dzdx8Nb83oDgOTGtfYHOh4+DbLqB9cb1aSnoELW5vESDTqhnWv
z/vsmTmLj/ywblViTgV16M/dXW1YJXLZDedPzDXcjG5CSRVQXrq8sF3Tg4Bl62qlcoGiICUIyKzC
90kxm2YnZDC6EwvtEuwHbI5nq1t3FqRy1ltx63T9wU9RRSdlk20JqOdEuA8+RB3Wy1M52f+Z2CV+
ktVddTGCTtTNXHHiFpHQkx0dmHoi01YefsC2xCmh0oSUTVWuoB01N8LNWy5RL/Lk3Fz/J+oEmlse
9p6BPDpXAA35FoQzWXC9WR5fC+1bXz7NDaHpbCkpPNRn946jaGj9+dBC3ay7I8VLcq+9wwzwvCxF
Bx1C2pv9el1OCAmjDwN30y2YfC1ukCJaH6rhaDGHrGI6LI/OFVJdbBk3jSegacVI7/ELLA1ZvoOn
uk5xBD8h7YSVj61cfxnEg0C8FJYbhyPRLX1a6nB49b00gON6e/BiuzH/Adt7lYuLxqwhXY5UZ7Sx
ozIMVeF78Q4uZD3f5iTbX9ceKWTJw7M2OfGaUi1TYWrQn26x84MrllLQf7uQvVIrG2fJZPz0d4t1
VuDAxXlKfJRG/NXrZ+p0yNC/TH3e/yFd51PXdloGHiQc98ODYO4Tv+xkdYG2owatkAwNpL88VXk4
vNgAoZUYRVc1zfHtASIrC2ytMSv6KGsV4W2nkwjWkaP8h4uP8M3P5T3ksnwwqNlQXsxb0fY2Mqz1
h89EkXK4deurIfd2IUEJmqU7O0g67MArvHXtdxakqSICrDkQn0F2YrPlVba/zZdXuRXrkraIEgn1
uSuTc4l5e02dlMYcLRbCPdKxHKCB9Gtau2iPUuxoK4pOGC9Shz4v5h56g31UBha6QWDHnp/2aoDf
YG/+W+V6SDh/3valiISNGfgBaKBc1C6SqZSZ258eRaJspo2MoJbgGj23ynDpSq8aa475HFXbdUdp
OK4WKQ68NuTSbJv4YtKx4LekAPIVtKLHq5bFR/mfSbV2/3JNAdqaqAx1QjslwhYi8WbmBnzXRdNY
cfjkzHpa4JaVotTec23p9ASHmXq7337pPr7htqZykTguAfwmZpVBwMFXyAxRozi9zcTpdPpioazX
eLs8EFPXux8iIO2Ygkwe+BZnImluxHD093/gf6kCizUsQpu+kBsqdpZKgBV9UNNGNCETDo9AZcIh
uYWDjGqTn5EHOVq1NeXelo2mpI5TeJeF24QUtXsRzUto7lOPacYq4Sd7SoyO3UOP5kCSq/a1FPJO
lPIJdBJV/wnysWAZyFhPTumbGvKIwvKWXlUreS9UUDWp4iS0wUgUByAmhMGhFCQ+3AHOs87Plqpr
Ay5LCSxbqjxn8Cy/0buOiLr+8Oi785fBBOgl1K2oIQ+7ylltvkQUQZq0gl/F+5itrob3DV80NLD7
3LYgpiYHkbBbXn/X9rHYta7hVdaaG0xPp7uo657FsoCSPUQicL9n7WHb0fSpwB5EtHPTn2/aotmE
EIUxlR6lZzACChSN639isUslMtF77y8IDUZ9+myE6zVwS5qcL20Zk19qnZe/FIv0B5flaWs9yLzi
SnVjVKAfI2l/66BPFSFx2IVjeTWuMVvoBo8hfhNe4RNr21WyFUoBPl3mtONy2Y9/5IMQFs8CCWwL
nea+86p8cDd5sQ/CAQoBO5Zb9JW5X/xDLhOMfPv2nfm9jSh5xZijiT9dRKRv8kh2Y/9VluidmGOX
V56nSF0Q83o6ajdM2FeRv1dLpTMKpo9/zqewHfJMou0BEZpWnOJ5BYxIJ9NxCFhkewmVX1SQS55G
URM0gGs7VZSeStcYVOYdqKH4miRIclx2CYjLoustTk1zowoQyITQMefSW/Ldzgyx4kOAOrf4Ck4E
dA8PhvEk5kpHNjFjQBg9zrRmpBqpEpQfOcWGHdLRZyDbQtim574j/nb9UJMEjfwkISMF6LMmGCEE
ehKNfkV3dB4WzH5RN7/zQ6wKVTPqfJOluFWa5TvBLsdvPVB81ZsQb6OzkTaMlTHNuhIydUtQaMo8
GL/E8qZwhUEVFMJ5BFjSxiYG5IIP3rffFcTt614CtdvsStYw3YB72yL5cQbxEHJlJTFGyeN97iNt
19wNU3Jte+cAvzU/EIGERzTN6Cr4b9m0rgujsTBTlj3X//L44v8OXKbJ1hhPWJUfU06d///g1rHT
uZKK/PsTOIixArxmPuNlVtrxUQ+wJO5Kz2vse+7U4Bj9jTmSKfpaWiuS5kkgwJVx5K4jyS1/SFp9
DZh0gKNRAOSwEyFe+7jfb6wj1Z6cq+8s+jF3pOOPT+VjmZFzVODwsPdwPEFmH+Jnc2Z65ZC1sOMb
4741DE1u7yTsThBub1KAPcJdHktPa3TH+Z+zwvAGSHU04CEqIbenODnppVGl+OtnAoQgiNDcrxwf
x9kj6n2JnfZ4tCrnmag6FhKdw7akIwolELgU4ipcxpDBKl1w3snaqzh21YAy+PqmbzfE18JP2Ywu
VN1+4564xJwvUbB3DvGZYCmpwtuQg0H1M+2P+ZUJL/ALBXOMvQHXTn+0GF+BxxxWKP7rXxlbd96G
/jKnrb3bmxqUeHJMOUfUrO3W8ruPop4meQaykgIYaboJ+27N2Dsss2Yj8VQTxKl51RvrIUWKtQQG
zVhYtYrcoguLztDPTVzaWyb4oY0STC5RmTS6FLf8QDFhOJiwqtjZ5Af8bsNA6+M1tpVh0gZIocBx
mRUGutlDQUSfT8zh22lAFJIzBr5sPlF681WfE94rUVpx8S+qbqDavbqHFJgvTPdNV7Dv4kKsq1La
/L0JVZTtGB/R0D1k7bT+1XquYh1iKUdVTv/lSmuh1IxXZxz0K7oSUuGMZJ0QuxqrO7UHcvDo0dRf
W/7G9HHz371+4tfv7CDZ+vOSVFSXBu8k4Lz+iCppXhCxWR5vGhtxqgO4GIU0hEcngSsJFqw0nxUc
Q74cqPCI1WxwWiQ/aiurzTNC1TQkhVx/rH/SstQTHZuWIMMfehmT1pqCOSMyPt6lm34BOcYX+dWe
HxI1LMOhwmC3EzsOU5q5uPJ5GQLPgSLCCy3g73sCEQCMn4HObgx7SEyILykSe8l6Zh3oGEC2Ikpv
U+L3Cv+7Lnadb8DN6vlbcF84i/kQkgJ/1cjCND+3cqjKwuonUTUXzEg7s0b+o679KNv1tMpkfQTZ
IcSFwPxGsf+17228lCX3FyJ7k6CWKPrw5N4RfM00meFYOhjdVwUex2OefB3RdRfHJFe/7WWQUs/b
fzemaN5ktXG2mFVSzQ+uGCyghQx8MxPyDBP3p4ypCL+oSe9VFh2BfuRtUFUaQJAFBY1lJmNs+IDQ
4mUStOXUL1BkYiUE9lDpJuzz9t4uiOYgO7K4fUUHfTqtb8ZP0iOAnMKsnYr7FyK0bzTSxEo+ic0J
uuydvk6EO/dOVy1fD3Ce3TSfWhuiSkTVJXl0+sZMW9SI2MJxVaToiqOA5JQlQlxGqgrkRiF2+Q+l
1A7Tv2SQU+zVCB25Kfy6FdhKzmNW/7FZhgtlSIBqYPXkRK9h+nXliIJW9avBvetq1QDPEwSK/UaO
92sY5wGCywnh2QsPe8ZyV5aJfaBa9XvNBjACkwUlKsnLXYKxZhbCs8XCvhduNSp7RtMfpxRhm9BU
7V4d9j/xt2grBJZbwEcKVRr1Gv3YuoDb9iMw10E6Mc1d2yZaGv/EdEFMqhPDiVFYNWdQF/m1vmVa
/M5+sAGLEMPdY+3sNXgSxEJ9DfLnfMmc4qS5G8QQUC3iMwlxwr6Vf4AKKzBqshCiozXi34CbxCrq
b5WFuXV4d5n1musp9aPHddeDuUoVeOTbggr1SCPAvAh6EclaboOqmfxdG17rpYls86fF/mG9kxxH
PbtkaUTg0tHiFoVCoFNN+GLF3rL+o74uIeQSyWnU4rZfdZdBbLv5s5/krRVsZGW2XVqqpl6OOzl6
r69ZtmjK6UlRM3II4cbfAn+bd1Tz/S0JCJLcrQJGkb06KnZ4eANmT3psHypK1yuH+7mVoy1dE/hH
B6pa1eYrTshU85aXzYpCvXNf4ydCpWo7WL3CUlNHaUD6HIs+3YvNyvtX7Up4c8de4k+V4lUNVy5l
DuGVyljGSm4dRdGCeRCbNuaBo8jDnXo3uch+U9yp6WjufNLhgDQa+G4/6HzwTDZSyVy2Zs1XrIM0
IUzB7Fp5JKJ52jvsQFeq3ELbZ5dEZkmIJxMEJ7noV6oe/rj2G0WFkZT6RlFEY1mcYxka9VivnCiJ
/L5FnMH3SV5SLhDLiVd9eMBcg8hM9S5AHDZQVHE5eP3+GE2UbRbZXxjc/UPkI3gkCNCL/NY7YTn2
TKUghn5VClJRPlrqd0cleb5eywz5E6irBOipw9NTOCYXZdE1OfKf5Ovjny9kpdZxmFMph19bhJyl
M0xgba652ThJu0jGwULMV6IJFL8ifrxTttA87N5WFQn0OXDAtzerE9v6NMJ4ULzYuWapvzgNmy3S
RYXRB++EF9MaSV72Itub0zmGzkiU5WN1494iDHSKAsFHPWfzgAsyiwrz6vDIjn+jiw8S9MpRqGuC
qNcbEE02iX4WQQIq28Fiq0onCl6tH8XwZlk9n7gdS3Aq+Mxilhy0OndhuwL9exRbKEw2NzujDyET
ZhMMoHO+U17f9Imd2z+UBVOdb/X6v0qXU3uF0sweIHJfPVaZQRKMB69vzQK64OMtwIdUUtFUoDB3
0YCC9XRcgQMcfMXjwpxKn1A6XaqJY6x3VG1rletNgGanqY/XbQb4ulqfjcxNcDR4w6//35ilA1op
e/Mo5Z87J9Oe/tGfgpR8G1CXV28ENDIMTDWUgjhzSjdXQYPCevAi3rwhjJcVKvy1OhPQOigJZgPo
eazpVetBd007DyZQnz4jVZ+P/RSGYI+/veF4DKeDcBQr8GJp4werI7lB49AcxcwlLufA8+Wlmh96
RIz2MN206sjNo2xU2jMEK9Op8sAc4YefchLvnN4/0mVolzGOIEqzlggXChADfaD7AoA89D9VfQ/3
0BR3pNrGwS5yx1HitvMS6b1Vi5i7Dd/MPVPVbXZM8UZUFogyYsPTgzieZ2UskaiYFEbugUYQGuCD
j2nfC26n/ic3bDEIJWpp/p3cO97KryeXauSzkIt0pN2v7CAUvbwGolml0aKIwGp2TkBtEq3rodJd
zMPEYOGf3J7uAshmtFKYMkJr1avH2/LvWI2mOE8eWZierHIKZdBWJD+vgwCro2cnpdBZpgQH0B0C
gG0oV4ixVNf2ckQEYYIAzTqjwU+Uoq+5FYyQePStwk8+hLDnn2soIONKoCVgiGaQtXgYc7Z8TQUr
1XTyBtg9/GKIWLz0wJDLMxRHjHpbhLgx23IVhZbZWMbINVrxtZABPx7am2KirGCPs+JG3psI4Q2+
x3zKJ4DXWBR4+n7Vt0jWJLcNeiHKcyfFQTiSPxf3RST6tts1/Qx2WhjAzES1P7CWJovtxjo6NGpt
4DsgElXWK0FoTPO0LVfhs57zb+0l4Htoq44fHv03bHFkzI24XyOelWGihDKc++EYLv0bnTtTUkZH
3/eFgCnS0+hCV5lLpyR9RUq2EIBK2GpPCJaZLoQy6h1pnyl3YXIvTytMJcj4/9qQZJ1MWSuS5sNM
lfaM5guYAlP0ZZeGhJBwqysVPPQDR0WWjzEAJMLVgkJVmO8fDx7fwfhd8M9464N/39Rq2+T3SimK
WE5kdGyafV7PuuzQirZ8b1oT4pmrBMIkhMx1RSClMr8493yEmr8Cl0CeSrajC9Lys2RKcBN6sqzX
+c4hEmwh6TS/v9BmGxWURaC8gc34n2KWHsku85PTlah0oc3TpMbCTh5IYferhBlcUZISUMdIJ+p+
bgMRv8PbQA8YNMwUUPZZOfCrFx3ToNew3vI5YnHgawzR+b7By4a050tYqjJ3kSRNvwoi1xq73rgY
W2zCJ4Id/mku/4yQomyqtVn7dudOfu4c/0Y9M217jEaobwdNEOdmBldyPX2GifIutk5Ue1QuAwic
ZyXYAmUk6ZCjsZ3gd1jsM6Ogx3cp+GBQiaznsbNswdOaQTNpKvuntwpUtevu4lcdFv4KgW+m0W3u
6gsW11BrtBBYHhBWL1YUAYyHllunZcdrdCln8813ffcqJrYev3DWUAZkIQ3YhQ7uoakszIdX0Vdy
KHLQGSG7tunTQ3TqpRSac5EaSgXwA4Qq61asqmoeZjvxr5xpKQZL3M/dMlDOLEvBkqHdQTb4T1uS
SwvqRs5nUgpM9KptKtFyfDMVaJBd+9HeHIEvrpDOSFLuKOHi6caNTSbD4vfi0tDsxiVU9wsTcOqP
tlz2sA3LUoPlsY/LsQo6YRzBcTYykkzTwoDs4qSqU+KVeIkRxxWXaR1Q45HbCCAqO0drDgZuRFNW
FxUjgNp67fTMz4B5sOn1hEl9n6W6+lOnwO3hPGMMKMr5j1dztoTwPBpaSwhJJ3lD2UBv3uactNhJ
hISpheZvDdrm6cg+/+VBBomg4b9dtsY9Dh6HeKqdajcizieEGdKWxBS1QVGZA2udH9BUkyoy1tlN
65LsfHqkJvJ+Xfa2jtBzKIB8Qh8fK5bBDN6jPIAmWMO+Cut6RC6l0hBW2J109Q7oNxRDZpPxZaVo
Wuq8G/UzbVmM31B0kwnGLBJCwzrhj08CpL1wVwGil74ZUScAkTNJ4I5/BskzdxaC4eX3rx/hS0yH
CLDVQIBQ2xk9/R3UDnjK8L8TY3TU+B/cQx2q/AXQe1jVIilG4P8Zgbr1/wKMxzMffdGwlC8BLq96
9BIAuifTyDEboRiphbn1rQNWeDFTiIZ+zUwQ2Sqrv1LIn81Lz+rp7eqGgh2gOCcOK+0FndtB2DQF
OdzssG70Xjo26D+vFJmiPj0DvcG1EcucEeUdkjpkRY81pimk2OmKKATDxMZ4Kksov5IAWKgW+bWE
6E48akhx1qUdEfhee2GTZ5OMQqWNu+HmfVq3+gZ4BOKfKilOY/fTTakU0fyqu1/yu6nP0gTIEbyz
W+yDRsPgFlSmkAA4xR2tGdnE+Y9UOUlOqyY8X5YVjsdUSz1jVNGWVOVwAflve82CnReJIIhjuYd3
6GmGwBygYVFOTXQQ0aLs0zu1F6o1zJ06XwzcUHeViAXVkb9SRjEx29xBoOmUsgmMO3TqJZ9iqanl
u6AzwHPz+K4r45XpbFmrVpvoOB91ndjLJSuonoLj7l9mvtfvA321WrFj/1y/10WHqYzQkLSotyV5
DfaGtcOy8wyYY0JC1QENElv3diw2Qr831T5tjU1kRud7lh3oMLyyOQZ/+OjxA1UZJ5t5Ez4kN2WI
4LH/wWieu+wAnCwaWFAIFpjnKkondsXVfQlruVp+g4iJxJO8oO1c9DBxUfo9q8bTXbtFsPtWnxk9
VJfPknzfn6SoM5IoquOtJ7BaTSG3RYkdgxBlNNnPgx90Yqtb0uv5KXTAqSGpSPWWOuDzsJ9dZLLT
3T/ve2RXtxGGF9B3pHO32n5D0o6Vo8Hc3lSdUJbiHb1NiQp/y8a6BwAWsQjwM86gwbjGhdJq0Zdq
3t1hujKwoZIzRmm+oUYAWlHBcZaA/fBWZnK70PC00nZzHmGJcnTxGtIWP2UZnZaLCowAK56ZP7dP
jkLj7Xm1kQvyyLVwzHvCpAh6qFlrsUYcUuklojHAMTkO7aQuwWWNwsBLwTQ8mNV1dg6yphZ27L3q
IIw2fBFCGpxjZqRX0j8fCS0v5UDlmuAEerAY/ka/XG6N6bLAqYQBhwwP6fIsoGfEdYr/F43a172/
G3HqTrSWCc30/nXuincOgRNc8yIpPIvZcatCy4GeW+pObiEQsdrDkdVLE7kVzxU3zFIJkUqSBnGk
fer7g3D1ECcOoZ+Twsz0ahgqZCA5KEkVwLoiLflhbWflCwSiEzNGMXBIWR/7/EAPP9HY7wkviFe0
65s4+V4qDbE9hmIgVDQ9Q2dzbx55wAY7RCTW7Ck6g7GJJxB3Pp/m/U9Guy0gsLZJNwMQX7EiIBHF
9lbYSSH74QQTSWAc97/LtfQ7fiA1IZDQTrQputDCTY/dwzpxiXObSKr1wOmOYcHLVXEUP0hZREB7
3M1ilV5PyC6qPErZ7TyqDMdKg8YLRMHKJZKUefXmGFdIxhSJ0V5EVXTWymmue67HkqTPeZeHYp03
7kMGDO3k5nlf9X+mEfg/gtsiHMx3I2zcaxZZEDs7UrdwwqyL5kbagfubbZf2Cq+ko8vc6HnRFTJg
8F811lX4aVriD+DIzM3T/XvsVSBu3ffkXWgtFQcrlbP4xuDQ0+5Lajwo2QrLSKHyoT0ucIdPxIzh
RrYyJXwBYKuHlmRtKIEE0HIFmg5FF0F1IfGw+v+KbMePn2pvFh0oCYy3Eec8lzRyURyCCUoLqKlP
0GzDjHDmBgQEURsJn2TH6wVrnGnXni3ymwX6GFfW71w45H+fBR35uouM8HjWCdFxv7ACXNuMZrC2
vmnPnPROSZiS8tLuFe/FIHzD+yuPKj4+Ycmg4lYu0ZcDYnvh7VPDqLQDqHhRv/WWc2IeFJ01P/D/
6SRStBKKHSlDj1d9x1nhrrEX35e32wVlM1dINQfX0GDzRfwlvguPe+mObE5AO6hnIkyWy/gerLZi
VjrGMh4xIR1vEzt4ykoYdP7hU2zR997l/jCqz2a8DfMtu4wQBKEEA7EXHl8eInAu0VWlvemmlGiJ
5ScgYK0R6Ln++URQDHkLeFa+rdzV4ViATNUfXgbnOLs/jXbsZdXvmL7YVWqknLuswEdTn2vuV2eo
rf7RfNxG3gD2t4a34V9Wk9a+Ms9iG2BZa58sGFUrsaSi/3KPsW5eql7UYqn/laResVJMw58vcLVE
vmb9iCg/dWqmQExRot97DfbJjATNru11vNZIXwL79kOpThunmz/mVh8TNIwg4bn+Bfow4x1/gkOm
M4SCemkxgiczwJ9hYxBOlpCTX6mDECaQEWKLun8RbG4v/zQr+K+V08L7j9gWycwBBJ8/0nl80Gzs
HjJj1RZM4Eo4KK6D/f+N6QeO4EFrXTpmKc1620I5sX98FkaFr5R1cy3W2fSrS2Q4oPiz7UhP48FB
3LdRoNqAFLZC65FwGNn1fZxg55gQSJcQxuoSy7n8qT3lcRNfNu5+NwenDW4oVvis1b0NkOp5qE0V
qC+ujdTxSYzWwlzJimUCQ/3nBgc6Aw4JGOWSkEM9AFTETtlIXIm6ygEOAk+mvzfIgatOAFArXxvA
nCfrGvjgKcqMRzfV590pKugFhGPYKcWCBVgDj8cAuLQzhZzlx5ZY7ezykXwhbC87zNJ2I/Q2FNGA
6TGrAhaL6WY/kuTQ2f8T501U7o+zzmf+p//ve785PqD+QcwSpb06xUGF70frB0e8h/lD8Dfggrsz
9lnZrZSWPR7OXoEruzL9GRrQ2ccrCqB+c2oVP3n2/P7KzZtj6nHrdbMBKaI8ga/mChyUQXPIfWmE
BwnQyPREANPXrciEb5lSBrG7wwTLbsEKF9518EsevY61ziD/tLHXQZ+bOJxXS1efMIICQX57E0UO
40sJ+GVo1ZnTx7wehhklAavvomsFlUZvZyem/x95oqC0U7Yb+ONQTt1Q9w0rXLzCcQ0JhCVDKk9q
UVmBRZTwovaYqG+O/YCZNDRvEefiUFH6/OyZaXNk+ORq8/QI0wWaB6riU7H4XHITVxawkujCBRg6
6DI0X4EVDzf4sRroeIor6KeQIYot1qMa0EouHcx8mXRXXooG+AomRXyBl/23Gn5YryzkOGlCS/4F
/ZyF68y0J1VIiyQVxC75Mbu81wGwcr4Pz4Uku+Eu/PWAtacFj4ESDUd4ZmNd4eM55fGufLTpKPSZ
txfmPnhfZ7DEZ6bCxJB/uuZehVCgTbIGCEGvWq68RLb920cGa591rZn/cH8n7dLKOICuRpG0NM25
bpc5C/vIpwEBDkoS3Asvs3w4XuPL56J7GovuMPVUlCuWpGXPXAdRXp8cqCtNsJ18Ii51biaRH2F3
WjYZmWwabcFgudMLYNsHqGrguwY8c9p+uxMZ3kWjvXRcIQ9cwUoB7mzO/wzzj9ibdVfTujKuIgSF
8k0qZh10twQygAMvpe3EaMWGvXl73SiaeNYZfPOPEAhcA9WB9/2wX8+R/cG/CQRovBCgs62S2uwG
W7zg5NzFQr8rDmMqwvcBz1YTSZSgevPhZZ/P4fEz8l997rFVPHGrnisg4I1GvKaSu1sesxDDU6tN
Yt9uwq/JT/U1hIKOlHCe9fy4Tp0KVKOVM0w1he+oGMa2D1dHNYreQMObaczvlb2m4eERA2GTdbTP
yEnocDuFVdRu7I38yamWTCN6mwgT/IDh0B88ZLGdtx+6UUmgmnNp21PHg2dDU2Ib99ybUCb1nBf2
tJkLLPYx0GW8iKyJUpXo5wBG5clMPSK+PaG9sPeA+zlFCIxXn21awwxZi+ZE2A7savYjED97z4Ip
u3L8LuXfIy51wwnYeKbl+sVd1vuPYk4KieJyoxLNT+ETfhAjcNfYWCY1eQ4iGhcttbiB9xxHTtzH
kzuI2pSsdDI238gRLjHRvpLueX41k0UPiqAYBuSG7XXhU65D5pLK+fas5AbbfCyixVrm0iPQeCTj
tfZ7pD0EsuzfMOt4HuwLidkHKvaQrDosLXxnNB5bf5vzMjeqKBbA7XeOrY9h9Qs+Hiw5YKufgvSP
3vCp1QJgOKS6CB9tKFITfh0bLc+uZ6PRAdkVjGA+0BQ9D4mLO23vUIr4/eFnzhwbeE6PU7DT4dIj
jPMBdVatosSdn3Q+9T0gcV42BvdS1q4Zx3X+tGDYHdodmLodkpUqGz2O+BsHYO7+/T01jfvayUvY
JqeI6qo3zcjZUUrYSmpNeRouiQqIBxHrAeRy+PvvW+T6AqRk12y9tEiu5lBRmyTdApbCYpL/AZqY
oin/OV9mDNfSMiFL6Nr2F2JNHNVJtBLJdgMZ16iGLm4eKDUUwes9Ij0hdzID31HSvvinixalkHSU
oyObVY3cVz5t6pWWy3Y6DHH19A7u09nz8NITuZdwN6ZEl5ARpnFlGUocGsb+MDiSLa5XOdOG0Lno
qndTkKiEmSRAjoe7prWkqeamzVTFf3HwqTmhWzOPhy6u4sIqAYUmkFO/6i2Zxh92mAh5J/TTI49F
hsn32cEUFheak3jNqEf37oOrjGbGZKkVpfM848ftJYdKvYYbl1FhPyNo+UYJrMmFmNISQ3D0SgTm
Qab+3t1oAJYtRYp41GWcP8GelIk9a/r+P/vJNFOiPjieFrH9bvMg0RtfgWIz6y3FnxdDjTWAT/mX
7e2tGnoWsazojX3Yh4iIHqMSK/Gb/ETMHBkD7r5Ls7W8ANOk73VpExOA0scLk0P7nPFD8kV+nLRO
LQcOLTqKSroNbURWG1BGplAvYPu2a8ulnvN3US2zhR/lIWNB+2w8EVe8K8bA+4S6OxBvC/jDWOMC
tFQmnFF9D5WQwUefmKvddTNnWwWcxfQvBHs17yefU3dZufLCqPMBmHzjQjrS5Rz154U81zFLvMeX
IEFQO0bGmiXsKIOR/EK2ninSOlHboQ3savIoxoAZp71k3KdNi0O3m+ah9Q4eF5VDrvGXAUb2FnLi
AqLrciC1pIOWyIeHiFWi3o+l8wi0opNJB9d4lIKtGHua80tZ8pRi9PeMuiSBvyICn9jE4gpO1tzF
sbuLhl+zr6tUJeSLrIFH1yl3V13RjNGFjfX12EHCvSBf10UwbJeLqgDY89UUwGRTZUf3QAed/oWp
7TqVhvjEL6c8XsZ1n0mXBGPBbHxychYF/We+kpIPTkxU79UyIapud2p4sA2E4zMn2X6x05A/s9h8
c6Qkxn0yo4xKmTPjzfih0vi4PXRSsGDmdhAPwH7jOANpfbccYW12q1TwVvLHfK/8SXh6mIm9Sziu
sfapnKf9n0QpsgBhIFjWeGa9fIoVsVcpVpC8BTE9lD98NVp+5naSMXde4SyMb9l0BYYSR7bowobg
+RJgwyixWf93uzzTOPJzfT31/9FQmp7rGAVaNqR5xeqFqB9uRP+4xUf0OO5tYop4CYVoxwTQ6t/1
9nL0xxsJm+yqbkX73OEVRIDRAgve1BlEiW82Y1PTUwna0gSdVM+8ikk0t+6uGY/9lELtH27nwyN+
NsBi2VKPXsmrvKZKfqTIQHMjWk3USpPgW5WT+K9kmYmTXQ6ddixj+CTnC7+eFTt50YKxftqBo0VS
+FzADIVpBF2yQ4ZzUUg5S+TG2RYnuezpQkvsvImqCz5IUYy8KbBoPmaEhkp/B5ZJsy7y+Rl3zcaa
DT75G4ygIhJxkMqBlGz5rxJwYFeYEWElk6y3dpwGgCS847O16HP+T09/Hyq+HHCE/4c3l9TWDM5/
Lbr91k/d7tFpXj1zjN/FqXG0GEKlmDRH3Gsvkx8SEnmfZKH9h4NIzXHakNkfAp7+V8ggw6yWnccE
JJBVEWorLlzbDpymbTfB+b+KLRAwv1k8OteZPhwOhldqFsc3IFKSM6Q7cML7Lbzej17OhCLdHb/4
3ExhtEy/1a6+sojg8qeZmgg/fVY9Jy9o7XHkzcJegchOdBMne0LBz8PIdY6LfdMQSVCInnl9mZsE
NXem7cmvnexLAQyUgP1IR3TfQSseZf6ngFb5ANyJGG7BJ5+8xGNx8jiewd1bx9aWIZ8e9O/tmjT1
y19/6b2kBCGmsFSLKxlIzweFjSMl59A/6M/ev/6yPWsHmXI6Wt/Lyhr5UJxJA5KoyMtGJM/hnHL3
+OgL2YTosmsA/8DQu3un9+cxUhiLeb8s4kWbIsiH0hkqv34NVKsO20FpSKwrhCOe3Ey176YTPMJb
bUfO0IOoPFhOp20aiMw9su0PgnrSSyxBqaajshY+KS18IDC1YIYI+xjby2ryxUk+wm7fOAdd9jOm
bgY2yJW1arMjYtyC12QqYWUeNSLvSzUm796XZxHpQFHlojhwP/ncVU9Wyqv+OJOpVemwFB6L9rlD
ZUaWTPwXJ1g699XRVISuONR7txK3U5kO8FDUwRBU/jvbM8TuoA5NPRsrPb2X2/BgpuYqj8DXKXGk
4oDdyBhwYn1gKSBTJaO9fGMdXH/RrMRYtbjyqy11Acv4oi/ESBzd95GxC6WNzSXsCrRk7lBnQRbP
LuURhoGZnlIWPSFMdnHnF/mWcRlLsUUzbj1T5YcLXftqqci7RxPkVvh9OCc6JOPY0sZDwHmlEz7B
a9dC7mSeswI4TEBLWMlQbc+Xz2z6rRUx8kjhIl/C0roL8E/cpElQ4EFpgDEi5Ndysv9bsCVn9nVf
XPQmxPAWBnFFIRu3gr4LuWv8aL5s4rPkyzzl2BFHrY6GI1O8xIOO+JzntFx/9ulXdL6NNGOsf/kj
Q8tBM6nQrpXLiWbPFbD/M4DzW3yD3yxHEzjTqxHE8FBzkwT7Di9s7Qc/mIiu2Bwia/HyiCfrBNaf
BCiljmGrpXMW5d47GAYo8VCRqLKriWX3omqGXioAket2nVClQsZqAdEcdg7SHfcZk/sbI7ZSyFJp
zs0suc/xUlQOz0AAMsWvMpJpXLG86tu1+W0oQmNmsWUGsPWlsQQrYsHXe9R6INr1NcJHjcnBA6V0
X/FD3DS8b07lw4LdE8eX5FqzqQsybFU73gJuMVfdX1NwbWBjcBcRV2oiw1U/NqEvT381ki6uq3Au
FWwrsTotZuQRXgIggVYJcYTI1H7/FnW2wtCCbq/UH0fPCft7XuzFqDczDvjmrgYUAnBwdXf7Ciu1
e++pv4bI5vpIYFGmU5ydLuwrh+sIUtOKHdoLcBjOouyQu8v5NxXFwtgEtBPt1UxkVZKsz4MVxUZL
WAriyBxGrJNIfR9Fs5zznqIJYAhmXAgbOrXP9Dxbtvju46d7aSoAAV9IMwJarYo25k7kaL3EXXhx
CsIWwaVNtSPncE/NdKCVpyRCiXtB3zWP50BpAQrF4SXfVngJytzKXbsxt/rjbTKOTAWC0ICi8x3X
Nx1VmfQWH5P1W2EbtXua2h+YIti/5BGOvo5SWr6GGSNC7Xn5L3jt6kisvPBLTJfwlFfQVm26COap
OtDTLn/tzEds0sRt0PKOo6MzxjuHSE2uSCFg0DM7b12HnLuLNY/LKzEOScDXHnVstAfERxh99lFv
WS0ZF1SMTjAI7RAIFgzhDI/SKGNo0GaA7sJOCAivwEbg+fA5yTQluhYgWic4bTBWpgUgxJiPnP81
fEADm4PMO7XNl0DLFtDMjr5DBWDlcO+N7t8R2itn4R3zS2r549YEPgoe7jt88EL1Hq4Z7rKCtk51
jBvj9W7WVuPZakyHed2aYAawHXatJTeMx+tpMN4uDqqSYRConTbpfyja2oRqitgHsz/3VRynihkK
V0lyIKH1p8tAEPdvpZ8y3fMMN+zLd5yV+r31aQEz+Eml6cBmFWGhLqWGR40sQI+BHZszns8S3kT/
s/7Hi/lKxsaVyoyq22vTMtNgvLVo91nfxTOe3M4Fk+VR0RDauiXn4DHSuYqz5M0sJ2q0gbdIaTwp
4OFyY1tB8MMO/uAJc6NPihPvPy6iGnz5rf7CheQ4wSaV+ar4Y9YeirlU67WUzadaDQQZoCM+s45h
ndmBtwgxFF7l5YuFECPNQvWnklns4DrQP0trIdus4Kk0n6Jq43zGZlVPINFBF6aNvXQoq8L219wZ
6haQ+sVGDWKvEaryIzJIomug9K05ZNg6rUv6BHDj6nlkBYi8sczdLVGYeR7vSFw1Ui7qHxI1AoWX
HbObtAshVTXiDmSfJp5ZfcSXJbBiF8Mu3wKGUyaQNslr77WHKFRyW76nYppL3AmayQwRcWDZqk/L
GpuSb22OGa/bw/pmDHVP+OdH+7z1NQ8cGlqNVqgp79uVn2a/0GafCyTn3yN9tegBFmF59+LJRNis
VHLnXYmyvQ4M2G7cl9CzNxHDJVRzNz/1iDIWbZ4ZRjU9uy34nFNj1beam8mVCeixyWzB6Tq9TyUv
d7JNej7nr5k2quN+Fdct1aJ1FmZ+Xu4GUO31niK498rm33TdB7nGFzaS2YGyqikSc0+kqhuSuUA0
daQ9ZDGgKZOlxpGoya37fztaoFoU/4XhEk01+jospn7X33ObrPa4sQjhgHm8lXiAErQVC4E2X0Up
NLg+mYUTM3MEkLhBTraIE1e22RC3xBlMttgveqxOTnBObgAyKfIemZepuzCvOGwfqX3dWzj4+moE
GyTXrAYbPqiyhHn2djXDxuqVrovDC7zvCVPTG+fOpru+qZXaJZT9vXhjLQNSbX0WwkiePYMZfKgc
n2MfsgnbAgHdTdVtaQpTRnmJZ62JeijvroiJ5zHkIbcXCp2pYgEmmt0sOIv5qGFUoyPrpHfUK2wi
t22YHh2AKreHkU25c6zy2bx1jDB4Y+24oSR6b7iQMM4IHv4PIjpbCkm9FW+8S2GX1HpiuVQhYLHB
wjePC4q4OBcGXSPUt+wvKa4rnSVJCHQeZgKZ6Z81/pNl3YO83qpWcStucbTUKMPK9eMvSsaI7bI6
0zSkg0FA4a7XHaYRtir8JbJcvwY8pZuGW/UVV8s0KC8e7VxDEzSPUscdmA8ZPwyIRjGKZDyxs+MI
kQbAKmkrD2BK4jDSHEoN00OpJ3ATzHxrYPc8hk8hcRK1lb8rUrKi/LaObLcC9Oh5gIDksahHhKOD
knQzPRxCbkswilPbsNvjKa0VQk9f8lOmQr/WtZ3HtbbbNItgUZiJB7BiQxMy2lX8ztIJpo3p+z+v
JH7ZAxLDAiFdQiN2/dDTPIswswr+h2Xmg1875aiqL71uJJIrjTs+DpvxZN4GHiZaRn+Q6UWhm9Q1
KWZhtCSPPhlTi84k3JseOwsr3ri3jlj1RR7RSFnLl5g86lJWqkPa5FqXsoMmK2uTR9g/T1bwm1Sg
xkz2ME38UEIVZWP42doMBy8U7Y2Yr2g3BtGDdPmhbGxHysxb86CGps4hfFN9vq9IG+cHT4+m/FMu
C9cuxRQudMucKHLZKZOItavsIyyAWL3aizdGjBYaEJiuff/hkkQCqkp7o5EGqG7QDzjQLyLIoJie
yDiU8e6Kgq+L44ltfbOcr7zlx4KSf675j88bqT04z7zksN3Ytm1iCh1HCGEENc8VHSwTDgQkvvUb
XDYJ3vAMBB0tU9vawWya4FbmTIChqkK0pdPdVoAmSLzBf9LSAeO4Cd1bs4SY1uaJ38S04Wqrin7R
vC34ISZNNcN/gi+D3mzWTRQlJDn3gUOKD0g/DXJ9OCDyQLASpn4KiaI7UVIzou2vXENWDB7SwIc+
MkGaQoUPUUSBuB3iEJaMzDZRc8Ss0x4y0gYKrWESOK9FEwciNJ+5g1GNP0sbATUXcmhJl3dMaUzf
HsZEt6Q+R5S9+vCTdP1ea7+sj2et5EvniDFWPbqPR682xChZuE1u4sUhveQUFMkKmZg3PKyrKh6V
4UNFa99z7IZ6Pe2eUAdpp5jzT6jfr0fkSJETTGmr5HNPsl9coS4QsoqMu1NIJX52Sw6uKkY5k1LK
zECJm/0NN/PV2UcLr3Yo6JghlMx4E8JF/f7MirELmU5fYiBocTFfU+oaIBeijxj46y3W9Imjf5yO
skYdjEiFRR7cBjm34U1YgQMTPjTUcCJytNFO+Iqd2JO/t9diMf20cRHgHETxzeeW5IOqYrw2Jc19
CvfafOATRBdpcOcVlCn66KZia7y30bQjIhNTGgwSshNTaeJ5wtg7uJYQLy1kd57f8JwzNhgf7PDT
o3PRvNM29dugW54TSYaAWhmoeotRqFpygSC6ltHFJrJyiqF2k+tdumyVHVs6fCoWi11JD0XtbDjH
lpei1tTXQjkvNiGVen69fc6TZt5hmYtYlsZoAKE3JPFxFJ7stM+PghknVRoK1ZOA4hPux3eddo2T
Q/6PCVgrjhdyCQs32meDAf5gAs7EKySuVSyItP33E54cJRZfig9RdlCYvF+nOXoMxs7DtyOq9Pf1
lRBkd9qu+n0vhUamc/oGR8Lbrj6RmdTdnXzaktUZGF9DFsjT+//tjbk+LHdpuMdpHkmgCjC8hDjG
rspcZ3QLYV3rK0rNPfQs9/FJo9UyoTW8FiKoWzHknOVLI9Mxi73DUtugaMvxyUfBQtOMIy6xa8a0
PiAFa7K8YupsyqOvhvR4TthXPAWkf5lQyN9ryMgxlPGa4EBKAgqDPUM/8UrWjoO+I9agQ92shbT3
5rZ32XPVqbp0ysATEtPorylNRDECWS1cGMrOWtNmM97SqMLHcmDUzlfjrnlIP7HCWw4mLV1B7y4d
qOOJ83pJSiBvZsa5Gl1YK8KzVtQeh52IYeJMfLTLXIEelWcNEF6x+wa6BeE95JKyGtQXOtTTVC4Q
1dF5PdptjL5E6b4ZnDVOvVp9U0eUIEoLrJCOOTL3LZKuC2kIlHlxgmfeQ4M+fB0p7qy1ZIxAJOvx
gaO1BYtHkl6c3wUZjQFuOSmE603gRX6Vgx+rbUb21UPErg285uGI7+0bF5sCob0ccR2slWT9d6JB
9MC+zDB6ateeLvn1k3oOxJQ3XFaSyLm8LzHg1IOsVt6JTdFihwKph0GxaxUMiaWl1jZR1dVisZEc
FDZrhanjFYFrBjuTsNeQludHqlnPGD5Y3nP2e15nOtJiKd7E5zcH3ndPVXTij83Ytwd+4rqWTGtk
kGbK/I2cVSE9eHfA6n2cCUf5q8qyIAZCeVJSsmv9v7QHqR3s3Y3ftucVmshpCa0BnhGyD9whvGJw
08DGFMFWv8PiJVGGJ2MF04wWuxx3xla0v4pnadA04xdxxrOLhgaNypjhfqRBwIZLXq4cTR0I+Xfq
5r63fSQAtLMcIgJpTOeymi8cf8vwNjxxQbNgLD77WPfvMoyRpf/NiuocSlVrU40EoAggsqSFhNtv
ap2uLgelyCLrt7sxQwHWILiq412MFbymjgpuW4iVEBccg+qmJei1EkAIg+SYN4WoJHbYmmMdNS0s
4FD6C7YwLtak41KYDGS2nTr615usrklafeaAszQ7BGrUBNjU5Y+L0p9m1WSkLMDid5y4g7j2+vCK
5oKXqKA7Y7R3VopKTNmMyjvCbDnPdX8H0lf4I1q0GjCp7xpV+1qNCY5MB1XnxYY42RFnf2OcXk/h
XdHqT1woZzYgQcUbgYC/B3XZZ6sDgA66n3EGihmCmpV7VJDdDZ5QSHfrBTEd7eRJbv8ch+T2sBWT
iYft1dUro79EeYRSVTxD9c/ERmHhOFLVo0invgzSfGin87ZllDC4jQ7CtKVgITG1izoOfrNxSl3E
/xarXlsuoaU+CehzScVl+oGb5fPaanyjqV3NzjvkDEKV/vsxuG2Xe+CxHO4hV7w5m+iYNIhtRup6
W0tr7iXcWN5M/gGILlZN5c6WM+vXJFD/ZgmMu2210WD4wQPwaLzWqdnT53W96g6dKZ6ZOkUZi8pi
7ZOAKwg/O5on0yo9nSCYl5xni/dC7ERwbIM8aGM2c5bHjoldhMV5LBa48JcQplyFYX84b5NiHv3c
LQKDbTcUM3dY6ITScvsZf2xDt3G24gAspYmAUxJNNP3eNUjARoXBnFUXkkq9wjAyOMy5e/+o8pdK
UnyZ6VKo8P7JS2NwZJtMxu79YKRYN3L3K6Ls1+HOq7MtAB0YfmQZ2EByVCBC2xn32z86bkeQIKtz
WpEmd9VuAYOZB4JY/WQO3aj0Hwm3Fl8wAXuBZsfHLVIH4ax5uMmCzopPpPIkthW+N4MR5M8ZFjpl
WID+dD6jxxvT+g0f7Lq7pEfuQgspIeWyEGJebuAJQSL3cZBcAuog+PAzJWhxXI4xx0zFWvkTzkyZ
FLCAlzBgfmuMUKBU2oCn9gJgZhZlp3217smjPUsbwy/xw6hBM/CGxEYKynPVwWcScrWVnyjrEkTH
UoKT3UbetdfydOLqvFl73pAoSIi2NMKRBm8ELjX+HaJ3iEIaIm7PAV/HO+tRxBb/nxwSiVtqc0LV
kSRtsDZFmN8mPvPrbG05amN/p6MeBXM16R6ogg4w6JM6DMQ2agAY7ztbvn56EgZOcJJJpMVvy2Zc
afY8aVjD1gjr6mYyDZGtcqp96pyJvnWNH7/LKSyO/Hrzh417mjJnbdRmykZFRGTDXDe6binocHw3
O2X+9RULHt1lB3kvnWTZa1YcOX9H6z2njMrnAW9a5pdYcFj9NKXnOWWgD5m3NavFe5W7DLZoRYYJ
bBiKIXdvmgVhGe3mtNZVP89qkevte8gb0xRoYV7dLXjNikmqf0Vy/ecjgTQwTD6aoMD+w9BJ3Iga
OtXcRq96WUHKX3uwNs57X8XS9EAzEscf97k1aEDPe/Bxa1Uy+QBZWz8IFsUQu2nRo6LDimQqkGIx
pxRQQ7eLSZapGsCiJUqi32NXofYrXWsJpwa8ioKrnU6KZMqzAEB6Tl/Bojh144eSpcoRQYLczGvy
UXuNxM/hjSqjWwcy/BGxEhnFQ0yI/3NrA/nYrQ6/awGJZo3OAq59BJQNychOFjhLAnJdtWsVu85v
/GbCHaDWb9RrLpNjqKAqAyRPPyOJSeJAqMLeZSJEMNinInYAOZY7JMtyONKXr++INAhgRdW+020l
uUQe6PonvGqt6qyRskb9Q29+Q5JWLIE9e+nPdJl5NaXdJh26tUW8oJc8871an1m8X5FOyvBdprPU
3iKJEuXsoTE/YDjdRLF25jCkXVCZ+Fc9aLwwTi/qqZ3yCwdPMb3ZsnBs7F4FmPc0P9ZuHlwSxPoi
eImD0bDZiTQBYeo9/Gj0JgDoI3acB+TMIqtAruRkU++ms5iEyTNmB5VjKImh7+QeJpHtksiT6xIG
5k7zkRCaENPWgo+OM1G0nkAI2npLk95bpAhCt3FM+7K+aMyVkcaVgfa2pjGiPTuJhyfM3n4mXRbu
B1BcyGqEo65e9E9hXipe66il9IAaQ397oz2rtw3i4Z4gYYBNWNP5zl87qdX8yr3SRPOgPGQ4JMZs
3wXpg0X55+/r359Acdm2iFg2L0DmvHiGnLwieV3aClwIZ/Bohwd4JrRCjqjoW1xrAHx0o6lvhY6y
cJcc5KfLBz+C02BjCkvj7QYT8U4eFPP4i1wxEcogUrMf6zSoy4e4AUON+dzerkNJQ8Gi9/WhpW5N
CDR5d1is2T9Sz9tWynaB/SZyqL8AJsu3xsK1dSUx0WEqp6DL0z8nMPw5JPb7gAeeJSY91tqr8mi7
RxIGzIebg217A6p2jqiuzYcodk63Ofxyk+5yYfBLOr/auK9LAH3yrl1ah+Cl+1dC+jIjw7YhX7Vm
LsqRIWlKjLhJBiTlOfV0dlv/9FnXy9Twa9Ge+CDqIFMnvEdWovg1CUCon0HAGmRlAuhB1Cjt03Is
/DL59WEKoWCLwWOOATkTzm84WVTLat11GRpAS8i7ELFPZ5xkmVFiI7kyiHcXgwfu+b/0U7RiCaZP
ueJDVPLD31LDL2wn9kGhZuR1TTlamgYk318hpl0Fj07gMhVtO5yp9E3Xzynx3HsTUamHLiWPXqEp
n0Zf7FVYC9jshF7wrmU1/DV15oqgDMInNRG0uPmbmPfAVmVgNyZUYoxPFfH1YpILOnphcgffgUe/
ravaWsUtTojEC4G912GZy7Whf3G+8q5YjuDLFOPME/bl2xCCPZIaGsIfFvW56rF2kEzxRkGNv3LY
FydObxmHI5i+Eb3TKS0mmZ4PlKuduAmjTrpxKx7LPp1GyvIJBgnKCXUnYqxSiANYmOLFVQH892Wl
vPFYx7sngUc7ThXdr3ZIwTELuXRR45QXGgOJcq6MT0H9nf0420kFkvp7YfJlmXs04reA7OorL6rD
1LVHdwa++VbHcTeYGbwf4nDl/v7ZEL9sU1YAfqFdlLurjKAPaCkNFwzZJV/+VnP/z8IqsTePEUmG
gDl6Mhhpn13mv3X2akU2HGaZGVpnbCdAIIvV8Et+9mhUyE9C1bmmBt9FLmpufB0r+jYrZh8Y51Lf
ceKckdwagZWcyIPUcpWa2/a4oQpiK6FzlM1SQGisU/2S09IDxcNKf/uQCBb1iqFgTBbv4QVzZuxB
9kBQ5bQuaW93YlvozwMuXYQSfwu+au0vuXwQLp4GGMdwal7XvxpkNMQXgEc9jIXpuOQhc2beixmN
PSDACwb2+b+V7IeQ4gQVZZAZkGrs88G6uAApeX5c0coJuxx8TEdEOSG4ad+gXfjwWAnAtf6i/Eky
Z6KA5lS153100TYcZoOcSh5VmD5yzixLuJMHJWJxNDbSwtpWF08mPwSuoQEE5JOYi9fepYd6Fhaa
GsueOyqCiiyA32hIMKV8xA0wsFUgJHLCE2unjScsus1otQ8BF981IOt62AuBJZ7Yb99mlMdahOvh
CczvOp62wpg/Ir41mFedhE9AGnPdlRBXk7PWq2vp7kTo78vQIusFzx5d48iM8Mm+u88KHeGaA+WI
1QIyOmfw837M/NkhBXPl9Qcn2hEx6TmmKxF57odo77rqHWB3zMEm51jJQaIpkZYPz9qgGdgdeq5W
4y3HYdRASEvbnv68GNYBZjsnYJ3Sju+PXPc6b3jqzbz4h47VlZGohW62kHInAh9mVarhF6HRqDr/
36X9wDeWc/dkNSEXOQe/QoZ2bd7aWlnwwLXcv0xjpibworpY4TjA2HEoEvWdMEPZyeCv5nU5KNBk
JZMlBUIIVIqCS09HRapUCdhBhw8q7A/jeywMGOfiC2vdBeZJA67yhecy2A7jMvm59ZGIQG2LIQKw
H/GLsFQtRIWxpYp52GBZDbvLU97vYwd8IcEV4OhfaKpPsUsJ5BTaAxjUjko1BU6xK/NLUpwbktBy
6gON4LuXbsRzcRdyx6U7Rvr2beSelKzFVvIvq7ApsWRETIXFGMuYjGvYPqMAxzMhkJsAzTyx0ZPY
JJi4inm9tDEL5e1QztK+MWdV1fSGsIoh6+6NPOyTFuAf5+JHemcCzVVop4QcVoFf8vWjXu3pC0cP
rSzc0u3/BW50jKlOUNMmNUPOrveKV8mUD0n+gU27GEUT7NSk4Mdl9m2g8BJb/45O72riyWHxwVGp
Dy2zVaEfs0R+xLpMuoPIjNAO4Zqy1K0jYCaZAWXuVPwGmUxrGle0Te1oQxcqk5RyFvpCZyGWBhLV
Y7V9u0MAwJJiRAGpLSC+u2R8aFuurGHcJo9sPVb8m37trScZwEc+wW9Wg47UoxPhG8qfYkVsTtz/
AeuxFIw47yJ6gzyg3+bpK1iF26KRt0I7BMOwXOkwGSymGPWyUeND/UPVoiXsD83joHhQtr8s8Dgu
+bRP1EVEYTTDNU7foNBNYiVVmtGWm1HL92GF4+oinH6/Jh4/WTLwfV9VCMp+TOTkkDvVT8uJpKvf
NnHzrluiABRmDYWn9UczwReNTmvm9LgshOdLLj48BW8Tr6f4I5liEtIGo7rMeZ0sz6GZZb9mFNkH
0Kj+3YBCoSKAFgdsrE5v1YypwMoDHWRFXg9gnJncTrWD63NfAdpVw5Ln6CZfk8uO9L5ytIIsOFZ/
b4wR7WPnyljVQ8A1gjaqcijJ6/7/lhNZDl+UpHIo1X1hvQTulQ7C7JnUhyAJQKQtiPP7HxLioPz3
AfH2vPnB2uc7cofmAMIRZumUHeKTiLHGLyF9LwpMZ7zcwK2zMSm0Xg5N9KaYrCb97EmsHsaXdQZ3
5XB0fleKE/nNeIL4hFJ7lo8iaAU9WGqcy/g2fsdKSg2nYaDZWJO4x+WctwngwPF2CB1XFiFb0DEN
Fvrjx6lB89MBw1HRk56Pyj9hNc+5w6spyGs1QRQMUWhWNPh8C1qohA7meEf0jcnRDuoBux7UqtAR
NYg9ZbD2HuB+L4SA1FDoP5nMwr2YxKkSdRUIPl7D1zOxxVgpBhTNusXiOQwQ63jzuHRAZMsaEGIr
479URSnm+a+h/lBH6jOJmwVobz2ApUJEDTa98rOv2nEyYPuUvF7F6SrCA2wG6cPamV/1owyHZ5bE
y+SNkif503NxBN4pAI1n/CqrBnFvbfFBwgRInq0VslJPAHPlXHpnomqL1rmpyRBYPEwV/s4HqZau
hRQTvbK/zYerggWPjujPsU1Gy4Y3kzl9a9TptAG23X2BcVCF81sQLD1u8yErc46b8CAvaIEdqHx2
ukafpSY1hxwkDFGX7FoOauzVaBBJH41bjY99/cFB7eMB31XPPJxx3YKC8F/tS4JZJS1eRVQt5C/y
XW0H65hVqJoKbmuOfTf4s2N2FKr3UsLkscRFI9p8Tz3ZC0lDUi8PgemJJ/OFB9LHr115f2evHLhd
k/8jJI73mH72iXuMEJGNyPStDDlANg1eBl4NwDKWrX1tglmfmCfZaVCqkBD0KH8UF4dlAmxI3Zpg
fUsBis8o//Wyp3crIou1yItRfgl8CttsKfICOz+9fslS/pVduhyJ6St72maw62xaA6uUokDibxWd
Jf8uhMPLdINhiISVRWsCAkU/KSB0kiHg/lmCscLwuvT39dPP2YQh2CmPfiSy+I4nWKEEQaGwCKJu
b/O0Sz0Z+EYjghyRoWRRRoUIQDF/0EbM5L7wWeqOp6wbM56jN2fdmpfo/gxUnVf6K9qASvoOUmqb
8zAoD0Llewpx+CMkDWP7t/RbdKN6t3eVzlxPBqqRmhzmgB+MVb3hsNuFnqYUQDhBRl1+ihRqXllV
bi3EMZiGetVGEkdKe/ImFyNdEYtCvkdEOHpA5qMXl423QePgFT5iEgihjjFgDRy9FUKVcEFRiyFz
abzFYfy7HbkBUCmLcvejk2TKaDkeyYows+ZhcaEzsDfhlJvK6LBH5mYddbRJrSJ3ZtpF4G8a7Psv
dimTvzSP0U7mzmxsgXwh7MC75PB8Cx1tILI25UgDn2CovrNP3lplmMR1h0473PLrIg63CW3/2CkC
/xaU4NagrsaQgJXX/G1WwdK5F9Z+EnFPbIxiJGXiOKLuQN1DfK7mNeWmQONxBGoobS3LqLl0dzKp
/SoY3yOoSAndvWwXDfDQnX5bxbjOH6nE7DTFY/Xs6MIpcY8w4nJkIR86somRSZVnc0kmV8E9RqCe
ehI5nWdh10C+YctePSwqmfAnLj/DR+ae9OtkRoy+cLUEKtTfbqvkbslWn/uzV+3GK12O3ONRR7fC
hWy/EKm1UoYvfwPLpJpOR112sW3fpSka1RGhTcJ1twjVlufEaomqAH8vaGCdOcH68CM2wS9+Xrdi
mH0pMOUIy5rXGzWvSNDxv3oOyeCzGv1nJHOXI7CZgToekT6z91pWntUjlZwFOowKAjiAmZBhUGQB
p3KjMKk0lwi9V0qqYw08mpYTN3nTnTWvOSzn3cxNU4lKRc0PDsRXQx9hE50LhuY4Beo8SNPHC+1A
AfRD7c5aB46nbPLo5Twn5RMCAy3n5N8voFCCUKP10+2dQaipNWDiJysmHYOWCHYkD2Fiz+QAhDVo
1h2o6bww9MmhHm+CSogrpzbtMhmfpA/D5dq/Vet3fs735KeIMFvi0lvywfgXlPvvd9RX8ue3Hhpr
Rf0flY1b9U+UHWACkwWHCcnxt3Ls+rEjZ01z3zecOw68Ofk2j4+/bOhyNW17GAdNQX8uZl6MyGkN
+LHcDrsKPBbwrYDGcW9DwEOf6qqBMcxz/B5OTmHaJ1hgs4Qs1vb7oLGzcmdPIAmfPMIJup0mBpUd
cTUTbEMIxNDj7/nuiZNya2XQCMUy4YJHOkg2/ZMygDS1xsldNUbYiQaynR8iuVS7f0pkkABbunxk
gzNuezMA8ErplIytiu58xjjFVz6DxTYyNHM/Aaj7ozJHKyJqefyYKTFlZJWdF8G5T7jqWlBmTWph
3MuCtsXyGei79Rtv4hjk7a4BHmSnYsMn5bIdUuaQAu7s5gtUhdC3b62jGusDyG9ZYdHv4tY3/VaD
RH8mKUvgEmxELsmxjpB6ovWnNOpDSp13dGj0v7F7ii9P7o6dWHJR3SQ7o/cucTvjv8+xL5puwZo6
PhZAlIzP/eA9UtudFvIGIIuHLTkU5sO68XH6fP/85L7mvRfGHD5YWoFBHhcTDauEf9TEBOLizAL+
sJ5oKzisNEM8C3/I0XP/Haqwmo6AF91peUR+PRgJ6wrvtvBQY8mKBVwWJf5fm/O3qpKUfffn8WYB
Zydc0WBs8E4LpGWZ3n7+bIDIab9I/k4W00wpq0rDcHDPfYBlkKEEpRAyzN7VL9S/Jiish54u/7oM
m8wg7TOz2nukPeKl/FfNzZ1UzlEmMmjiSVKzF2g3de8u6x3UJHCxnOxJg0bidpmShl0Hh2KoEP4V
fnudZKwJ2DnMh++1AdBtwEtZr5jQ7b+sglKrBGYHovcW1HWKYOZMNjK24cmdl+nQl5npjp0awg5v
uLS+OQDQGj1g74U64iZDRcugSkfodZitV7FnBgVnBnzyBEI0erFiCIc5pSykKsWEQE7WEdlTYdRL
LcT25HP3rwRg5X1VUd0BfTOVA502auFK7iPyg4yyU/SPwHGQAxsU8E7R3plZmXtUR3IIt3Hsd1uw
U15gzGHYaGessSQ/rSbDzTcjt6g0wHcFFimTuhqYO/VEdRf9+vZI/ucdbSz0uumt79p9GPVSez/m
pOgsKdF2WvyEDBf3x5RP0sKgfp0JNZnfjOw0WuRnCzmQgtqW/wW569aUH6yxmiswdzZniyKZPDR9
M26nH6zn0PYJtRoS9sptR0bHgfB6jvUV+EvJcGG5+icFXqy3NMxYsqBdjP8RxOkQ7xwj38t7SCY1
T+Xpd41EnkvAcsi42j54QroKL5MR2pEck7zs4SysalYPLkQVhxA/zjIRIVmOCPUMZf9iurAMwCja
EKxBqnHwwrJCJModAR3ZziGd5RHb6J6Qe8CrHgj3srSoj/ulR1ptZQCD2nSspzAhBBlFIaSHPCYn
mfvPsBdPn1lTeSyxmY/6n7c/4f/Yx+OeG60tlty/frAH8dwvAu45stGZCazrTfVJmDlsEIL3CL2B
s09rrr7bBFV/gVzgNky0xPwuvCk8CekVDR9pXk6lzm4vMctdn4Z2Ln3ra9TZ/uZGPDPlu0TL6+S4
rnCVrlEyRSf0RdiKmxQHpq7ddJbUvW7zAEfaDdpmP5B4pBY2sKNtPnnhAX4Xz0tt9c0JqNy5jssw
IMIgAcDO50Fdp7nRAXsuJ17wDKtqrHMGTB+XohRvsDuqhrltDame7+pzfcioTACIVAUdmbJsfpYB
ZLKBygDvGzux51n29Ik2BGDvAjo6znMdcGalFg1MgEGHmFNIi9nE2Qkaqkn9GZsOWEEk+0agVPx+
UI7T7iFKHdS/QLWfsZmoQ1SbKNk0duw/prga/ucaVO5dJTf3IWo51fhzCpp5x9FtMW3oYWyvy6ab
Mw4GGIIXeilGduG49eGD6SvkjXF0pa0WQERRgGBnj2fG8bYhijTKTUJ34eH7rWNTxF1L6u/YQJEH
3IFGIxYshMNT0rfwjX1U01kbMQ+dSA8xa6igwjq+ySMqi4ht3CgOXaR/vzJmeBaSLtubZzUiGLB2
KyPvJ388tHDqXsAGmjmQxhLDlylMu28t575lTfIzNPnPG+FyYRdGKqQm6tOwgQR6rbonLmurY09O
7klbMraCtXhY6dZ2tCPRoYeb582ykXXvIbVvl8A76Br6w80wqnoFQQ0q3+Qj2iGCgKnmK16IunVS
pcp/ESRAHpC8h0RtqbKWd3BlkaUUl0GhoZFCVsGglrNyMs3iV2qXqPiLvQ/cDiD1bAhtm7L9g8sX
fjrVH0yFN8n7OuKxGaVwmWia9TfI5bMfnpKsny7MG5JTOH3L+HD72e/FMeHIcIakEyl9W+POVdSL
betqsFKKaVFd4HND91/pdEMYPDEHXYOns1pTn0LdymJugRBLOyo5fnxL5SU1Xit25xwphNfcsGB0
wyC+g/dVhEFSV9buReD71gP5GZYY0hVSPcyY+e/8TBfefCljjyD0CF1ZINY/1n2/n2iAMzUmN9CV
UbP4KoZdoVfaX/os5lyphbC/gdbIEKb29Zv2G7GQ56VouDi6cGtF6ui2CkTLGZhBlgFo/mqSI57v
pIVdGttbndGqGA7ivOEj33jZWFpr6rn8wNCB8/K1+xmesoBj5Q6Tx8nDccXsTXMaI32AR/Xp50WU
yiTMpGU7kxnIUq9rAAVet3N3ZzXOa7vfqVD0RaQABM5HlZFpj1M2UftQ+owylQhfUCf2+aN47ovL
Lbt3tBwNhsnHncRXs9pnl4HIBKu4gsVcGUEOqqXRvy4IXPxdc4aBJbO1xiGAkRHwpneKdXu6lSto
yUYTm7wPTn3Cq/mSmM1kp4ZwMqG2moYf/6h3YQcnWH9raNorlQ20AXZAEt6pVN3bkkG76SaBy+e7
1OLHDVQWM47Pj1VXBkE9RoWstAMRNC+NGZVU9kcIGvLTxJ5CA9mkJ8JYGkMYc57HuFPFhqz8exnu
Qq0RwheS82Ogtp/4PcuPlx3lNoN0nvOZp1V5iw9uGFA4jJveZBLcP/xhDlOJ+nKHt6OHPByjUGqj
RH3padtLH9fXlTBmrMWnivKny/Db8+ug8XbRzEXTJzZjmbbhWUTotEVRUpyTxCKXSbDcvw6LHwaH
l8Y46Fpi+VBoCFCHK8fJn/M5ec2buYvXvt11ShWkyDa/aBQjLbtzq+5JjbSicAVflMAE4zVg7bSp
hl5Ed1o+nIT2uUHXJ4l4kHm6ZsNElrKjL381L7wY7xuXeUQAfeuuaqw4M6Ic9ahF6H2wTzCL8mZb
E3oe7zdWPbKItUKLsbk123eTgsTzXbrkzM06cV8SpvWbf6kNp1Qp/LvXskiLwUurHM/xloDpfS+K
uICeH5ybZgYXVOg5oEN2svRp5jCPTTmW6MM12s1KmRvB6Z9fyRGAZx+SRnQB488kGE+IlQHcktMQ
c8mW2yKJqCLLmTMYzbMEOvaq0toka6XnOP4aHGWICN/eFzaKoKJUuO/pO58V/0SAr/IcSJ2/MW69
VMUb1C5EDB4o4Sgp0nN5ifiQHxINfWqRYB1Ma2s+mhE5nHIB+5eeC8lICsY4pEZb6vlTpkaqxbZM
ta9oxSoXuGTvuaOZ68kXck09v7pG+jZE3IXGqjznq0rvUHEvX98muEEqNcJ++0WCKVttc/KhB6uC
9GrQJyclB+BzVu+oMUyo5O3SkRnbmLXmas1cyKH165bAu8z5WwIt4ByuXvDmkUKS2n8AJBRa32zw
zmWzzh5X2jDkJI8FFj+h3allTL7m7mrkxQGZ2LVusmWLfokR3XG4p4yzXxnll0dSw5II7vNALK2z
t3ewxfTXO/6ovOMPxoWiJscsO91lp44Lf1HN+RuJvja3tfnLu4XDvVc8l2hstX1yXM8pghDU449J
hukhc6iuf8JA/ascc+iZcXbDFMd4OXbYyO9VJtrENYcmNF5J974kOYSPCo1haAfFLXjy7dasrgVC
Th/LeLB0kV3uKq8VdCqia2proUBZiYuK2p3OQPcgbcjNrS0xADF2OHD/bXqmgOUkWd+BS2d9IVEg
Mcn3uweEY9srDT8cbuE3VVGFhn9tXnj61degJDw2ZDTjWYkHwh9otQGz3TeawxmbHZyF0sVxXSxr
KenCl39gz/FLamGHkqltpAPh4fWMRoFHB3PkS6P0CUGUBBjSTurpZ9MDsdFzvHDv54QzBSgE0D6t
LU8pouWLCYXHnxOw8dKSooJCfRES/ER71E0ZN1nJWDT7AHEtifjkHHcBsF45HzdfcDOO/laB3jnm
LnHC40ku3j6X58VVA9rJnO4mA44bkI15f8r9nCnGHyGo/lmv1LzRt7UYogsF+KHW7dKes5ll/ptQ
l2BzTS4Bg+jcmlaxnX3dUXYleoRxQHcTBhb77WrHNwn5eoAZC7JXsrfs+L8ySOgQJvr/AI3zY+2e
PPy0HSk9t2gT4MweazmdzsaKCL5OGfm6aXClqSyThW6kgLLn2nuYo1Y08rktJYIlQ0sLTdTXEVt4
TESbNn87LBYhTKNg3keSMfpLeyy3btxXcAuR41px68/wQNVMVbWchnhUoz/u/eSWi4ArIx8T7rUN
YDf07KAkeMERdA2QnCzRYgIS13aBQKpbsh2ePnaBoc/keHcw1QyDOZhu64yhMRyq/aAwU9dGaFrp
1s6B7d4KS0tgoCy1WjFnKSzjR0/VWQjHzpLAKYdiooR7JK3t8w4VHA6hS7u5HlKAutkGN3oKBcj6
hhnJtaPu0mm7Si+MjB991LMqPxm5mEm079csGrOYA6VtRzps+itKqGTABZWrNQ8YtK9W8kBb5ZMp
b+IJhFhjCEpfZGSDrLbV7FIiJZ8Jn798CeZ90/2W1Ts1UrhY+l5nGFXa2cxCMX08hlNDOeOWJzkc
Xuq06Try+OMcw4JP8LlgX9dLlVyvJNvKYw7jMONVY8zL3O6aNz7pwKj9n9Ds242v6NezU6egRlZw
5J2L09HAn12RcX8ltCXQItS3lcXIXqAFTkw+qtpljvIEVvktParKxwYc3kZExCkHbrlLJ46OniKw
5XD8zzI0YxgKEeITGdUmr56MVM7mRgiNgf+NpHXxPRvg5OJPfnHYhyhpDFSG1HpmWHDkdZUOzoab
g4s5PUoeBr0RobrJBNBeWmtsKBfiDl35I9R7HE+5yQljZLpC9B4xehgog6DM2DzVfvruRHY5pOid
NMggi5DZrRRg9OTU0TIcwEAPY5BJgZA8oxMTBSqzBPa8jBFRrlm9ZyDqDPedEayYlZaU9DWaNsVL
qbv+DPJYLdRbgeNpGK0ZGiurg+4YZL1GHnHAyvj8/3xj9Huj8gkBJ7v2Eo3gn6W6YomiWAEL3sac
jW2xQVeD4LIEwyyQzmT+Bp16cvN+rOsnCIG1VnMoaa3vLRNfFn0GfGTKZ2WhVGUel4Nl/Xd9SFbw
M/gN3RtOblTgPp34bD8TsA5QjkrPak3yGiZngkjxOfL9j+VnSJwAttt396R4TMhqbA59ZD9zm9jx
36ox5YegaCLaabR/CywR1xbSwa6EbRnsgs+bKEFV5sTO9h8ff/zHu9AizgenCncYpNJ7z5s4tUwV
kAGn0NSpf12x00R98bGgM2+MlTRfIyeTSHDbRUGrvjG4IGrEQLR49XKX/a5lNvX4I5QK/kb/bN+a
BWhUQLA6cIM4B/Fbetg505NInz+7+KjV1LHFSnerrWjCI5sDCIR3seaAXquZoVinjzgFDehH8MNi
F23iYae2FxQUMJacnNiFBQpk6+FLBAtewfeUsD/opy0jI6yKf+qNgXceCOD7L/A84peVCI9yNPTg
2F5QO21optflTWkYClRdOuJO9wBdkUZzU+ejhbDUrsBnKL/DdJnxIwEtmCpx5m+hDwARxc3YGxwk
Cd6Bwh0tN2wUCq6U3xILsgMk9+ry5zaz2fa9J9KUhKxG2/8z7IaDdXHApmy3BOAwcB59ZndkgYK4
cDNNoTo2CHxgYUrrtThKyEAAr7f9try8jc3+c4229I8rW5jKgqEUvC55YKnSHCkwg+3rtYaGOA0Z
GicHRSA1doJbPKs2Z4BRGbjQJKwZR9BzcW9axHyWJ1iv08/CnagVYILu2DEVwUbUtEpCAUSF9+d8
qr8AQw52f6XZqPphr/dKUT2ESExXx5Hccx8MPfuIkMFMAXFpEMYNT3uxmIAVC7iyUunnixXhfKKh
WZyLfoWO/vqHbJeNvYoMM+HLvcjJAyBf9nl8nqXpK3jlFsHmYgUzHCQA3EeaHs5cu4oKyZQCpWXm
RPOwTnmETicNv4phh2Uj9kEBQPwCNtUxGVEq2pFC1kfWx25VgsWWPYzOKdlP2eCRZn1RZYRvv9wk
LbW8RfRNZw4fu/KJjsRrgaGDG5qHeEgCcSsTY9T6Re7sb30C4+1eK06s/jfSBc7ElVvm0AXsfzFT
fxv+io25lPHXmAfKQiOFawW2ZrRyQEYheo4B0NtGgED7t8ktn+IX182D2vlFCzp02Uel/D/MTlki
10wlBvpZLqD9n5WVJp/gahbSe5/rSLmdjvM0TY3pynGThNMtAYSkszaK1HVOMIRfX8e+3B9jy0DG
qeODtIyPfb1fMiCrEAhvtqNv+KgGtkmxwmFMBGGc/XhXJjv9LrtAAelqjpqpPrFA/2VJLH2GHsjr
+3pESDLBxqhNIUZTrfhhiS6upjE/B+DqV+y+QXqatY+LcbBgUP1g9o+xwYVwUgdU3eSvzSafdbWc
cQmLYSxojW44M48vKJsvnDjP1P5fqS+eZApdsAOlIJH+4tMneDlbV5WgE9+cozMxnTfOE3D/SOA3
Pt/zlBfTjTrZV6omgMBURmVPkCTzAId19LxasZ4unDXwly1jTXCmKyrXNjHgtDJ9c1PQ5yXjv1BB
DHKEeF1uJyGRL0vrmCSRMH5sSradfH+zX3E/4TUVJ/EB9sUsvRQq1ygfLHxGayxtntVTkjBBaPYp
9pGSy7TtIrM2ZOBHaR51Sxr+gINZM0zrYCABi7Hu2cGuRDYSzMKxnEOKYP4PWF4xPWIHRwwru/ta
DMbNonMc4mPjC6QdKvsSO75RePVMVX2cvogoolmU3ciSo7JnN/ABzYBxzvu+ggAzO8WyarD5WMCM
NgpARpQKEglJQOeeX1LSx4WBja2eoRDd9eFhq0fotHzb14zEypahVoCSARKRh3d24VgGzRAtQQBr
rydB7Bg5kMJtDFd20Mfpuko3YDGezTNmit0GBugbunXbd3VFedzgsU+Qgw7QNA9Jouzfz2Rc7y8P
OM4JUwx9bMVfLKOFMIhWm30k+H5ly4OuAFbS7cZA6leqGGprAGrSbOdIzzRLAZw2xce7cxG3Rgse
FpBSF0AHxyfvt34MG45pDdIpmZthoDNU3BTNairuQMVjpADBp0TGSgTBuXr3l5ZfEgl3KMA2yznX
1zinwGpFD7qh9L1yerZUGqXDCEJckigseCpDCZZVx2mBI/sAO02gUOEwWWgQz0T4J5PgCUnYKdHP
sT8+z+vsSBiBEwoKmb6dXTOhNFOTtHy1jkjWy8Hkojo0M5hMLaWulMd6nvfL1lYzWDJRITA1T1i5
6+h3NdSbIU30+weJJpHitqG47Na71QJJ4WWsUE21ngSW0OikwieEfz32f439YOawLGWjCTU43HIj
e9U9hJgTJWKegg+eaR+TBuA9LbS+w6tkmb2+frkx0OqOg2zerqiRV/fINJ2Q+fkuU36q3BJShtG+
d0CmkEcFrXl8HHhPalZx2xEMwlm0iabQvlauc8il2Svk12jw0+vtO3oocfO7uP3H+XOOQ+rQOKZI
Wq58cksh8CXGUJ2vdbi7reRQIj9qV+ATEZpsnR3QaJnjGctHm8GkoxyIvqlhteUILIvUlJ30SlL2
tMt7Sw9pl6N0gbRlt3gJWHiwAciflfYR3W5KA0zkFba9leIqdsTBkSYTuzjfmFezr+PC7Yrs7uTN
VKFVik5Xlm/QpnZX3jGrBq4RAJykh04ZYbNIaogmFtktjVMGJVzPmCAkAq60AjgZm+M+UfnZfrT1
G3gHkswDcGj40c+bHcS0gcoy6gA3wHA9/eHncXZscPbuMzEFMP9gQMyE9nSI+33DlcmwwKWroDiZ
zlT7CE6nVGkUapj9Syq1rh9XeubV6ts8AeSEQtAEl95AmcOus6c297V5Em6lq1RLQUu7I/zp6tF0
bq2FLH+WxFp48srJ0KVIyrJZP0te4RHHReCPS+cO9XkDQeKC4yHdVBGbQ0tHdfKTFuhBkfRIK216
G29sKD8S34iQtEuh7npUeVRhcK5IxtvCbnYN9p4C3YU9XMUG9D2TyL2/7LIvFEmL5swx4o5+mfM8
gRRIlMUYV9J30qwl0u/ZnL6+/3C/xQ3qOSmGoojz9tmo7673V5vM6hWGycpIVTgaFs3LdvrEnW+5
hZy7ItkdXXBR4wO7GqTtWamL8d+PQ4NNXBpQ+Yi+B/0TNY6FY01JH6NCztvMjX2yVPL7oSjYjPWn
/Bc5gJ1ZcvZEuCWa91uH/7HwOn+8uFc110Nvk/jvpMtxtotujkrm8fayG5l5IexrTWqRwAzC0Wh9
SuQiRyCqSJW+0rsWtTp2hCbV4z7OGxiBvX7Z9QLHG0+pFqGObmxW8LQl/zyqdTbQa4HlBHyeNCrm
NwtkyXRcBkhJNvb5HM9mPCxHc6I+N5PGEOc+A+n2Txz1Xa/4Z2ETXLdkgOak8AM+0mO/aLeyd/cK
23VXaW+6D+dVM62C4iIVhoQYNDV2Dou4WN0zrc3sVYnzAg25XK61SQ8KPHlJvU7K19FL+Q5GpS3B
/LfnYs5azWYbwypywvbD48K5m/xPsMB139GF0Wy12noYxsCUsuxmBp5AD9qfVLsllamuwVa3ldul
gaqWsfCqVccUTybLCRtc/1xQADVDrCdJ7abvnqkg8onmjwQijjXxX2dHa0QiDZqqImTD5LWeI6LM
fUZKPEXq9WWJKSEwhilWJ1lKC/y3Dj4n/kACZ5xAZ0FJHyIZH7xDXQmvzj1vnA/vCnKWrt0GVcs4
+Q1V/FGLERDvHNfI/5dWsYVMIDpkRGHXMrGQw8NUQ7k/wbrufvy9UnL35zjJ4BV1Dy0bTkOtRuY5
l+XeBaYg0YdsbpVkErWZhCUqVR9NvHg5oWnYB33pOn7nY5tZ8DonE3WN3NoyOm6U5GBC0e02V0C0
G9E5ozTrq7JBAq33SQSlAAwW7qhi8pbiWMDByNXAYcm7mOCqoNYxcqQZwxYY8zlGi4dlPMkuR0DJ
76PdZOW4yrW/ksKQ24DNDsVwD68Xl3Pf1nlZIl/WLo2NZSL3N6Dbudp686yrHA9cJUAoWJnWKywS
eIY6E7/0I2hqf6yDAPbg1GnVcHI4knp7VSjhAuN3JfYrylvG+UTa/rZecJhqZVXyq0XFuxisJxrK
PQK46vC7+uyljdtG+hHWvD8GyUdP7uqya/9I+oh8IyzQjkmjx2dv0EpsuxbE+VG7O8xQcrJVX7h6
sNGut1bbQDOddsqPBawTgdgeGEAzrqSMv1W5fkP+GuqMs7m3E7rIE6px3ZfSgLRFAG8LyOsjQCbD
/20uMCPaTJAbUVCegY6KiBez2F+ULPWZIB58PrrwtxGSLx2MO2SYxqnRVNGywJAgiVa8+gVHOvCa
6f/0rTBP1L4jZxMvkdrZw+oX8KdZvxXV1dX/2t1ktEsIT0X+BuVTTnbMQGZABP9dUEWeXFBJIjf3
jZu0jMqwonyq7rcTCMcB5x8HEVlx9BVAsPw5yu8a/afH9xL5ouwxD2kw8/jkqcIEN3XYKc8GxZrd
L0FRpDC14+KLycejMrwfKwBL+xfihxzjEkD7yrdAiYP1UF6X64JOJGljodzPj4aoYD02u4k7lCOH
SrXXEdinsugYaUuHBXawpirJGLeY/XCLXVkXmBsD9gC5gKAG7HDGM/e4fdtvkQDNVqshdoCXJjW0
VVjw5fYZV1QVKXPHYChL1b5bN6VMCf/ny7Ee4bu8qjavrfui3oxYg4eMWZy240QptdMii8euNtW0
GAYMRFoMdI7PhroD+R7O7z0dTNecqfIQZP+W1Lo4PXc5t0j+FwluGk2yao+Nb2RKrSrCzwETqhmB
CIDLazIMj0NXjsY6PcsVY/50wLFOYbXrxguTTGhWdTPtGqIW3V8WmxHH4osz6tWQ8FwUzP4sY2nA
HjsHuDT+Wzx6RwJ2eA0rgA50U797skFP/PITkObGR4BWFDTsgUwaysIUc3doTXav1Wezkj2DfRJY
Hn+vD6FC1q3PL/9gsbGkhftn+npky6R9ldxEKpUHsMWUOPQrwOsVWFG4BTGs15wLnQpC9t8A9YbL
5RKnx0AnqRPjH7LHgLklOwgVU7ibq4xEDdHf98AsXg7px3TxWfiogN5k6aZIzfSIt4ynv3VgSBTd
Gt3YVteMVQBqM2AKB9KRsbZr1Mf4O4qG8SXVGBiXLRNEpf1Nrc54keHeLVpTCpdyrvu2Z4O/Ek6i
wPHvDqy4RPdvJU2DJXVGqniTiJXwpyxhLBLKPNX9aOH+HUbmUu/SmO4mwabVizI2idwcIhtMgYUI
8Z+njNvDQ/VAfqFNw4FJLuz4jGh3MdyooGDX9Ck97BEMfRYnzdoZDX3yHpf/aoQsZjT2/81B7R9g
YMC3CaHx6POoxW2sg57r7fRJ3wwfrHUHbHGav2/P4U8K5ttRhQwj898Y+TwqAvEIiIJUn4pX45rA
6kpZlsjNGSpEYPysnyBatLrDJxsiT4hkYgRCKXB/93G/h2+6t0AE7Ubg1Dq7ZOb2LhWeCmjL8jJk
VCr1afcsAk24x8uKBVlBkTaTsklHs0wavkUXtCGMOIBToLxniMYTky+zT9BHzbIbx7MzOJGlPeDp
AuOGMcOSY1pbkvS9lTJP8UQvVGKfWD1XL5Tpu1LEDFAdHB1HBtO7lVG/eWvQlsg6uL3qPbGPVnAW
WOXz8swgMD8FmiLXXS1QFi/NIQW2yqe+sCJopOapKIHlpD8ctG6ET36ZTmsv7mhlQ0CTCJYDaj+2
ks/PZ6Km06uU3FMahfeO4QGCKDuWgKfXN68FWbx/rG+X+4uoMS9V1sk+0I8Ixrjfl9pXDE/BQNbO
pXanSmzxpvj5Jcj9XNeYaHak3Ktp6WAJ3q5sm0Y+mdg3PtVIXzip0INLwkuaOb8xfaypJWMoKeME
K7v4f1mnT5Wm9f0VV8/HkfcDM6HjL0UN5nN6u1jt92nDufUPSS8y1dfpswYhqx5aSDW6DadQ+Trs
USy5p3ut9YkPmhVki1P5/Oi1OgNe6dYsN/iJOqYGJ/3pRszGNUd401WRzL5ZqbTTRs6XsruTh5Re
OXQ+tKhhp8CGO04FRxNy2hUmdl23f1TJP+p/vbPKgkAC9raQn9mo07a/9fq8l73iOBskm5v5ZJ4x
29nze0c3tHYnJejFra8N8gZV8Dx3PfMbozwY03phcekeALxnYT1PPW+D+JfSUXmTZhyKB6SJKk29
QI5tLuMrD14xbXIjWOdUwxn5xPwi5rLcObjOSpYxeEVgMHtZIekCp+tfAsP+iZShG5vFpeTbLU0p
bjLdDC5agwL3HCqPGAun6Ug+EGhovOW07oo25DBpHPGlsbUBMEaMNVO8ebuKTTesO7YB5CzcO2x0
n2XOV1mvcl0lraDRlnmsGqeWmWGcfkOvuFP/QO6HB1+u+MhbTpm5kRN8nfP8MweT9UljTiRH7ucn
TFZEXYfbTsN7V9U2pBenBWgx2+6lIJ/j1LS2fSvTdJM7TZGnTnnY1H5zrjJtSftLGwnRpK74mhOq
chbAiDYy0Qbz59XxvP0rjvwlQqdUreAIgqjR4XQC/ZOCAtbx55WYqcibnQHf4bv0APnINWsoaqQH
hpWwebYoswdIm/wIuxU1Y6b3nDIibTImFRc8gYd6rSC/uXHBFxzi2qC6Y3di2r20KXm46WAcPSZK
99Z2lKypYQUXWxHN1O3ERprk+KoYGd3kv99waShR0tQrQHVII8EnOWmrUfQVJPJK6mbuR38kD3dv
f3Iz0xIiyKiiDjyS+VHmtdYkPeHZE37XHb14H7Vx6V1dgveZdSV1ggT764ikpq02XO+boQVctBNc
U+F3iFp6ukN8YyJRxAkN5+Gs5isfPIJH+9SLo9JJboqh1/0yiiUtxnhCiOkVXOuSl/CshQSTBqYo
th+98hICpUzYRhY3AWF0HQyNwnf1GIlBC6KVjc2Oc/F+2OqXyYPvVw0OkbGnF4DMJmRyXUSYd7sB
lovACEfyaVeYp7a3Ud/RfE8TI0faNZIUZCWFIQigGapbMUXInDCYXkPr1h9wBV9D7tZk5JgMpm09
qqOSKo/T/Drjhp+ptdJypzH+mVryhtAucdWw3j2BvNzebtYsUReYVbYiEsz2ScVZivDVbzQ3OlnG
OMQRhZ+BYFeqQIFJKgq4usdfAROonfvb9XOGiaSrBkpWqLFl5GmSFZ9U7VKbeEfRtqpUDyuUHFWL
zNwN1YMqURI8T3iGcQWoxc7uYEVzksts1BqmEtjvFLku15LeIqpueY9iAWD1ftdHq5wSzL2LYyAH
xxosRflDnBS9q49rFN8gJtmtqn5gWkjFitFzFgx/HgLDMzabgSou60ReHXqa32k2iyFqngdPXyl1
NRn8BR0dwT87wuIY3MSZgehFQ1wwnxYCdMeTmrFU8PZDLime8X2q1XMvIxeR2TtV/L85t3PUODsF
fkKkm2sj+DjT+4Xh6Iun18FxfGYpjtVA1smIJszYncn4hzt9r1H2u7CMGgmmUpfoOIClrlOqq/oP
gOQNbsizrJbF1LpE5JQRCWCCr/QuZrAyqwVCurlKMIsFPnYOwnZCdQ07huhUQV21xROV8BhwjdlF
TJXWOAE8aZsuevFW29byxunovJXtU+T1rkv/eBUqcDiMFI35+ZWdK4qCdrZfU3znlUTpKS4ZUPOl
Ab0/sjWySsgQb1jNx081zkiyxEcqfSafBuNkN3UpE5EaxqdP4iwjqJNdZTZ0BHm6zpfHXR29oCj5
mxlYYZGagYNJo6j+2oCfXR9IcHeswLAJnxTr6Bk2UxU++pGdAKYpsfJL4nQG0qBiTa4oHoxfeZs0
scwI+9i7U2j/FmGztgQ8TCqkFWElxXMev+WWCGTCwppu/YxhMSIFgsEPFvs8B8i8VDysJR6gYvDt
3RYEWd0H0hT36v5slIsZan/GD3Gu6m131H29+agvnmdk9w8ahn33gGElqAwMe12GwD2Ie4iMrVPa
3EZiGyBDzCsSswJo4cS1GQjxKi2nSD6pWCq7YxCsF0VfIzRT9sAR9t2I9ZkBqeGUciiNkGuLEpqB
TTJGamQS+lJN8BqapT55z0VjCR0C8VU1aMe4mQ5wvxqyJiWghLyG0iedUJB8xy6jKyb3IYU5dqks
zXpAER62x8TlL7gZVqZ8fp+lQNLxJ+EzRC5VAgSOowMhW4guC/6kBMb75l7Bl6+NPa3ZQnnFfOX9
CtkqPSFmDyGjBW2G5cLThNHdLxsuYPky+zpSjgHHsLa8OJWrIF3bCMg2BIGnSHfibtah/iMa5crk
WnMHGGUJGVXBwFsQDW0nFzAUc4K6nnhrqWUFMI45w5FAC/ZxWjrgjyUCCazSqzK2vNW9/TPLXddb
kbEZJiGJj7/zWmNT+Sd2FIMF1VOFEz5nAz03glCT1PznRxgl4024XFMFVOBHQFT7JpNvFELsgxuI
3m2QznPTgwZmkRZkvXLsvXHqCeNfDyPST7AUZJjXLQx1FV3XKi9N3G0fDyNOyJzcykkxHv8/H21u
+yTx1P7Gsfk1xek8OUJmSKkfZJY+zX0/vCiFyf3b1/NIX1DPiMlib89RqCtjbra4z0KRHtRZs9OG
3IL3haSW8cB75+RmKXVe5Lo7LfQENVa9cwLV+P7AI2JaeuCrb7EG85MJpFhWnnMXiUbas/5mo/fP
iK+l4lHPq++IjztKpuyMZjEmEC0ROKefsIOv7D+PC+5avBVlGFIE75jdCgSb3JYaJ23Tf8NGfX62
cYKbIDx3Of1MjnHxFRi1RZdWUoqKW/U9CS9kmBuolORGkQaiISGrf5BjlXzW0CoE6zCeZtxU8z14
YfwAKC7e7RwWAVSI8eq87yuTRhMspuW/Q3wpG9YH9NMaOqM7Slz8w9/1mjR8b1ndQncxUQ2ZLb5h
oKnOKDUZS6oxoGon8fYtOM1fu0+KJUkdl90sOykmcNBjEgtgPKlbvdjUY9vY1TDtk4c2FHRZS/M5
tPWy2dynRM3/kGzxYYKPTDVYaFG9hzx/dyCTqo0PyIywXDneeVugiQOPrPqTvO4jYxh8sJDxMioE
bYjaeRHgnhyvxmSoAwMM+u3Uh2VQxlR4+jskIu9QJCQyPxUrdJjRw33/wdUn4PGF3YRtaCMWdYOj
FTfX8KAecqhWJVpZgATS2s3Rqigj8K0phyOFc2Rtm+UUXR43rM7UgG/kcoK9F7GRxBMGEgxxLB9Z
87LWf/jS772DVrt/yD4Wc2UF5mDPszC5HBSs9br24Zbxa+LxJt2YsAfoz6cuYjkVdH08pdo2JuDk
aw3K+jr6WHx6cSOp3lIdcXGO/Ion3YL6s4lsXjMkI2ZiU7x9EWVDl5Jj5VA7slnafFHuXCr6EmE8
fzXLH3zFxFrlaPluU2FmpKuoWnNFOswKyZklH/ki8hKfNEL2/ePdFuKAxX4qy7i8Bqomi+VObKbJ
rBalmOQsrLz3ZSs1Ji76iV5SNQWYSi8DyT1RdQx7+ct/4WruenMQK5NKotsFJCXyKqeMMOQtrZ6F
4LoVSN2Dq7/IYxireYwXn/cwLO2VkkBjFD1KcqV+co7DD/f9+xBeOmNMCdOgtytEohKchNF9HGZ0
pLbHWFeALeG+qSr3WIvyuAg884Fs7C4TZMvUUgwFWgIUuj3LG1GR7PvrxGsXQeBpkwJ/QqZhM3lf
RFkdX05sNsXlDR0/juEAdnkSmED80eisiGfVuj3MQssZ9xcv74WYzPctVQ0ctjAGns1Ls9krMBji
8PqJOY/mmVryXziHrfz3zaqOljndv26DgyeHu+EID/MmcX8i0Re/1/4YOfkdLE8sM+ZJ41xyry4L
LtkHm951kyT5vRSSTYIo5w/Yov5vwzpoZEj8qfeRQTB3tjzBwhxc6MTRCCdfyb2kJIJNpvmdz0uU
Lh82p3wT9zC223+2pvFp/dI5owOX4+B4UZZxq3EGqysHXRE2MNq5Z32c5Crjr4AV/Qn9fBMXveMp
HjIbu378Z4dBnAbQcrM8nvSxr9HUgJFXR6XbAgUruOZvH3+YOKkaxsQwBrNCONBxhStIV1gY7dUZ
5Gps0e1qBbKpTmFNg/ijSv8lVZMQzdgAiG/57ABMVcKyl+LPavlGhPRU2/8070rhQDrVBt3q0yIm
kbYvK5mbIxv3YpAWLdWOUKJu7vETgi/lNy5DiOek0KjOG1bwZc4SFe7CKSbLZnR1Azhttt2MEjbU
RGsDoybLDcQ8PESCLsib6Ys2/tZPpJtBnI+QBRmbetM8rt0nt9LqHezltoOKmgt4JjO8lSb5xljL
hr+s4TNlURKy7rPTPPpm6I8tYs6x51ByfTzylD5CUrJ1c0OAHZ+d6Zl3Fbi7Z+GaEK/4UqNVr0rV
8ZppUx8QNPkLCe76oPy7un74cjjR84B3igEH5kMbhs7pM8Uf1SGkIywZiembUUJvIw83GXW0pydU
dsikU+VUWEZtd9/0O2RxDwrPKXEKPCXJvi+WiTWCthk1kEmnPXeZqCLoWuDRpyihbncLT24riwYi
JRRMW/jsVtoo6VjJvzbokYeoumzhQUDOze+EHe6rgUfkNGz7Ixmfh/+/Xm13sfp4fyz+HXa8vYBj
uBYQ1TYOHXlIL2/8GtnGTa2ob7fw8w+W/XGxiKXi1legM8PYXE1bW1xTcFOKMW7rp1ZR0PVHkDbg
ufIN3Hc0TtqbPfLKiKbXeiUgqTPBcUwpmp52q0S8qYo9EgdER6HUP3vVNCv2Dl5e6ZGqHlvByRHt
o3GvbFpV2xW35kk1+1XAQFUdZA7dpH71fveRRf7ov7xEb3SmqWndGGhGJfG7JjPoBcxjv65zqnk7
iq1rpzdBTkE7d8KloxTI9TjJkOeuwgTTU9yxIfrzvjoItMOHMbJQD69Qtyzl7MOkv+QiO0XmlOS1
JjkrEmTTrzaOB+GjojPukX0PJU8WUiX4j2jhbr8sT/2hYWl+qNTJt20GtIG/A96c1Q4BM867DY/g
6DlkXkmv57rM1bMnWV6Wycj7rxWfSTHegv+G3c8yfMmRjOySFMuq5+pxMaycnsOmRMtKpTFBCe9P
ph6pELRT+GgtKq8LBjTBSf0xIrV+Xsb3kFGHv3vKs/KrESVjJQvnq2U4hDVrAxOzS/tsJ9P+R/Sj
pIlZsvQ3QDwyNSsMbp8ekJdK9ytWXgojD272XmETe/uJtEqezDQyt5pm3clQ5ceoAbXi1gl59YkL
4VCeS/drI5VwpblnPUkOyE2w3uipP2FVDi0mGPuaeEIQfCtK4ElyYvf77OPaRePe+8ncdQN1lTxy
d8q2VxQOlPklOjUxB7NntFtyRn1sYNKInO0q+YLkQVam/jc3YoD/heIjMSHmRe//B+liT5o/FgzM
KemCw1GnCr2VXdN4t84nVef0OuCuIVGssnH5bDqxxk4HQvMevR20Do9xcaErByb6DCVMIG9nL+O2
zIhb4GjUc8/kUjSElYJbwWYq7AybAs6Uny7fWxrUKH745XZuxWu+gGBR2O2bVj7OycCJy+yZ6Vay
Bh5OmzZruj3xUhQT4gpF2ULwqpRGrjfgPwFtVLiMng2HNhJexQEAZijWr5SfVceWUyWyyjdczO3Q
F4rzWpvwmATgrQTgODPZkVcVWC91hAWxF8e4LIz/XaDQ567RfAEW4dIHZxq+hxZ6QCSANQs991SW
NtOqYwDCPEk/W66c6tj7CXWeGiWTeE/JBuCv4EK5xWWdq3WvgyWHsl2Xf4/vt3roCIaasRQ8VxoJ
KR0srIbC3rhuiZL9VQNc2P2GPzi9AL4pD6rhD7rXE1dI0C7//yrTXNAuAbJ0MM0mswY2uE4YBaen
HBNoE7RDv2LgAa2lVaxhh84tVT4kRQtSw0p92Taje5KHejKx2qw+vcnvPRisKctE+OrgkQz6wv3V
oBl/RUQpk1OLlhnQp73xlpHvrpKGVUYvlkd2JQ+SUrbb3+Nc0UQE/VVxx6ukDPKkUjCHp/EerwZ2
vUAVLHnzj2YFkZnFi/2RGQOIhgram2H+oCzpsiTh+CuI1Fqt0NOpZibTiGPZI5WljmiHuxGKjDsI
RyTxh3ndyoT21IT2XL+5tp5kvNCSiwcaf2VkkeyTEc9KThpgfnN8Owf+8FTCWdnh5JwcVi2LP9Pg
V7onQ7/e6Ro3irfBCZd8xv/IMUR+m94vWVnTUAw2/6mC+Wv0KMRcWhsT/oYalrQ8i8ZxwxIpB4Bs
QbeeuQdA3cKkmn45mbxhqap4Zv96RcY1WtlxjIc5WhciOoDxuruqhprYQawfgpvxy22uPPjlSHK0
qW0TEa3RxbVFZ6VnY/MjcQXdIl4QV03NYm4ztrxH/h7wZL8oljNKVahYe2BUYzkx+dBAk8/K7pIm
/IVUpaLLnuzCQ5hZ9gSzh0LBdwuSWeTJTfJPunTbb5fGwCbHuCaaYcKKpar7BkDeYQJGLIobfyCc
X35OKr5OdG5IiKOEiqTgHCWHs+n9yHQW3DhDjU/DALZUSDM1Gjqrj5MN58cl7ugcXGUmhs88mgYC
k1u+6dQ0u3y/avlexrBm8pSgOZLP6MVcrccdwrFJ/9+a8cth9s92WXWUknClH3HNYDWUhoe/51Wx
/A3iLzzFk8Tas3mxjoLBKBjgm78YOhN0NbM+sbz6zMKMYri+SWIjdA+tL2PNzSkA1Bsn021opF8J
aOC39Lis6ShT6taXkGtu/Ov4iKvLlRV8A49RTSOPvrAvb4lW4JaZiwu6QTjVoDlbkL8IniC+eqQa
p7JuXjPOxfDcB/dZsmfqFc3yBcHXic/VicsKsf2WqE3gRvSYUuWhTpSOH9XIPCgqFpa1Mtv7/bFh
+6lSNQ4NCHG1Jw5DmsrQBQmDDQGrehIC0Ih1L2dVRFF+hMg08xfcfYXkmcAQHFGCl2tN+SG9ZDhi
q/Ussy7HU7jDEnq0enD+dBLG1wgcEJBRZK5eI32cvvKmFvFH2VXDV6wBuGpQbz3hJsCTSGi6B1K1
6ewz9SSqtRMEV43OJN1CCNLeJ+bkTyD1o1EiY6mNHiK+Dadk3VTJDGoFfGF2KrJcBUtaz8y/2UNZ
l5LjPp0n0QnlzH08w71t+scfQuTqNUpFKOy6O5qRW/fTEzbxXHvUoidHS9g6HOFJlDgxIoU4U1EX
Cpzj7+iScSrKJfbLWoNEyDcjrCCF3htQ7Bjpz9vFxW78BwD1AeoOj3Y5H5rNmYi+kn8u32Dyi5mM
hnfwKdvZoayWk6MzgA0tXy8MVenJEWcI5QNZWzGKwB/6Xn0Bd08Yacv7qF5QnsvZvgMGBlghlkfJ
zX9jZJgJTwnJ5VlcWyxbZAkMyHf3IgFjOKcvIl/DdS5nuWeEEwjVIQ7SY61/BCD99zXEJzw8s9n2
Ckgs/rZC1kfvaHYAvDUKk9CW9ER3tR1YjUvNvFkyXVCW4uAkSTIvDf3oclWR3yw5w6Tdnv/f7Zzt
TZnEgWKP2gTvJhzDQRGGh8f1AOLRfT3nOuRfuFuQ24x/dgrA13plx4tr2Y84g2Rgqy38/wIPPW/s
MSV7ykGgwqo5MgHCq33ZWyfc1AXf4AkYt5swXxUreNMcCsPxB4/lrN6KppvKK719pQYx/qNv3Wag
gQnHtIMdd0q7uHZMudHbQEPox0i9Rx11qFclI7fhRggIDDA84Bdip0FiUYQx/+PQwXBkRPIi+bZy
luJ5CFoVpeeb4FnvY5pNFc0hRkyjKyC+9vwpNU9dboT/KI6Go6cC4DlorJ6lrPSIQfZtoMvr0yB6
QE/xk/jpfv7nUCXCfN/ng4qaQL2dnm9DnoBY4iLcgaV99LvZimhb4SQE4lZbCGtg11L3CDjXdq/m
3nmM2Q0EvE4n39vbEeRpVjhpb057v0Dl9xS2KtwTQLqCBZhqPfnKfLaGUzSQjzhdt1gHJEaYBXCp
gCHjJBsbTHdpl6o8AtaxR6O2+nH7HsiFmB2+7aW3CALo0JnqBksZZ+9Vts1/aBboBT5eLKYusNv0
msMRKbfl2h+Yvf8XQH/1yQE5h8+CifkzFdIPV+maxZVEuwT04wkF86dYOOJMMWmX68Tpn3S6jcUo
a5MYdodKmSSnB31+B+tEkJnf6gK0WElLDi8HkTttu40An9YREFN0tnun8qDts1umYsxML9RBzLqZ
HxTujnbNcb4ln0DgNRE0FBY0Jctoxf0gOf5JXi9D2l6lImTDznl0wUAEW8zeFQ/lOs9BOF2PpR9s
DA2nIeQb0S7miYkHC8ioNlqHVVuug4d7lXD9cnUMQFni1U+7WBz88dAg/siP0LgV8kT7iclkyQdN
a3hunzXQE0DKDqmL6di+HiK3MqUoD5OF9KDWhowz9Ntypq6JW7ZX34b/7qktGUFsDXdHFzvvpTud
33t2AwuVYIqAf2PZa0WUaCps+KAxtdC659QESIqia84rXLFTeBohXMy8oUVn3mzy/8JaOrxtyYtp
RlSn5c7dp+zXKCVzYyeL8Xb0gMK96i5o0BQdr5EX2/rTn3gy3W56k4njFNHv4GwhjoF5PA415Bt0
OH1r4me8TtpW9SytjceWVXW+KpmG2YwpB0YbShYOOgkyXRzOGacUUHwsYiKgTarS0k7IKD9ma68i
YCijV12/k6HkMSO8TnJg0ANr+EhI4HdzjvmGXDi7RK10QngpwQHpzcW3tPFOzPoWbWcGoxsNsy4E
YKxcKKHrA06TFMgx4yqDJhI10CGoco/8UXMYYUAADrOP23JogHZ+1y5qxuD0q515k5Q3ma7604wU
Kr2izkW4ATvIQIkZXdLuoDxwdeskPXl9KBYWo9GN78iVDx0ti27EA7r5NYgmnn0TTh44mMvGi397
oJOBGziaRN8fKJnHtqIMwVXuxSYrY4bwzZ6yrMSxlCTsCkOUMJV2KX0e3O4a10q0cfqUBdSCai5u
oz8DFVQku6qed7HegV0gkhzvV0EWp0Ym4bv//Tevl2qW88domFuoNoAd7K6kRc4+DGJQlScuqp5Z
ZaWAwZKAZwCqvbBEcBnLe1+IaqrhI3TOEIFKV1MfuI9p4DLyusPiyLlBfXY03vfOGq2dNHi9Mmrc
HqFaY21KSb34XSr7J+HsBaH6b/oneUoojJdeL6AB7msVFXny6vvl7p6zTksiqJExRXiTYHCCwxrA
fIb1X4Z7/GuFqkIu9cigJjfGs1WXvsnfrvOTU6vaWyw0LTs41hk163iP/e5InINHWnJU94+xOqih
eJKMg2xEUm9Oypb9QTUxWV7R2JwMbLEJbdeHRHcau08m02c63a6EJ5yI1SL0wn2DWN9oDlG7kCjL
2tIk52oIGAd0mEEWn2bGYIb2OQYF7ZpggwJazJQZryqsWa+Zwge9xCD+f+jM9YR5VUQwbM9d/fNn
v0+d5XuKghyeAnPM0bgnr/YEW/qlpWmlrSZsvAC1Mj6izP6j2V8cYp5/EBOgyF334/O7svDxMNnm
dsCTGPMr6LXf1Gz9jdQual+l5XpzOxGSjnM3mAx+1/MnMr6m5VC/FarsyxhjVs6DRHsXPzL5H4KD
i6QXGgBn6JuQnzB3uT8QqJKaqUEhbbyjIjuCGhfnFen6TOwKZH4kEOYuq5k+fq3kxBflSC2SrgW6
0v6dOnQEifVgjVnsDd+ekC7WFgBbBEB+rXBc0s2IQKhKxALRqyZp1oHuBGw5P2fGoBdY+tbFON0L
WhGXnxmQe+rMBZA2J6Kc2UN66E6jzrr9pxl9Qu56+CCW44XX0/S+2Enak2fEkN4i/utzFTWo+4Rs
Vx3h47iorMuCBPztEQ2rbfVkqQY7Vc4X9Lvaobaza7nbfQYkhe0nNdyF+00KW61u2QKJbpnq5jes
T0uNA3Qvr13B2/AAanHlr27tcO+scxtcMVAqsduIMfakQNHpAmJqnP8FKMXNFVgfrZQMDcS5ZCx8
4VKTgL+Pr4kvBsStH4vKRyAFdsYD3KNso4XVDfhr4DoTS+55WJhvFVdQ7gRDXM1xCkOfCoOZ7BMJ
inp8/V1WJnjemJ60g7rRRyuvO+smPbZVBHSjumiS15i9Glz/0esDFa+sShYiajnq8Utyn/s/r/GG
C4tKxzYDWWZ096EcpxR8f/2BirnK/eyIwcQ4jqwNqzd9rzbiJ6QpEwR/y7hw6NH6WSzxhr/zradK
hhIj6DvGVoRNpwFP4MuaJxMYAimGYJ/Rv9ppDUQyvbH0WnGHPCx0XC/uIDR/QZhWniMYcpq3L6kF
UazLAWjBOjyT7HYfJE8rZGuMStZifCUBoGBt4N8sevJR/l3Oa4qtysR26Mqws9MPWbYH78cF3YzH
Bzdccniaoyg4ixZtAdo6udr30A/TxK+y39sCJP89UCv4FC5toa892g0v1ZbYGocg5roXuDemRWD8
hqHKv+tIDSjjrsTikklo/XaXcIuM7oHYE+1PfqQUl+tjHUOo+7nsCSgx2BfXRCgkYGAdQr/pUkcj
UdFqc8ydYlgQhhFdmv5dx6eGC6zY8CtdrXSljywxVDMgM2JbMtABedIn/6P3KUe0CHnKfFADBUka
47bcOHhwHijZxTBBC6Rh7BC/kzAztBcfTVX4Xw+TiEYlQNrkZoaDQ42th8BgPZReWZ0VyZ0EBjUd
RNyufk4vBND0nHMMzWvzrseMSOFWZLZ8V6ccxbK2ICtGPwav7O/uAtXX8wpTzsx6OllzxiwQxIkW
Qm8JoL6Ov5iVYUuMBG+Cz4ZDbL3Wa1ibsSGXduJWlg6cCpA5MYLdLuVkxakkKvqcz+JjT2jX5BM/
2u5oGuBpkWH6+Sx07ol9PHlxLSO+0KPgdwhuwaU/409HEYdsVN1YvvoK7M7S/7hyqiTvvxnrL3Dy
Q/i2R73in2yZ7V3x0YSznSRlzvMFfFY3uQfkW0m+xqFGhHHb1YVlOBCeI1Vyvue0b8sVF+tUk6kt
T6sJuUw4HozyBPZJrjQ87B25/btzD05fveiu0fSdybbgUDHy39BCokxExQpMf66dAl1HBhGXpJHz
H++17dHXA9Xat1N8RGCQTRWGesQvCtTbOkuMD57FhFAjieN4udTy/Og0gg3YppUn70RUeDx1Qi78
wTVPOXDkF9Zh/9oXkgRcZf+zK/GiCHnYgST+6htecjHSvqKUA4FNudWu3R5sxI6ZPEdIiq+a8/aR
3QKj9BP+kQldhaNSax99YWG8ewNe8i8mpRoqVyejrZk8plaEXcULf9xHwAQ/CVmeknNEUd/4KgPm
FTIWysHbzO6yUfsGi3CcGgonEPngCtljB5W1fiSNKMf3w6RWuaUxjp6LoI3HJ5g+TDzRMS51s5OE
TW3dYnpUYztIMZ7+DLikD8tCCydIF+o+w/QHlGmzQOG/xO448BZdANpnFbItjhRzQkwwSx5lpctg
+m6W7XSrsFwVL3JlZwzUSOUAJUoycd1kJq0abmRDrw3b7p7srhbABplxf+ljVG/BwlhcgUzRkLwG
pOWfKYaDgVaP7Ni4VAPuM3V1p3Qa6Txbf2qEGQGl4FxFKkDSvRAYI5GOQ+vMLiHJa3F6KRZv0DzL
2ndfTv/S+6AncEk7LJjmyU2dkgdnj5iToHWyGQstv2rL8gZKcbucaiMlYD/dwhOYffw9HSH2rMub
RTLrK0YUk/Ns7Wj0rRQauGS3J6U/bYj292JvJ4XRi/gMVhhZHf0AUtoCE8/mkS7eM/yMDVbJYsrg
CDI0Pm8/tVBUTaBzEnnL2W2CNwWvODGyzkRbIFfgNB38pxg6ZzyaDgFqHWUm6NUfgH4WWzaDEqva
sbcLnnepkSVfpfuoETY5mm/VOdDPIGuA8YZjzyh2R82zGZC5bOU3ue+I1NqbpBm/vr2poG2Wrhlu
A0ltA3ADNnfYdbvcicRVy5XFMMHVDPRPxmgvSCqSLblPCYGZCvYzcG+UKiPMqf6hiFJ2bkpz8/LG
qYuWyC+eg/wO9XhuNCjw6aIRKregLmMb6NIpJy7tNiy+LZzfRXdh9Iy98LTU11hHBi+dZqXOgZgg
mSqJo/hDqWoeBmvJ3p8jUwt49qml8AogUqe0L+cvVw2o6HE4uEcJWwRmmEwFQtTVrVD2N6LaXkmK
uAfD/tiZUl7DaCyX5dVca4eiRYpbw85yQB9doyWc9KhrrEE8FN6HQdaGbqTXcnKoqRaMIW64Pb1D
42gRMhQfWnPq3UufGfGS8Dgam/ErZJwlO4S/6iKRjVPkhjq+QntxFPqOP0PYw9OcRVWpUh0avlyc
ygL/BpAGuoqc6OiGABT54u2j3ue3vtDRQbGxhNpOpErRJtZY+kX+yj3QJWq7H3gz8BiptFEuldZ3
pFjAoAWdTakMkFF2AxrsiV9r5l2A6LhmmCnCGt1G4w6L4TtVFmhO5WhriPjWLblo9ecIZvAQsUtO
078zJxgOwSxtZL4whPwtFrzLh9uzhn6nz2wqG6a05kF7FjE3zAsZvWLH6zW6wrzuD9aGi4nC+mHW
ryXJwOKATUzoac6PxREKBgqar++RdhU/ndJjfAHcHGCnCoCtBTytPTkkpg/8KoFGlb2yHyKnHN8k
7m33lbexB7iULmGAAZ0kMKbTHEBh/Zk59PYC+FgaAFIrgOLQlRpazUmGh/G3IggYTLhlNqEFksZ+
3zx1HzuNKM52rkcukUF1K+82EuMTVPL7jMwJ/fF2wQSj2AXPuNmvunvdZet21i4urTu1Y0S2PTq7
od/T54m+L+Bg1CgEdEs3nNCHvgARYPj4pvza2SWAmWpIoTTRpih0gQYKGKQmTsEmteKbBhSlF5xX
kG61M23QU0sW89VfQNNMwVBSpJWyhQOBxCxVMmiAS37f2ywRLXI6u3gtnd+p0RYDdBngeTQypwjG
6kF/k8LRKREKv6pXLeYHS/ydv6LrGc1VF0xycK5teauwIKKNE/Mjh2DakSloSPWA5WVF9RRlCr77
2RVvlu26YiL2J7Ih2PGqV13TjGzeRgnXSCmLryXJqCxDsU9VHX34Aau029ypRudJupwM7TdW6m9V
Y5YFMXnUUjKEgnJeHG/XImA5JwIP8ZXcMQ4bH7RGk2uNADguvXYl6/CX32kEx7NVH73bBjE7jrmf
YcEamfArDUn+g2dl2x3ykrTrNSGp5hzNW8tm6d1ONPaCAAM/jxLLl9DvnbHBXYRq9laVmjIrEliH
8lXoKmleLtIijEKC8wCwXgSwJd1ZOFjIZIafOeGLTP6Kx4vble5zW5cPf6emOAQ8yqELhX2Cw3RZ
lKdIGDLY1Nngtg01Ua/fCrks03S7EFg4Z0DWn2Qm2hlb5ZEoZs5KB8YR6056Ou0PcF6HruJpeJtU
eTFzUK3xOHiP05PARokBigsZfyVLXnWAyiWg4wxqmbwUYlvA/nk9owouMG6YzoMVxJHYB06AQ1AK
hntmqcbbgIpicWu2clfqsE0xdkuLinFP3iHVMSnRelTZh6H1hdUwJ/JWD1gsB8r2YAIXHNHaacO3
gN1xABaaZEMVu539NXoYkYTzcjE/vB3WNNRwvskPApUEC0Z3fKnUFWJ/SI3RTRwhGQTqwT1zcII7
hbsvEcnwWrFNbU1Mv8zmfBx6bd7rTm6WhHUWG27orw6ZOXhmkesUmFXhN1vS26Icgx6HPz5IrIpk
L6Pg3B+dE0D3uKquV2ynQ4Dr9gPc5PKqxIW1hZUqyQ9ngB/yAaotW/Um5TDrmqCr080JmezBCXUn
nA2YbNocxoWIGh9TAlQEsgONsA/KykSug0SV+lb4nGaMnSMrFNr3tebhrOAqtAgaOyabxREKpFXb
ng5u4CkfZSjpMx+erg9PGGtTvzOOudqLPqrJ6B5EpTf90OPnXNyWczAjFUIi5wLBwHCKLCO5KNg1
x8zmCrZU60k8YWwM9dDqSBwBgwr06riiNWrh6AVvtFYikke+iKCH2svZH9Xdb0zSdyCY/kufugrO
EHzRhw97wQZTeV8pkPIJAgZy8aZpnaafPF2JerafQSAvU24nvH5/kYCn+QACn0xgf7c9yYUd3vtk
PR5rhOuyUDO5qf8pk8MtLEAOXyYwNhsfQPPeadNtUnOGr8QnTQ+F6XyKmfQk8VhIEe+Rq9Muuc88
I//WRWeA0onEws3bx4J29heYlvuU3Z/N2t7kVqFaBqgeEnE7lU7hCHAt09TN69VhEs+l5P6oPH8b
u36S4FG9DKnDbE3sPermUUC7++DklCmk1QJa5h0J3UA4U5oyH5LVxCkxFk9JY9EV4e64XygLHBsB
fD61gUFYeC5tWEmVvMzVcBTCWPM5xwtHBSHD2LcYDPpwqb2bY+15OHOeDc6KTtqA4k+LnQCyO44V
Hgwi9ecCZ2xep3a4k7W5XIqqfsI7AGZa6g9u4tQcDsVHzRHeIt8BhMFA1HD+BxwCbnNs8iJYmN+k
rXNiKP7TAw6Xr8qTzO0m02lkRyeycfmgX69zYIXSEYx293osbQvfWnRLqt6Fk34LSG9yUoorPWJB
V2CgmVzFkmqXzexSvi05N21Yjl9c+RMWFUQ2r+NU0gdp80jiSNriv5ypRHYbo7f1thqVWPWj7Bou
TkYRMdb1BtzSQdZlVi5W+Gm4IoPwl6301pXsyAxnjNb43aq+LwP0oyMDynOjqAIpwuJu/rc98Fhq
jiAEV6McTrau4Q9qW+QB74gu0gzbir+laM8OS4zHcE5GdrFG5Wq5sxAeyB/AkwIiwCHVji4GlZ/u
HMHhlSiLKaQH34vU+yNqJBHs7FV4LljyfIsZUxBuP5hX5GjrxU/o1LABraayDPfXJLciCll7EfR6
poyl1Z0KITeTJ1w/OvwMPNY5bv9/c4NL15TMqytRHgHH1ehNvajxc+77dtqPi3CEp0R7CE+WH2P+
YXVYmg3t7BHqlvWjj4j0H3BRcspr3zenvno1V/6pQkYQyWLl2AgtN1A1SQi0QQBuxUYRsANrTL2R
a6nhTtvBVoqePhK2xky8mUO8g3Rt6fWtfzfwTUqSf3744Fm3wIC46qGSZzZ1lHrg50ZF3k4gBA0U
skuE72HOU9SDpyl5fJ+np6f9ripKqJHTBk378MUivgC9v4Qr1A+Y268zf6TnhwVg9V+TJ1yssZi1
9ifwC2NLfLDGO/JFVe/TXgYQfsp/+tFXcM7GD88YToDjYqJgJ29fYed+jXhRsYPrEZ7VAsq5tGXl
Ow8eNrnVZ3LTlhWBtiU/zjmxplmoCDXBw3tHOT3PSGeRk3mKnC08gOcJmOhIdmHA38TSZUntn91p
kXjiZeg9+Cj1sgoegzc9ZBY2mahG8fDf8/3f+U72y+ZyEV3yaOCOpQqatJmdTgQYfLsbs9Uo7P0Y
X8UDyP3XfjIn+4Gf029+WjZdEcsYFFGvb5Hk3pexggXTglvdVxl5AoyMu9oUopOarc4l3LXiD+fC
lX7uV0l7gtoJY7ZzoqheUIi7bGLhgtYUwy+TfsxMQEhl44o1FCgzFHGvJ8DwEAVcNm3FrswWtvZg
f/Kfbf6jkDYzpyyiZmJFD7w6E2/5TqyY/CVYOUVPoFJZBqMDdknfl4UOv2x0mG88VrnkhDxz5EJj
ajGJNdHJ4vrjXEtDdRNMS+qhI0qJ0hLCVVGU7q+rWD1J5fUqG2pVVSUx5n8Agq2OnJXFFx90Mw59
foFD0N9IhjCDfpJOixmM7og32h3vkHyYY1X9SiJ+4YwTUxJkUQWYd5X5NvvGEMGY0xnUnfiVuTGP
Q6H3714M/b1np4G5R2wmhJx31vDsf3bRypG8lXU0O5yR5tzOunfH4NjgWuA0HvwvbExd9egE4ahG
1sCnYKgaZmQ6TwqFdOZMn8Cy1XoCeVFY0g+GQp8iFAz//+5t6jYD7w29XDyElFs4Xw70VdTCbDb0
6crQLo8tdfPpBnYuTZRflo1nTzkQPDZMsqDAQevJe9qKgHmGfcl+DEmEBxnHcc0CcTMTNaZdbrZ8
BSs+UqKSOpX7qt2XyFzMkdgpErZoFGSHu69mWcVcU2FBI9hyjqEIpJ8OHMknoY3HtB5cELo2YbTm
SOhQ4rlPM3KtquFrGUEXvFP46tze2TJOBVbaa0tPmXRpiayN9gO8l1dtN5YVGh87WTICIrVSVZ63
4wMRJiXEA5yq1Gv0/8+sx+N6kjrPdLpq58uzAaXdzsroKlhUlQexZD8xqL+E4WBBr6bstW0FKrES
WFncAGRF0TfLiWlY9sfmI8ouHFfAerG4noI6raWxsDPBRBlssV3zFs0eP5guE1hSkDDvXuaLdd7r
0F3zG5Erqse439G1tUKe/9gPd4G5ux89X5eadvAY66qWoxI49K25Pr17NIAiCg6cgpfj5Ro0XAjT
eMgzBPSVFmTK2F2jyUUtX2ae4swoTBlBiG1ihHNnijAzXP9Mc0lRuhZ00iE5yrZrNX9AAtfpv1vV
DFOM9/HORBUbAkLlQkK33UPWncQNUIvAzMDeIqNgQfQq5O/0LL/DQM6B3/Yeeobiq7Zu99mOYYYi
tdscT94eul9lGV3ZqotuIegCZIjiwmjY3gzMqhJZjLOV5LcwOO2D3SD0LbM6x94uLsW6CDvwyeKP
HZFA+CpywXctYtEfcqyUCzpN1SvElBxEi7fqS2TF6j9rD2m7BCaGltoLkKvloyAxKXcQuvAN+rB8
qsE+HVoRLZB7OrQ9Yr/dj7D4QirQclm7AyZJ3bkPx/6OP/U04DLcku9X5ycW1V6e4+DWxB6oxKAd
r3+Ghbuv3YGbsoPF512QYRrjkxkARdjPSrP6e2yVVecubf2Cn7imrvd6lXYoE9KTTXaqQviMDayp
2U+Gp+37TIyEwFGGrgbK3rAeOEe0iQSR8ZQGgOwke1YpMF2hUYnJycA34ttUGKcr29NilIUR24p0
gmUSWSZ1uEMcElKmhXy1Jx1oH7fal9IqTbhwEq9sgk/vufm3+IV4DYUkI3eWxESFnOb2xAIAELoo
PhNkRpZ95czgLfzEMWIu8/GU1K2yLeGp9he1sjXtcQOJ2HDa+1r3DgjwXQQcIECjhlc6oefZMfak
Za1NXdPu3K1K+x8h2lrhk7DvjcccmygfvhGOWvwKbdkKr+U8rhIiHTeUbPeJgEoDEWXkyuJjotuE
XHnTduixl0j4UVhQOFNpBWKOC3OaZ+CwndYEYXSFZs3PwRxGLZ5JlCtqc3UTOdCwcivwLErIBTQq
hHbUceF/3tn9/CFvzq2ePpgcFLuelcXhttvbnAdZsJRe+AXZzWcUbE+tk9PzG/5E/Vv113Xt3eA7
agKWhVRPpFr1T3rVkP/iWa/hErXT49/3DXiDFB5f8c14BavCX7WQwXaY8L9tZhb7ez/+BHfAmhND
36xMHgy8ZHGbOhtVazk6bqAf0QvISbqPr7ZZsvDvqsNMcCTtILJ9UgJBWyYcr7Dwc0W7NGjUjqIW
+ng6c+LMM0tN8kOWTkEN7qyw18xOiWKW720z0TwKu5tJ+UGPBfH2+YZ83nuG0yaUOTqiqnP7y3C4
yA+cGjbnJcs5KN6cs8mhy7bM2PzJ0kV+At+ID4TlTfzrPubvWHTiqg0F4w5b+u/mXCiGYWnl+upy
bdElVg4TpsNYWy3M3DkATfWFZS3qReFsg1pqBtFslKCifUmm430/cHvvr23sYA0Ozkod5YsDJNYO
L4d1nKn6zheoBXteld48f8ML9cw81DlawU4eG73JqQ4uR7WPM1vvo7nCrITqNtJRouBFuJyTKNQd
KnHtwCR1hkJnHewDYWHD5Vcdv/xnhmClnhZSKDWHSAbzHmWC21vRt7MKV2AaKg1VHgbOKeaN7Ej1
kJ7mrQHekI933kKxNauApHcW+7k47tragf8G6o0+iyPn4ZvA0F+KLiCX9UTNijRyGWp+QfvqERzr
bPwXSaHDSGeZBhWkMqFrlyxUsJ8fwtFH/wx6JgI+/Bx50LwBnKmhAypgkJUCSQvPGuLkUFM51/eU
BdZNwYpwdI1xsBPBjHYLT8AQXKyhjHXQaT6bQ1whTXi1AUapLxBVhLCEIt2s8bo7v39cA7HBbAxZ
JSTvxEbHFHOkQnCY+h35j0S8UGVtRboY/yPPjE89t7SU14DbOLr6OEscyP0SAWUG5G7AGLcA5PM3
mqp3XgbA3xSq+OjGV29Yn/WL0JIR0jGVhpal+muZP32hf9XQrUaCpyxw0JCsdDGwfQ6/psnKm1I4
7EVsvdNzO8GHZm9TSRGAsnLV6hsuR5u9Ekyq+bEckk7wI8PAr0SWBr0E9yLz9IbMJce5q9j0MH9D
6HVcFxKrG7NPwq5wkcOQMp6kGmhXSLAL0gnW67audJAb6oqcrOdwQuB9qvH8NmcDdUNCGXD+PW+w
Xo0FS6FCoBxVZD7Uaop+K04dw1ezp1xtCyhsMf/c2WRG3h4SpoHHc3gGOKPUzqMexMmFuVw1kO1M
2/JJersQed1S1beU8Nk4F5V2kxCZPgou6Wc9+eUmkTv0ssLy6zstQi7sBcqNhRlDmKEB+TGgXI/c
N89oiDGvjE2OHZXwdYxi31E+KstYGMpnpTJCYj7Yo1YK5fn6p/21VU7tcAsn15WU3H4kGvUKadWa
Fmfdjh1VyKDXf3GjxZ3hZRlnOS94VqeRgMiyn2SbWmBuhDIoxkbbBpC3zjAsKcYX4s2ck2+JkJAb
y/owH1rCxLaiu8mJzimWaXKcGDOeU+Y0ogoUP8iKWDY4nmnGY6UbIy0sTDIG0fOwBUSUueVwxxkO
HPCz9Gt0cG2gL25of6+QeZMKUNXJFp87vLJf2bLW0qg5UW1w6c1tLiVgwg6C2yo3bzfscvCD2L2y
sYlxH6n/Exz0f0wUjyYISYRolRB5TwBAgW5JQPMjcl/Tsd1TZaBbnw0yVfv5/iOaVHCpTvT+zlTh
Paunwk+liBtv0rzUN68vCRU1RMpdPZRt0BXDrdK3keJRrL8VJOT9vbSw47qoK8LHShMSlHmLWUyK
E/mty2ZvjYvJsI5opdCxduDkVd5wTDVOTJ1EW9NTb5WnAqKvBe086SySYJDDRbqGkyKSQWJhpvRF
pY9M547Ko9mFNNAyS1m36rPe6ZWXLjwHL5RLRW7eDdoCdtVYDtdtjDlXbsd0z8y6HghOqsnYkRBb
tJSveyYBg0X5VeOSGzNJhmh0usSKq9IYmZALU8lQ8Abxf9p3GkfWgJFNKTqzSns5Qy7A6ug4Jons
4ydMrYnKOcWBRaPbYoZyCdPGkfpAPAaJk4/Ka5SVqBPxzmdh8rcKVkj2OjFD0ssFVjVXGKu8egeO
A1I+t3NoSupOQznVK6NQrVVr5pkXN5hqkcjLaQ1tMIZN344UlsGWAtuFsV4olVFG55JImI2tbkb8
be0FXozv4W5BaBCDwr+jJJ8F7YG56JuzOi1cHpzfv7Nb6O+OGuAsoZWd7y05nC+rnO3VwsoC8uEA
AGYbIQfmdIeAeuDamZUiIhlxJ0/hP6LNJffvb8xOyql/67PaHwOHIorlK4PmnOQP8UVpmk2pkZr1
xPy3BdypNhU+h4gz6O2p4KmqMzxRKtc8lpLPGbwZluZSmeFJWN5VaWTmtEw7rixb2byDRHviUFQt
s92M8uU4l/D8yLPFhUk3dCHCBQh3C9VcgjIOEqqGcNL5ElsVfgYTX4RndvH/kMkqZSQtd1Cqk/fJ
Pw5N2rT0B5bE6+Y6EYSChmXPKsWrKSQo9uoBO4EFFvwqW+b+FYc1n4Fm3yLeClmECoC5wAXTY6Hv
CSEdR4ZT31tTjKoJX6aiHWFKYjOp8LD6Yfjne0XQLc3ksGWN1oaD0OkGi1nunQSbN5v/wgLhtQ1R
vmrmn1ypsZlPUcyliagYbJATbzxXBakT6Z+1G5NglxxM0QshXzf0x2PfN/i8rYGWdA5aKGhT3IZb
Lsz2Gm4gFTgD7asqlVT1b58uORjBq5psm8joMkJj7GvKekbEv8bSQdacAD9r/36MXbEDU4CmMGwM
4A3Do6BfP5lwuP2apRDNQ8pO2L7GB96lmZFoaqfIHLU+ChRuZO3Vo1N9VLFiciW/SNPExUqzZsnd
t2Mt3e+arccueLCDmkhc/NpTmniwKzt5f/9Oo/ORS0cdn6LgaFwanvC4waPAQLMrfSfzVdYhHiRz
fjRVpvQ3KqQ7L0MdD+80tenvBEg52g1tu9O1cM+blmE3ZhBq9xBpdCr44cwBlqD4nRaj1YtsMdkG
BQq0Ayyqk1JM1BRCFVYLuXM7WknH8NH6hJb938zxOrEnF6+d+UaPWTC8HLqjdz/z1o4Xl3TzIaZz
5mqAT0nMUKlBZ5n2a8vKEgiIJB0g5NnaLPba247uggXX9xIMCy18UKK6vlxEQQqK2x0e0NAm9G/b
wFgmUadA5UdOTZ8uUHtzzRqPdV83FlmPLbyAk39oikG/JeIiqX0qyV8TkBZ2jDIw0MHTriQ3/7bp
XmlTR9uDL2qvBuSFZ6ZgpgMUJJygWlRKGUNjfkxB43nHVOwxubVPyv1qEzUPdxJrDvTmXstDxzCU
WdqG0PDdZ4AbGdlSodWzuCQwV7nglhNa5GYRixEWqrOaFJ8lw7pc/oU5YCq+/m9awnN8UXcAlWPR
nXgkXRv6SxIodN7FaI98dFdvJVm5uvQVCRhHXg1FgUL88otTewUMZ822fcHGC2yG5lvn1C6j1n2S
bYmLfObrmdMWWXCzmWGmI7y6Ps4HT1A9CZIQl+5Ia9Gq8vvK7VGb6iUHG3T0s1t3I4lv5De7ypKd
d7bpvJBaENRTXu7NfKfRbRCIf3J4/FkUvKSV0WtuV8lNIbQ8tYentcXcePInTRUyU8//rH7UowtQ
EQPhHnsEYMLTjzxwgg/Usn3mLKM5EY1cXw8EEwvnVqA3mOU2uGt6npxiBkdHjQYH5vLXi7gt2nU3
8WXz5KBMKvC/tN/IbNRBQwwFGtY2hQL8Ek86KamV5SfYYpxJ/X5g2yth8DKMyAkBckLk2/S499ls
rja7N3LVQ9a9GIIWLdAIQH0QohN3/1okurFOVd7XhJb0fqiIgQTcvroGuwjXYoGHKaAewNKCA/sX
+WCuHrgAYeeHDJ0ZvcwLc9vrSoIXPfdShQkGEf6F9+FnyZtVkE3CMLxynujAzqKrqdQ4NNUxzu3b
HqnV1ePyxRomkcbYO8RjvNgVlPdgIvGRTLACAY1ZirAAoTvGjUY2o4yBh4nf/sR2nsEmPUQpcSIa
QIhhZeWeI1tvoaEZYpuw1yQi+s2zHXKP5t6aXGYtrG9qDQL959bpxeIphk82GW34UHCRrGd4olmg
FEp0HrwCpC9ZNvl+wgqatMWkwqme7npm7KHE1d3yoI4c3CM+ePmJOqmxfVfv52TgPOvXKoY2ScvF
tbNvfV0UNamaxwlDExioWQeaa+qA1tvtRT0MfQ3yUVWqLyQV7PiIgo3PfV3l3PSoXx+A8nWdr8jY
rNopzxyX4Sa52kCuvGiOkMov7sstWy9EVCXXxthgn/8+UzneSz/WQUohyrj8oea3Dsopg1nuwtjq
WmtVB3yeoQXuSQnXpH8lnWD+U8LJPUJWFAvRvw37lYrzWdYbU5sCrADGgTgFF3xyQhfMDnabok2s
6cOGVAt+vN7AwaVOCX9IC+WJ8zozyrbux+aCgbnAfqbeWlU5f5SjpsOndEd7QdebPdZpXii+0Y0T
HgsOX85KMhls3oo7/qctHXa24kcZhKuv5cyx6AUIO15XThmA+IeKVDgU96Re3MBAF0V0u3rt/qom
+OYgjs/EdNEvgvoIWOvT+K5ffbT+aM27Z99YYtaerw/IJtz3QLxZVu531bROOqTbTO7nUmkJRKyX
2FUwEBmCQYWM52jrAGYBPgtFqXUrOcid73mBJIQoYAy1nIczmESjV4POZ6QlkFq09GGeePBRB8mN
WQPQuX3In8apKPJKjNjM4tw2SFcX9I31a5c4P+68maZAK0Cn36+o3Q0Rs6cNudPq50J+9fMWrLuF
S6O6isDSM1QlVpqfrVwCKFpVqS93SK3a/A7UghwfMebJveTfPL3fOySjzPAiVXXfR1gK+fBhji6w
0IoyHuX8jcEK0UyASDY08aNXYDhctCMyDl1PzUZl9hn2szZe9kXrL7JuOTAZvdcMugtXuEMulLvh
dV9kl42FQ/YiXGUJyfccNspCRVC7UrabfpyZWzqbFWaCFIplxeRjuRILgMvBwBX2ouQrHlbtmaEF
4iWMTKg6KnrV1VufgdtzxRf/M0nwCR83ZHGT1l+MfPPQTkeBSNDgFeHf0VT+/9PiKfCLdtGKqr+X
4Chok31M/A/z+VH7/YfUbW8gLt3C8tq7NyzxNULXDB+GqpMrK54vrE3YS5CmzEBf4pBBpUuK+1Wy
Mk2eI05Xz31D1rfeNDrOXuDHu7JTGTZME2x2tlL5AxnLK/52bjdhupTTnVL8ZYXKNvXl2N1ApGem
QCWj3+gGYuImmlfq7VNNRxu08Azn9pzLoZ4hKDcbrsuqfrDQNKg6qhx9EKNgj4qKMVOF5opvp8nt
Qcd9IIvUXsNGcqnschRcEHkg6oUGc2KFu9U9PraIwz14XMXVHnGJ8bGLQqFFoA+8CKPwy3X9Vlx7
WMGnm6V1EMdpZyeXPAkNKx1suX+s6xNgY5hM1uRfnpkNChZZAX0HN9vkF3za23H5Em5nTANZqUHF
PXJRjeg40M7lSldIaDcR8aXjZmJ7Pg0uBeWs7WTBE3ulg+UjYyv18lzuFilVt0KAXXeLoHYaaYly
m9xUEBNL6i3sXKuXM9kbtKXY2lF1B3x2GxoXUExMDIZZdB0TgoT1idxL0sRkR6NxA4K4Rp6IG/IX
GSdvZi017X0NBMBryJny5vjAHjSEugQM2eNPGqu1rkOpaOpD15syUTQ6WgPBPBc5i69RN55qhrEr
ydT64/L1eBPYN2yY06Agtn2aFGfoneiL6QFoKFnloKPNG27DY+zr8ymj0Sn1RokJMGmU66T9hn7n
2uGSRUBeJpYTwWhF+Q8/SPNHIg2eC2+8btxfKsiCrpZ0XOrRzV6fG1W/C90U3dGGpuw3TEHMBQvZ
tLd+PXB5dYlTkRyRDZzWswPG5rOoxZ8Wk1MEYfVnoSMCgwR+4JZ37dJr5EPU67YF9a/1Ce2P6VLg
kB4ym04qZp5rrCb8O3Q8Z3pDCqufprShh07huof+JE/3DNyg4zIj9m4ZZWXvd2u4n8zrQ1k1NZ0N
3X8KB2ZId1XvMDxh8HNpYGKPbhWMT2oRkknafjEd7AygG1l5HXvKsfkLsY/vCX3LROIiz/LFe+Dr
c1gj6bpSyYlhOQBjZoEI4s3u/0bylZ3sjqAFWiaD1wKSZzv5XyAY7UdvtPbtWlXz3jT8AXjRU6+i
KV5xaz3NVWkFcfq1XxBUEyZggGiKcaWsYlskmKX6K1dC3jce4tla+WopdAOPfhDIxc7cuWDRO3xJ
nQJ4Ruom4T2Ru2Dd+WP41hKN8LaHJ0OhAJpnokFLAx5kLk29RiWqGRCqUGNErWpvshsqAi4bfbEh
ZDZMALo7GqezxFyOgfgCOEj6dAF9gyDob7VxSUvL2Tw+a1nRvh+vjqN8udNyvcAUDWYiwhXQJrSi
IqhYhqhZrYEqcCq1GBJSaBe0X7AunxybPZX3raYyT+q+1dn+sf/peo3NWF1vXbKLCSOIVF9Tlu90
GRL5Q7zxsxu62BMfE5c7L0/lTLjkAEXS9+akzZzdPh3c9LIB9nwDboLF5b7nHGnxGen78fi8ldzY
2lNwH5QnsMWBpZOPSLCVK4YNpol6C+//EZPIigOnuzXA1wLAS5oDGsEY9BivRm7y3JHoYuCpb+vn
YrLtPX0BKJU6PvHTc16F9TnwQ7SP2dEXQ1SO9hu3V/lyqEvcWgJEBdqgPzOnItCofE6wT0qiNPHD
eKQwGiwzZc/JIKhQ9kQIuKsJmRdpEqlLQ9mPnyOUS0gsFMxoeoNhaARrZjTrXVlds69XCMZ1wibm
V0LSdX9l8iKMJVW7WAFtF0+WQFgQAFv+a1cvu62jT9cUpGH6xpzuXoa7qCIUiYPX+PSwi01YgEn8
ve5UmiZsybYbf4CKzRQvqxVTElMxnjUuz7/yymGO9UwwN5mFc53+5qWkokJIaQ6xwqlxMXrwkR9I
GYUcG3ynnwi5u3Lr9E+iyHzrEabtqHwxUm+o8ctPrf1xVQrb50TiTSWZFqp2RhXPHNX2HC8m3P/e
poQnOgrmCaz7O1xwt9dOD2xxiWV+ijeFE/jctKdEUczW+VonndICqNUq2NSwUqZQ6RbsB1OEdnZ9
7l91JGJpT/IYrjzeON6ulIfwyHa0cKYLc5vxmBj/BXDNZBxo3uleMSUJ0dAe1+wddE05jPYRDkUh
d7OMq33ajkhn19wPZ+C4QfPGVpsr9FMsIWyyw7PznG/g57HoEhTzz2BvCmikKmJYBIDxwO229ogN
Xr+LEezq8VxiSqk8XNJo98et+Ua42TUaFPWOPMOoPyLgM0izJbZDP400ZBzy53a+Jtj4GM3jDwti
Qc6RenI92pRak5x9f93xRFSM++YhKSJ//7qq924IJGvaCoRXvoypU1kchNZAuQ3s2A7bnBnnxX78
T0h7QrankPyyfxCP/kr7oQZxTtiI2k7U7aNZqhI0apRSf9Dnr3te2buoV6ewB8QnOO94Gsky1hFY
5yGcgn4xpCmJ6Y51Heowj45UfnelfeQVN344oruf39f2SbLHlNJh5wN7b8UrQfRyjc5y04FPF4MJ
6OGQygvOFX969CG3MYdO08iLjkZp8eagDNCtGcfYS62wKMUForvqjo0MFmgNpc/gzUAIYw7eodQN
sG05dLi5ZzCpuvnvrm5V6uKwLSrshjESpUjC2ehIKh5u2gNE5SqlXf0Vi7se7UPxoUzopXfBXRO4
209BzsuQZVRMpJ1LXBLTqk+cigixZ2Mn8WdQOKiO3M62HcZQ0Y4gKhqZbd62JsP7X/vpRco+GDBD
r7Vu5bbOVbQ2zTqvw13gcC1brk3B75gvpVLu7LG/FrDOL8Oc42H/zRqFMqYgAMluXC5DZnTEojAQ
ypAAGqn0LQ6DU5IA4P6rWiBLR4uoTs5jcM1KCnrr7dHpW5yVM9g2TaT22AzVLWEyN/1+AM/sO+95
qhOuKY5lwwVefhwk23sbiO3EDt8GghZDjHEfCtSYapiTM6+v6eTijgO9Y1mhEznWsnGjSZOIL0Ig
GpIasILA9Yo5WWDpzrb9YnD208KPkCdb1Z3BXYt5iBNRdWNgZiT0BE3+4W8PxMOZIqvJEAJ8A2y4
TosXvaRhI6264RG5jp9lG7BU8Pz3JNMJngF0UkGRgpVA5nAW4TCm4Y6Q1+Up93OONlk97T11g+Kw
IFMK+xIF+T0v1d4RsWTYIbZo/p3Fbq1JXzdAb0RgFXTY79jC/SdtOSBDJI4GpOMDY/yBEZBGs5Wr
UpytUS3n+ZwNSKaVHKlM3O7VZMC9ym5zkqnXTIPHKVDzMfUFcUsaMlvK9R1MsBx1Ez50bVEbbwm1
i1efHASt6OjCL+qJg/dirXZJtgXPhNByWkUuFmWeaXsafd1cimdoZ+XhN6qkHqUy+J+EZRdeGjfR
T5j9OTC3AFUx4sEPcl8MYDctqGVfnP/Wb+tPv1Jgj9lVvt8aIclSCesYe+C0EJQyzF/nx425oRH8
bDoCD8szI5p8JFaG+ckGSXC1XI//+LP8JJ2jXKBsy/Rw2YrzY/ngQzCRb4SFdsepTN7yAZdh7+az
/go57s9jx1wNW2aT/boHTke6qHu/Bb0Itzd/aIYznM+9eOco9KMfY/6BuhBUDa7xby3B6E8jLytR
xGHrSkExgCk+dLgQq7tl8uoI6/fMpavpjtV9wMs9Oo0KQ3dLSfd5+Ssa45t6Q8QjGo+qVlV8WRjz
bB5ZmwECEyHilJ54Br787+G2KWM108czOsrszViOyt1ro2y3nxmpRqPLoAqVhSxwMD0bGK51Og+X
4RadmFosWvpizeGpy/kr2s5NhAN4jRU8XLNtw/pORzGJG3eluKtqvpfQxhJlPK2Tavs8jT+q3yts
HGTND1VSw2IX2O8PNJcrW1L3YgYtq0CXvllH83uq4UZAvOKEXU/PMsnuHH5cIHDj5TI47k9PWahi
WuMF15CmQ5kXIgwdbzPUcKYtoOZ1mw/TOKC2jsFNWWjM+BkpCYtsD3zQlXMfPho0K7Mtsqe+vRyx
+l3LQHdIFo8tMMFJo5Q/4gJyWyRxaWdpP+q+VpzSYT6lEumQTikJCdGFjx/HWa65bWKuhyjReJMX
G/3+jfjivxN+J/GDogLGrZlcf3XdYrokzFLWSkDRxP9z6KgC6xwAukVS8is7XITjUs3s6dLS56Tg
LbiT9qL8/XCMohHbzQfxT7fe3xdboPctj7ewI1du/Z/5cAmQeBz0m6pZRX8i5QVpibnJ1isEhCOe
LpyAcgbvaKIzOLGxWzBIHlftSenQO2+Rh9lWiknEgPZw4W8hBWGyscY7nAbnaLqHQALXgDImn5EI
i+jE0EUk5DN/iVlKXp3uSRNORreObZzgEfCsIIboPdO+QrZ2Rxe0S/sV72NQjZBTpNRZq1wljh9W
eik0gIrQBNDyN+ajX7p2abZyM2OEFlamYxSwPnZ++9TmD1lk0hRXJH/ZO43whnzLrye3oRRfORHb
z7HlUHJB+cT3rDOSBrrE7nD9Vo3kBJlbZ8dLMwz89Ko26KjIjP0EyS0/zpBInJAuod+hxXXDas36
nzLOg6tGMSCPoL9dz/F4cfkuF86OFNkdCOoKAKNBYBpOSED/56M4b5P3OwoQraI+MkMT+QgKvleE
GFt1VuGpWh04nzMAs5B/+o8sMdwyvHs51L4oF5GVdIrjL/1u3vu+41rPU1ndVEDFWeSJkdyV5T4D
kXuqItixUyVlDT7OGgUAOExFFcufcaXMYyPx67b2LlnHhn6CbpVNZKkwEAhK55tSP02MIg0OlyYe
TjpQ4IYeArjMNwXzoLiZD6jjso2nr9StH9Ul7d3qkAQiUrgDg2ky0yNpfgeGnfXjmfhn3D+6J9g8
kMRc7AzuQUmnuxCSh5e1TboGt0ytEV3+2wi7gCvW3f/CtMElxNk2GZEhZDM6MNeMgHb/GuZhqJTN
9jf0Bc92WBM17eRTZpRGncusiLjaiYZmPJQfaiNo13zGesfCqXTU7Mgs5Jlz8iedpQIflc+hJn3S
Ir8osGLCCPqTfyuLGXPrRKLEkCRzUwNHpLcuRuWtiyiiqKG6Ox3Wphp+QRybxy/srHFs3EF7PoHE
3Srqvn80i99MOLVE7G+Z1zqDHOljcd25W4A6z90pShjF5sHGh6nmF7IwvFp9pMU1XtlFf4/YlSs5
FTxRnGgPf4JwtD6YqT3Z3zC3p3vcRNIQ4CfF8+1VbZmTBHv2aVO/GLRcM6kkpdrrDI/uqQSjZc0M
SyI5UxqQJdsj4VfT3d4T786PXx6kxbK2STmW52bH84B/VIo8Ef9jUu3PptyWnV17HCuON8OLwv9i
kfhTFpmb8qNB6aXQNPOgDMSoaCGvr49rtIYYBfltk0HneQSNPqgrPpgoKhJoWS8fqw2M/fBCVkZU
8/HLJgJrO2KJc8SwM44B9w/cEsyBADA4wAcZiyp7GZvEm8fgr1pvC/ysZElxbXpz9abqWWRe/fA3
FuSXW0Zz2cjc7jEIJwTFIMlyaqdmF0ZWV1mBUtrQJbfOv4LDViUPN+8nWyJrYi0pHc21X1vJD+6w
HdjqtiWxUte7RthnGRqron2cBnAMJ2XeoGJQ8mJJvyFkX/Er8niB/La5zuZW+1wGWw9L0fKFQcVY
ZbGAvzzg7xmxKUqBNNoaxrx/cVMA9y+IvlZcXjxeMAzBu1qzcDnm0o4pw2UIDuIGadJRQDVTdetP
O9LoKXs0J7xIEs/emSqBgziMtpI1zAObrj0GXLAGxSMZgpUbzOyjL7MBVmLtES2kGhIlDBX0NLYG
6VSVZScI+/yVB8h5GHshsLzqs7Hdgveq1SR16tFqzJC9fGaCgv0Xk9WOd7tQdbRvONzTJ9R0uAaX
zjosghwfev3QZRwEiJ169b8Aq3V2hs9wp3Dn9gVie/LZ3NuLk3W9c1957Qi/If4vpwiHOC6fpDQV
pHGNw8X0ZqVLI8/Q2eN9BDA1pHoQbFQV6cvL6/2xzQjnGa9DVDfCwnLDUI2XkDvq2G0sm6eq0f1p
CuXek4wpgGi2xzb4FvHdAIlD/dp04KMeBIqJ3zVl9k1zTsgr0PTMSANirg8BQu8dpljHSC56mL2p
CjzI9QkhZ+FJvUYSChVoml2BiPsWyPEtA9f9LDJrqzhPPLLKKMRX88avp0Ks0zpSavubPo21YO5Z
pNRLQaG3JSopz3yt0750RC3GrtecM9ASG//LxAHzYgi6X10Q9yWaT7Z0khvrQZdXzac/Yes3bIG6
vgdDn9xEw3HhW4T11SpbB93Ih3kpvT725QbrgpdH7lVqPlpYxVTX3+epg9w9Yzz+PFcdQT0hO8Bp
FEowss/2EOJybao0P5/MBgTmUhGtoB9OI49e2h/iZe6nv/scyEQpLhmkbzjrdqJRRO+40k3vUgL8
UMaAeEATD4If3Fu17OQwUZt11aEUM95B9muoGJ0vrjrVdWE8qB/r+NNpakmVVWofVaAx0lR6wG+K
iz/EexU9YRfVYh2ypOG8U0zHH6Oq4DImCGEZZyrfwnGSuQEVQr5B6+5KobJFff05r8A/P41L+edG
daZPYdQ0tU3UUc1i2jYv7uoPANeOn5/JrXUPiOkT5hFJdFTB0R+Jxq4/xh1TTGiCYka6UDccvkG8
WZzKpRocM6zpSvP+praCma1oIjY9NeL3WfReG/Z5N4FdzGxq4MqYdW5CTaNEVt7TG4ek0K3vDtE8
aRBuQSTRoUsbucAM1O4WhxMHuJfBUK1eEHhPRsGzrmvFbvU9Blsmv8on+fyWiIkgNmKozv7F+EEy
aIxI2HWjkBWYDZzHUKwgrN7bx4fZc274MrdvVpPVPSxOdYItNch/G8xCwS+K6G7JzTZf9fqCymiN
O5tb9ziPka3QfyyC0I6vxZBCS0vAYeUqm09t3P+2JI6KEDcyzeWcjDmuC73umH+YQHCHozPyIUOo
LIQg//4j7/qJMLbTsughPEokaSLaqFQOz2VQFtdwaYr1znOKB1CYWW9UNYjQYK4Tgwhdau4NAT1z
qn/uXQhfVOUkM+PfvtF0oW0q+16rkwIZnIAurg+tiPrEDZyGlZBk7BSa9/PATeY9VlOs1QE0aSqv
jZyOC4RMzrI9lo1J30t8P4aXXu/Aauq+usWZ3fvHzVjXMSHnQD0QvPGeCYzJyozQoI2nmoPUOFOz
1zb372adHJi3Cn24KryjRBxsdCpVMyUXBqn3nIdLTTz7XP1wr7BeVpmZbXAenrx/O3xEhiNDgE2s
YEuBcM3AsTTds33LEYEJoxjYRmW6xUhnNgUP3Z9v/RnSGefiHQfRfy1zKv6KO/we1pDw/m0HSja5
km9A8eV6oyguq5JFdBnnpVzmTx1qW8TqV0MNvxxoeZDtuwCY4BxRqQn8cczsVQ51gcujJsrjaVAz
NL/Z/8dZHJXU+gZKTAbFqpODhb4kURwDng0dsN+/hnkWdr3KCH20tdUyvi15Sr2xQlXE0JSq5DO7
aE5jgtPbvhH+NeQjzrSXVlopcqQzLWSf4ctD7bbCKqSTHkJBSv6fzU79APRs1AJ8E3K61QDSL9Yz
LslWh6plzzz2D6y7lxjxqBAnuj0yxbX0rr8H+ebYnIwTce4hkMqr8T2FZa/7z2XqFPz82tvTnCOl
4KcH/6xfsp0aUMH/KGTUXYwnIpkOJ7FMYtntByToo+NDF1cAdIgvvU69ko3LiHM2zb8eo+2Dsc/s
yN4+U5fYIiYy+VsmoMNhKri9B2YL+CxSuh5oOWvUNuhcGcsPskO2h2eeSaaGaZ+AC4DyaBnthcMv
aZUKFaLydj+vrUb0CULBpTEHYwn6kmqu+uSIu6p2k9Uky0mtxFWEksGHmtLvTgk/EfSKHPUW6VqU
dLOWp39lLt+egzwS7jQ1P0L/PA24O2vW5Pr8yP3ULG+EQiPtpbHZRSNIOwn1XS8mx11SCTumS+PT
sIbrGV+thK4FDnnNQi+2HFGPGXXLbDt763gSjTDhzsjSAZbT+8QWt0A97JIL33oksWsAZIpWYvZ4
M2QcogHkIJl4A0O9KEzgdJyyTFEhu2Up23Ir7U9GSbazafYDEE5SzoQs7CgnW3sjD/cdHvz49VB5
b5VR50NZS7xYORCK2j97dCwo5HtUrNV/uEBU3XzB0Rr3/0wXOzGzHejWjck7yjvfgbz/Wa98kBSt
6f7tLEl4EltVcrPvaqK6p+WmpYvfb+EhT8nC7rpnY5hTVu/bE/l3ZpxkPLoYxuPARtKQ+/iTnhL+
eP0+mJgZl5RJUMUNcqe7V0kloQKKJEvPvPsuRcw6wuHnf/q8bkN7Ta+QzvMc0aY6fBzKblVX6lvq
QdRp7/e7wHADE3CttnjMcM0PVZLhO6l0m4/KJ6dpuZVQKWQAJVSuqVSZhYO0blHp4gdUZ1c/NwAj
1oqGhEoOGwmZVlpctUVphwH7uzszclj5xQOEiuTXdsbrMjXEyYXw/X3E9YNLP6nTdqa4z2fenyXe
szdhvd6XhcN734anl/eXNrbT9IWp6ExP7ylBB7JmGESmRPeD06VcxalpsptcgoZoqXfCHeHQnpFh
UOL8ddzFgyDEt64igXr3DB6t8KgimgS/jOW1Nsxdm1Fcj9SqhbLX5Qap/WED+T0rKoRHuD+pt187
6Qal1qNK04S4qSSQisg4/NJBkYMRpD0w3fa12ZeqPC3snXRBHwLFOPBATz/2g996n5keqaXHUxyV
6IptjtnXrrIcP54UYyjm5blqeKSEB3TyUwgefAvPEb0rZdnW1nxJK+mwixOYhaK9mKLIzspSDdtb
wLYGaLpAXtQTPyVhdmb4DD02Oz+MvF6id3VZ38cG2QR0PU/WREEHM2+1AiuSmuD9bf7OPAoDf0/R
cfmAkdyMfwD3LpeR+1JgHhvBxXAdIcPAb0xP5pZuajYR/TXUE1FRmlSVd4kFJpMYkL41mkoBjIbY
BypnCA0mVwCBn+TqCmuDMeeKICrte+ROnQuZkVKYN9nOoQlfwuGy+E8NHUph3mfd2hDl6Iobuxn3
R6O/zc5XD5SCtk13O87n3Le7sjVyvXsUWXMadhbF6tm/K1WMQJ5b8E8ITkpwy+2qZJzFu5+1FMjR
pd+WdcRTu0pfr4zi/SeEkNYOFVswt07RYB9Qtx5MkGgw/6uzvkw9OvaX5qYwDNH26lMo9a0HYBDR
WOcFq3BR3pkaLShnUAoVadH7ObXdhrBmvGfynOP/0gJRjIUVpMUYrZyOLDzKrrju63ihomwqXjgn
6UQOXE8plVBJwGS8Yv9O4nslZFH4bf2QYjuCTKrqWvBf/6Y6yfuOkluwp9jcCvlm8pZPNUIxl8zC
0U8KwDcH8atgzfqES6zAoQvB9CWqjDt7XX/hvH3G7KoI3RTYA6fMvxKwh6yN/qPaFENnYqUorH0f
F1zPXbqTc5fz/FuwU++VN5IbcgQYNmmjVKaaIUqke/m6gXINKVTnmSIyvztOSjkaRuW0OsaSJOdZ
kmj+YSwV6AcHM6QDYYT1+KXWtlmlQa51amuLS5PxXBcOUtnKZOvLodBd8bfUT2cU3JrDEOfudd3c
ub8hCZy2CBaeOBx4r0CTk1g1favIfEbxPk9Q3cg0pe4LPc6EsoIeyvo/YxNvjRYgGwUA7YCCHTxz
jK9vR7Uv6EacVqLaTrxmYHHd9Ox6/bF59b2l0k2qY9v08ESd8oMzS3BTR0GlL2cx9mCD2x7EHHTx
95C1n7KEcDHfeHpf2v2OmUW9blJ0u97tMyiQX1dqtu3Fh6j0w1+lxZ8Wi9zVJ3ATGI+Ik5IZrHgo
nDi89mZjB/kA3b0iuW8JU9IoH/sq2W6AqLWMRO47YcXP+MBiW+0/tKQx64qxWEq+7hnISVRFsw3o
hSFpXTUsAhPvMxwsCeudOhzsn7p+ixnQmbSCMVpom8B3O931pkvEGRBuHK3DUfheE5eIuGzPszGq
gtI1GEUQKt44WmtFXSVvcjzft3BcYVFHF6yIsSQfFg3VevADUOjVdkF39mAApwO9wnAroV1oiF59
dekGODfweJhJ6DsmVmrtP37tjkalj4DBRi+Pt7p+NtXi9ijG/uz1WxhPDI19tbDND4vGeMoWxqBu
ggEjnfXwJHCYJgxBQWRQGboBxnap230KunAZnzAsMD6aeCbpIAp1NnNVEaymMvoWGIRbQXQnUL2y
ql2eDEUEelr/mF46qehhyivD9uDVLDkjzzcSEaUeugbPwa5k2yWCaV8ODcG+RDFNfKq8Ii1G1hGl
IT/90qVXxXu5ihjJG2zPWr4MiE0VhsDeVRs5rkPehTEd4faoXDKP7V3kadd0UXlwBQ2bR7uEqefY
kSAzXLKUTIfDt2I1olFYpF0z+tv+8wsu0c6QvsFl53SfNXg7mhzBBYB879Bb+uvIIG8xQ2YypYsu
7P6Kc8xxR2WXkrtUy/gwWc96LR01bVSO2yEgUx2DpLyDKqmvKJpzgWXkR2+OCjYVqFf3EX1Vi1a/
zzPu43Oht+ekHTa5nuHN9bq8vAWvDSBgasUqw9R/sA4Kk0a/p4lhJqdOxgDDJLuY6cryuhGB+1WI
dYaHYv8YT+3LSDW7+jx+5h8GJle9btTdnNTKZKvdtE+tezGAVo7isE+Xw0kXTgoATLRxzdeipQuT
WJglFVYasvrURzHoKYDxiXAyP7HnC9BSd4fCStYO5ZEUNz903b9Zz2RLYrUM/7VgV2MFk5xAixbs
UMzHDzOfgW28yPdSbvfBG+4G6OKbbDEarTZVgFsVLrhoyEg60mW6o/1cD9q+crTzmVLmcL2VUYeD
3RN8GAjLxAhbiPaB42Qha/8E/V6ch94juwMRfu3p71drxwaPE3nPh651DNLyG61Gsd85gaPsVM/o
M566mYIz1H76w4d7p/DZk4tEljM5L9gzww/Qu5ZqwlIp3r7fvXx0qJui4eVhq6me3lxH46knEkuM
q5tTeqZOuKSei9tQvlmlrZQkEywzEx7fRF0sVD7XcYZENQbJkOUex1viLN8cr9mECN7LsSjVpeQx
29teVqCSsytQGJli/rVn4vWq7XDWue/V0WxOIsECTU6zrefijEiYCwP+dEZcUxv02lwOGkO36s49
EYoATVg9B4munvl/nJkkBLFQtDns/MLlSexd3txzchJQLOxNFUcnKxcywaPJVPJPyQRjM+Wml3Qi
3IZEzUQLhdpC8CuV/IVNvg6Chs7ui2fja/isICJxVEsGo7JLajFXn6ZZVBDCPMGjeio2UipGKsuV
wphHY11fSy8EtqRJNWnbXDnGtvT11G1ZE7utdRO07L5/Jx6yPZZ9RdP/RwsLnfb+GYT7aV6EHO0l
IWwhTdCtOnVXrvSWox+F7cO2BQe7F9USsDQGMuB4r0yWEM9nGH8ptB5nZOnMBuOhpspTCECtZZQG
DG2+J7PuTh8SfhHPC4FfDx6bpXyji2g6bD7qh523tmCjIVk8tUzg6PiIMfWxHKex9t5SRCtbskSe
4DhOCRDrahNEEYPRTEbkgmvghZdy6ox6PtvOAgdt9oMhHosQzHx3bGgOOqZI+Ea+qmjb0zvoNdoW
ngATQNTA/ReBVGWrxUemP6wC1RSKc+SUXlpdokwX17MlrJMpvMNaAaVqVH2nNPFn1gBRZjcXDqJ9
0qTvvlM9jOSWWWnhXPjFW1+XmbRgLrXKAXt7ht1I48f+y1jnTYlkFovA4biCYatG6IbBEcOqU/gd
5D4dnu6c3PtWgm/Thzwv1rHdsn5OCCgpTF+PN1qANs4TH2szTnuOPrtjP8rKQfbitQgd0xkrZbSY
5bDsHvCMayTjuiyg1oYaqZEtR+RBJQtixBNV4GG5uvqv0Bw/UJHbD/pyQJbUKsVzBTgQVvcZA3tC
58mYFwU1soR8J8+Jkbw4Dxl4qKlHZyhdkc1WijN62XKrDjT3g9OIiHl6VAGn4t54JS69LTAa/1Tq
KGu3sKoN7+TstHrauYl3ZjK+xOR4XE8Ez2TQet2PizUjCO+kIhay5h1cAiujeiZbpA6M6FtqQ4gj
VgwxjCwAZ9cFqAHofusG1vsAUenuHxZz55zPSCrhdgHozddvAE4C6mwDQsI15nMt6ExBo09sjk76
q08mc+zGdjPVFhm+fCT807f3BA4Ht8DePmABhcx9lr+h07xAXg8M4VPivLPKAtHMGqKePiT29Ihj
VsUaZ0KmzvLfZkINXC9PXDIB2c+OZ4Q6s+x/872Psqg0MXmbpxvLtPS1P5qMwfBd0oTW73v4Icu0
aZAZ71OHppxjt6Rh56jxSOfkoEpRRyWvljQ+vt+k2TP+E/3SK5LPC1RS7hqbrAl1lzmE7PA2axdz
QHbWAzVeqmxox38ICoc4wMv6K+FTz4o7R5p0n0JAbbIEb/oUWoU4W1i8Dct/ZTdI/nteEdkSCbzF
DR5e+JL8DWBPJLSEEgrMhZsU/CU3c5MrHoOAFgFjOAdf/bDKL3GyDhConEVP7WjxkRuHrAzsngPu
uLLhtwZXDYBKFc51mzp7lXhRDeKSVxtmG8293ELOJaWZQglcKcaEhqeZAQ4PM8av/5Vh66gOywL9
cmPF+yt38EL3Aq29dzAHgJbB7gqCJVZYJnJgKE3czZYrDt1VSVPMXZM1bNEZPRfTrYmPOEFyWG9i
fJHhcVZOsa7NTj2ljMPFbJEY6Q7vM09aEHtL72VLjmHe44JmEVtFXkEMCxTq1fGQIQjRGr7idlJX
ZQj5rFZQ4s35Q5vToL70ZkLl10yiGS09uoKAPUouzMherIDEqNmy5T4SIMxEhe04zWGG3HkaIYak
1f/Qlc1Z8/VuAMqAIt0gM0c+a3bjhV04zYvjiycWQW6LvLvt8GSzAVUELd8+17RBubkKnj+kU/hK
hyVO7Fh9+cSQnsiaed0n50TQ0xFYhZhUnPY5U9GnNWjEPpYf7G2q+F8CZ6kQHZVVVfmkvCahAHQy
LTslC3fBjFPGzje8IU31Mkrty9IoqUPHrfKvsXqBhJqHkZBU5he5MrvPtSaXBZpX4dnF5mRIKBJd
9HLFe+tIg85D5uC6U05kCJmKJmRaIyDYD3UNXvaF/7X25215b1FbhrIWYBPi7loAZtnxsgxx/pl3
F6KvA1F0lYHLPw/B2zYtk5zNgg4y2XlroHYZ8gMj4+jIXI82Uh0rdTxf/8YoJcsBqrHOwpysNJLK
3OOYmnYCHgAg1PQ5mZapyKia1iCz8iG15GLABITKZ7tSFP4bDqR57/ADH/fjmWKgd88JlTnU3AAL
3jzsa65qolQlPV93VNKbpNedmpiacb7q6kkd1geS/4db6tZijPLce99cArg8dDfgNnq4R4hg6lnz
sBEEdjJ81Sijfk0NyU1eTGI3LwF9IlyNorYDLXMZva2qfWttxOgRXpvCpN8STIyyMcx15kpPH8cD
lz12F4wJOgNZz4o63Vg7HqZSezzt18JUweG4Tk8869UYYflGHZI24WJSS6a0II6hnA1+iuqq5BGP
QtvdKq+vbbUkAamYYKJddH5PtpkspwkbD3Nx0nF61k1Oo7wy1cCikiKhPbxa6SftRbFuw2jMOkiy
LzTD8J9dSUdbWidQ9cDwRpSKA12dCrVXiIUldQme/E9kRpwtevDfsADzS7wBFgUby5cRfKzJ1gQh
dR0hfpMix/ipC/ZIRTXvBgfYbAhKywUtXme/li5xwnpgcOkewRmBrDd9SEuYfTgYFYh15c897zVf
NqCLtw4615hOIQWfHk6N4hMel9QvXqfIiIjH4tTPXwf79Jk3qL+pYGIttgNIp1RA1qpf6flLW2pu
wBu+59LCVcVJ5aqLT4PVzte9DQqVfgJudf27+GP+tIzg2fNFVlpCpMEwLMAMz4pwNwTSiX69opFf
u8+ZbXL2rpxfkgR3OyiFQUBF72tJh39znV4y9NR6glCnKefTPKqPNiJQT6TflLBzYzh/tLbZ7zYv
c8UMYXFMWHr9P4UzDkyZ0GiGsaIrf+Twdqw5CE9lR9SYAe+6mG2ZCg3nqSzfq8J0+11nAFCpU+yS
WL5mTXb/N/rwTjnsc90h1sAKvWNjBRIRbU3pVsTJBXbraWZaItYqKi4h24bFoBrPrfdG920nGWPp
anuSUGSAsCklLPNxU9c2OlBkvUs4/uDf1uLRbxu9XytlUKOcMO/o6c+GsAXnThLoH2QZEwggifZM
CPPKEqaTt/HJvaO3b+nB6lDjf/ErjtwITXA5LScIOfMBHfHxGQ4WipDsGtQlulkIuiDZO3B4Wv+y
5O8liLxEPI57D7nN2FEsVKW7+fL51gxcX12kH9rkY7Lx/BUyugS+Xc4pZ0Gcs0hoPw27ONVo2WkP
2hIiJRPu0cEKjUwHUEBJ6SggRNNeH/IQzHtyetDcGToxn3hCuhRnvVx9tGqVpCE0UMICCABOCVLg
3C+0A9+REAS8kstBbB5kQ26Q+6IjBd7IHwyHJNTi0OWiYrE1OiGEXe8JvJwuBlVajy2EhBZCs5au
qE5ynha38PbgL3A3jCU/8wlNMvV/Uoe+RY6x1gEn6n0/j2Wjsb6fytxrx+qZkWcJpicm/ZazFrsw
kbCwrYp0B3WhhmRli/PRf257u9A53AHpnve0Lac9Ik23mTetin7TO8X/1bf+yJwUlskV7cfVAJqa
RAZ5xk9MIsBUOx8QYQ5ncbQkF2K3/ZjVJHkSu1YwEgOfO7cu/X7LlrlQY22sum76ZFjC/WUp7nl4
eysR2VE03F6RqZWkODgxCCMqTZqwdyD17XDZUPuIKLU19pMTKFy2tOZZ/gi3aTRT/kglcs4n/ktY
XwIK593G5G4cRAVFV7Ofv+QnRG2LIOeV2XL5nqxh2n2fQI53lyKhqlvHUziPj2DG8XfuFbcTlWPY
S+vxhL/yUeZ9t3hgKlf9C+P+OzAwYoFvvwGN6mrGnTt1kzJGRjbKK9cEALeWAUrOImecFgJ0hAsx
oAp5dCtqCMACQj+1Y9nFftO4VyLr4Xe3JYk0ABP/hkcnZ9aaOiXAJq2XUFgaCdWdVygcozo7LUHT
49+Lb1B7tkDzCofshbAHqFWj1sbhTKuoR3J2R4fhTJt+pSTHJQydcMk6TzkR9wktobosT5OZV9Ub
cxRwigliPMo3aFeH+cv03w/53jHy0mF/shYGaFkRiW3deakCNg4PcbygTjoBPkWvmlr/Y4sHWGbt
tJkC6Cfs1mMNjn0R5geW8aXdxk9IVJFwjcE+RC0H0L0Yo8GHva1l91Wm1fP8vDzIVe+tlNuomaB6
Vwr85PA2UCtf9Sc5aL30b7phGecY98DHwKQSPho1qUfWqgcEJtMM7yynA0z17Sa95UKq63+Mw9W4
oeV/Q/of87SweEMpdNlLL+vZKQe5sAPpMa/D5i5/g7gL5y3jZJnzvFmFZ30hThJTu4UjMzZNxb8h
y4yl77e8ChrDuEpUxYllAovdXVQ/VLx4adbX6zQlsKx1L8itCfpzvKH1Wj1oFFPeczMhCIjy7E7h
V0NzzUKl76+M6Ws6Uo0Q0vhz0hKq5LzAzZaMSyb7VlgBkmHNURwHkaZfXC7wYf5y9rd5fdEG7MOe
eWAHKZHJme7D65uKdoBIog8JvoRW2bpn7hn4/O4LdNkBjMlPTeOrBYgg6aZqcHYvdOBSCWPW4Bd/
Yu/zY+TzAHHskNTpq/JFfakcWTFOYXzZJw5ELp1mz3qdfpdBIBpKHBxB+NdWtyf719IKBiszShGU
aqjqYz1gkEqRGBB/vwAd6dyLGo19xU8dFEg8prHgVhSNoEO3O9R/qS3ldyulUBcRVfSdE2SkysSp
5OsOhK8Rj40msxm98PoA4jmMiOVU5DpUS2KclrOclxhunaKbmC/F5e68dpZzfj+Wk9k9wf3DGwq9
LANXO5bAR3OkxI8aFXpHQJYAMIsyTRpiljcpxEV4dVs3sPuKyx8y+sq+VHZ94rIVInU7/oRn6cNJ
itrp6ItvrgYKO6VjLQMmAg6ff1u5GzXtjvBfOOOVnulbBFpsbBuTaH4USWkIO6Enm6nmNiyJFqm8
eglmhgXegsP4o+bhbvp442rbRmsRkaLBg56qobFZW8+zUtgJasX+khBcLvRfXMVtHpmMOuxUB59T
5+RBtUIzYdZVWx/ZK6fTlluZU+JzZvCVg0kXO/UA//CJ3m7hqQ8/7BMBfXmLgPfKDB0shWF4NA5l
PXtBOuDK6zjewt4QJIX5fdejlFSvhJ4XBv3M38XQtu9Zvk0yiCO0dBtCiIr2mNWc2DVelP91ALtF
vzvDW3Eb4HlTXXtwf95yZvf5ROME+nEYs5ku8ddFAOF2BRUModK3Vs7rLFeQc2eZwiXpwUH7DokS
OGQzBRr9KgS345p0f41+ikgGKd1P0ER1mFTgdJJlOps8ca9gYug7tRFO3uolX5vT68oB7ukf06Cl
1cSCdvpaeQDNwxlwpoHG0RgVTa247de8rhvKGwony5ptUB7cOXSym0JtQaEyXeVCu2a+9H4vcNyw
kyR86bnSCalfnN3x69/Wqe4Zr4MDfBnP3E0ZbSGqlmNFVAH6xtztcVucJGENw/0k5UIt0eZZNqa2
StRXpNORQnrvmxmvAUHwnsIxArRG9YBsLpkFwjmh+V7VOpC9IB7KRzll+oyN/ZCouP5naOotUGwK
lDlsIwJ8bhJe0nIfGnXKz2g1Ua0cDN4w3KOhCZD1Ao0076w7qom78WSLgQyBp+zG45+0oCs+S7qV
8My+ElsmsSbKAmVAG6IxlD7DuedxJlx3tG6rZWHcSaCHlYgfxaclnPeMNEcmj979GRnqrq0mypxD
fxJ795/C1nqTGLEK29931nuUAreXOS7P8wj3qHcUOBJW/BJx7OtpuxSTENLDHNp58gMuXOsL9Fg3
HbS4bNvoGkUeX9NeYOoJtYYTOiLE4+hvQs7TCGsV8kfSk6s88WIGFSIPf1QVAYPY4ROEs39HfFEg
2rgMPVjl/+UJDRAhYuoF/pp5QyQLAcX2s7PHobMfEHrOJCLmTdkumTk88x4TH05DshgN/qJMj3Fa
jr1036g8wlk21PlZrhZhBAO448FrNAlszJk733sUqq9lJE6Zel3BWslX9EQnIVGsyKzYtcEl5PY+
826N4DsEwd+71U7NN2AUxRwtroWA8S8SQnehwYv9O15Mz+JWaDMnKpMNsFEwfYksUeckETq4dRws
AzOsy8A6inHu5jpKgI2vKcuMp0b9QKJ3EvTA5Y9kUFHILszPjck8xg7vNAVu854286Ml5LxjxTUH
N/B542Kxs04zp2mQ5XnizYIYw2NB0X3/UHW+mTSqI22pOFE/AenuLPaCOozuNPdN/P9hGQfLjDYb
qJh1LySc8+LBB9e8L5dNOSzwrJ8DL2svbyDPPs2gKsJR+uK71BSSp1vLKo019cJMKgxxYHPImH3x
iUcSkt5ZAP1DFyKLiUtdEFtlT86vx1iOcg/yUjiirGCqh+hTueQSW12cjy73JDt7MjDnFqVGam0R
nFtGkxvVsEKVC2irBEiCislyuVMQH/OhsODqxUftHF1z0vjyMIJtwU83+c6ojx81vn3Dq8sRHylC
+e49c6N2mRhMb2ZZYmEwfFc0wMU8ujvXC3THtjXYzFCTv8od64fWNJFS7BLkiEM7JJHycVFVwusI
ugQAQLhxJYeSKuFD09hYWHtorLChozsMwVx6PUicw+VmXrvA+naRDHG93Z50UmP/cMVxzqJwoOUz
wTghtcy34M8W9fg7sgXRW0m4vggSz+QfH59Ct7rQE97UKuDc7RBCaNY2CrMrOqJSIEnYWO1GedVT
kFVBadyzGEIuB/f+9W9SWgQTSD+Gq/u6TxJ/RG9KfVsznTHtenthMHmNhD7SJfuLytJxWiaGewBP
yyNMvL6O+3qpuu+tkYxcKyXoMFOxtRYehXgyfCAQON7vmU1ndxp4KlBtjxhv1eFSZKF0MJ6QZhS6
Xk6oU1uRVnv8FiGlWlCFwVtslCncW/m71+Jl0azKghRkA2/+STG9A2bTLLX9W5vfHwZoTfWP4jLa
2Kql7a8hSvARCyWQdkGwxtNiBXrRd2zIOdR7gbVTT4dPqQ0+PJC6RCYIkXzXCq4hiyU4fa0XJiSZ
ryRuSBg/pitLGKZLbr8Mlwd3DKOc66JN5suV5PgyDwvrw82k4OcaelERkOrDuFHAcxGbur7TX4KW
QlvMfgEEthnawuWRiJIOEzarG9SHgcZiPnq82ieNPl/GWUQfu/RczDoEPVDiksi2C4IpmCs9YXDH
LOLL2LBy5FpYEKsWJYWPa+er9T5SawbDgZUp0VPuwVa3irQCYkdByaqIWRiQUkhYP8WpLzMLEZ5g
IY8hTMlrDISFEVl0NVPpMJ1+L8IQqFM0FzUkE6cEpG6ffWGn2JV03itH5nb/OmL9Cb1DIhbxWBpw
rvuBI12Cw7wvSWVMCl2ktjSKzdNtnpp//m+87F3kpHePAmgQ+o9lp/j+0jWk9Mu2NVslkWUGMO1Q
eEnbhO9UgZ0vtl5TymDw0ZBq+/QuovkRlmzczueVxNB2cg9WZMl8DRMqsBi06cwJvCqGgZ2ySStm
Vtnb/WOVRXBCOUyPFHYhP35D2ZNsYYJ28mSaoHIbm37OvoZtPuym+rm6h/zFb1D2UstnSAuma19E
hAvcuQwdW+IZxu449BHVe+oVpGv4Tv6bs+WX400MWAgBH05SD5jcxBKqU7s3gnjl0fVNwzLVp7vL
cakGqiv6k0tZelfhyk7VqV6TgqmJ4ZxFfKR244PZptt7+JjvvlzAD8evrzPP7qk6B22mZPpSvwXY
BntMGNiOJaYw3Zga2AFLWEXMHh2T1+xtQlMP5JQeiH/99DvaW9Z8OURKm095H8WAQTtb+oxBruEU
QzARgd4X5g/Pjrwk1aAUqyzp1Fi+GGpxGC/ITz6nM/i9j850NiBIoo8AF2M+5mLjGC17reInsK9t
LecYwlT8gcLAxkqMfHOUWPpcIpZFusIY11LAP3Ksg9qHf1h6jH41GsQvIM9zwv9n33GdZ0HvBGYW
MFH1nBSagXSTZVLkVJn/8jFlFuMxZ3aelr/G1/O94wcxj4YGZVuwDtiO8C0eZ/mP/EJaTDfsdLpA
r2q7LasrsH6qjqwq6RxvLMQ7NI8IC/RewpqUOCnrB7w6mVws+nPPxKWAkoQEFA8dHSlaVuvcKWK/
FwIF9tgc4A60VL/kaX9vHGBu9gfR5aJfi9FJHYR3atUwKK+f3t3t4ADMNvVpfxlSuzepmt9bgUni
GV3H1+eB5tu8K4UtvuIIZC/aLnp5sA+fJpI4faM+EYRjoCb/JNmVxwlGpBI/EMWhHbUPo4A/Mkcr
uB4d/k2PBme7YS6ZxD7y1fGY/++JHCDBGPDKH3KTKmL2jI+9NF08YcUhhHbwUzQiaWmzEBC8ZaHY
Yea9Vf+zGCQwUgvF5533gaeIfur9p+PQI6GAZT8USxVKtL/eo1jPpcJYO1JIDVp9gm9VpqgXyhpu
vihwVD3yZiJzmjamzg3Afm8Gf9g5xz+H6BAHTUChcK27W1xiHmRQDenUFdhiMJAj5nPkEmls2Ae1
ahn5V1CHXGRTLSSHC7WwRuOkgiqbTRKL9hbgirr2/ZxKZR3fa6IJBJXkYdBbgJkhJA1F0/5FRgpK
YNCFFOfW8jDbyxWbPDkPWrc60Ri4Vep8uiA5QYI/umrGsv5fWGj9dUngnZCFaoogwowZ+P+Cc3A3
l89aws9UKs8dhcDSao6YDk/uJSAOfmWUe8U8gSQHR+5ZVcTvaLe5MeGFXZ2X5UQLiTuApYIYbZ24
kFf3KprPiW5/5njl7i4U08FvYhh5P3QzSZ9ke9i7f3oPGVEAE4BZcvUl9tk8p3jpv1xYN5jbtej9
VXu9eRZl6mXYJannva+28EUAqCbwZYt+KqKgH2dUkThsgTTCV1W+0nPPNGyksAMGTB7ZOmwfbMaN
0s7YVaas9t05Dm8IONqVDLp4XVAHPxTA9NlPq+9EGjP6ywOMoK2kK2xGtmFWbr5MdnpKCTsfOQEw
HE6hvrVhxsJRkcJl9cNuXD0YTFj4SW0wt6S0MoZL+CyeDOQBHVk96pFc0WSTnuOqUcOpToB0fnwN
JY9PwNY+nbUe9s7e5PGx8kauMXvwEFc+DZ8XogAHrYFfy+bVz/9eD6QAUQ1cu7+Sof1SZKhBGQqV
P1saL7bROJ3oi1rTncHdGMWinG0ucm0HcdzswmCuxd1v1SSvNekPmcoBnEQqW2L1y5/RekA2QZyZ
BADczkXudReQ7+a0ptoggdWo2T9/WK1ZRQJUw4rG4DHm3Zk+U+mRRn8P5qYedgv13mC7EtFW6gCW
rWh3aAMez3mlHO034M4xg46aSdGI5ZrTMyCnJ1SWoWgJB5OcqEZHz6X4uJ+Yu6uz2HfWSUf9KMcu
K8w1YWTOse2JbBowJZkvIkB4asLvh0KgqeoguKOnlWf/+i9NAHRXQIiLYJgJc1iQwtg2HBl8WmL0
h7sHpxOU73/q40PXFyk/pS+I08pvpiEFBskM9oa3M9rjgp6dN267RQThRieg64GI6iWVbOr2xb/7
au1oSiuytjwxji/b+rSFs3aGPlVBbVvWKVULKzesOhfz+wFvLpVZSnuBCfhTeThfO/vn8aFSBMAq
qv3mEq1fCpzHJ1rtKknR3Sfm4wbxf2v+OKM8mUpGQVP7odr7OsEQADJQUPosYVdjrGkh3zqL6yBs
d68paT9/bkg4hewcAGASz1FiDLIbp00FKOlA5QYFZ6vnHz9ZmZJ6/gbI4OhlY1D1mKc/OQ6hj3tm
f8P6B1jNt/TaRuvkGcuNxsGinv0vseuJrm78w5m8I6Ma71BCmL0S6O0GvmlZTBMlP7J/zHuGNDcI
YjgCBv/1H/5Gvz0U6T8KXo7YgOkMLO7iIzivoap5Z44Jn5VzUmxQiQ8l+0KeHGh+L3dt5zycqOj7
GeuUHl1vUCfFeHFqFeUC7BGzy4ALUc4g23WjGBw3Q496PEZXc7+m8Hf2DEk3Rl7zJfC+0YG+ON8Z
6Ks+8yxTL4aTEzWrpwypSnV+FJX0n28GvV8nFIcjK6HC8J8xFKFQPMxsAkcC6KvzFls1KLNdjYLP
qr4hXza8spJzDvT/aNxxzvMahu5IxBg2KtJc2MoEplNcdmFxlG3awCbteINkDJTRczLBNZUsWByr
qlGFhwIDY8eqnpd+8y4xUZsGWxhDm3V3/2QLhyImm93PlS3FOlIXPkEeqKvjitlGAbqvTm3ETYmT
mBN02v7EtP3/jwNOFqc6KjRQOunn5xfBZfmmFcaLME9i0BNJFTDwaFsAmYSJhYnPuDk7ldkoAPv3
yNfC7qTOZKKHRxH88o0cYkIntTRBrqKAizPKzZ4Jmo3M4wkxsqjVhfN88KS9lyc+XcWUkIlnOKys
LB4duRpEYSE4TLZAmZTUJ/YUrXpQLv/kTjoZTRdy0TzUh8kyvDw5tW8Y3Sp7Eb6B/zfiHISdNr/P
tPVpwFyk7UWeuQVGT2j141VFfrJh5ERtjOtA/DLXPZ+79n+7oC7foaYIYQTB/3SnLV1E3aq2saje
dWbhAXeubcICfytE1rGNlq+zGyIkYnAhF/+s5lch0Rn8G2UF/WCGE5zejWx4p4fip3cmZA8V9P2X
zuxJMRkmDoQ8yi8kd9hAMV/80YJcCfsoHpUS83kWHN97Ljw113usjMEeueyHfrTpNfoE6Xoqvbuy
RBMN9thij1ckgWmvxJCVN0mnZ4PwI42vPXR3Vt19izz+AjjpfiG1lJ8qMLAeJU2z44MOzeRcvBoN
6yoEI7VYKQl0sgq9/2Ur8ItPV+9r5nxBUF1OyNipENPx4FuNNDBFgausIhZ4vzOUfwKr6hjTXRr+
77yhHU+E4b6OHhKEiTtrWuEd5LrIaPitk/Wl93qy2gqNdnjBdmCzW74zK2Ha+CEM67lEGgchg9gl
PdFZH/Gh1AL3waZvSNzcQ55Ofi3kNRiwMB9Rw6H0G/QnJPq74StITIyuh31fytPDr7Lb18vhys9Y
yRwCRjkwAVjBOtL8VW2nh3FoSwqJL8T3DYfvBHgu7nc659U0wbl+uGDmEiMCaWYONwppX3jLJfX1
DUHFrZCPV3axfO6gQ/g4vxNK1njHEKQAFjpjnINVpqKOoNd0+DmLm/C2DvS66nEz2BRXqOpRo679
5art5IJlq3ZsGgjQRVdC7TU9VzKrmKyMHehwHrzy1dhA2c15du15t4tvYOu67iNDRGm9jUwLsaYc
FmImnPYRDAFh2QKwYwCesarlTYtxfl687y8gewh1XHENVuutTtLgdOcoqR3oORA1f1x+JCWXCsfO
VHI7+VYZUSTvK+q9KIwnzrMnA6kjfH426/I9f5F2WgutvkA6t4E9I3VIDnG4ejSNmv67CdKqc9sD
ImHMYGCRHdrbjiO1KLTtbbjSeWYlTooM81qRlvzwVfiC9N0q64aE9yQlZwFi45WWTTzqVmEDxM6V
k/n6TVaxm+5opmw2RjfrvT9IT6plkMgppQHwOmv7Jmbw/LNCXzNcaB+RqqYZXJb8gVR3C20qzqOA
GZFsXk6VMyK8z3uz8YdcJJGELCaB4fYWEYrM6AMfZImpJaf1p51VtpF25bcHCe2fzXzI8i36o7LA
thX8XkBKEpCx3xZ8+bRvD72Gc0I0C79zSNPnhm1DGOofCZLJp0wt7MtzkmYIfOlueCStkThGopPw
BpVaY7lOXOKBuspCrBolu8USbQJt1TNTwbHGQRWwlKQ+vlMXzsFftKaJnhCQrwhrg7atJhsbcVN7
mPJKTFIoaDdTmmyCqrPf5vlPz+ebg7BlvKB6MrFn3B9wVmEALmiEOGkGi0wMkpCZuc/y+m58v1Yw
6JudeNlWBQdFgSOZ+e1sG6azt7MNd66SfBZyDXEdIR8S01RctR3bBtbwxqq7+/Fk2DUKx7jzdTwZ
vTQkOpGWEdQwfreZYNKvodgxSPNzSfZJ0rMxOS71rcPrFMDc3h5+flUEezFS4jhGHTk+ryEC2xVj
oBivDBTa/ZoP2bIh/0Oo/C9/TP+6jhV9yeAU2+oqco6ZZyBaDCoIyrOaKvRhE/AQyyDy0VRvwfX2
MNuQFDHrZVlh6J1A/L7BpXgqgKsjcHzpCZsAplS7HwUAUlmsLXak4MOM/BJz0oLqpv4PRsIb+PX7
WT+wEhXjEC8CZEhw3WdFv7LqAWjx0XMhHS/nPcDGWrtcsfVrMl2+95zNoq1ssrrPSo2H8XABiLfa
Jy0LuEnF13sbZkkhuQY3y14HZZh9P4KVF0b4T7YDTZJcKy6P6OzIa/lG3dPy7xTLazeCMMUL+7fi
g6kRgSmmoiCu248HnanzFBTqgPRX4sjKPZ2H49SkCwK7YhswWXndtFUBB8tVgfRSYgnwW4YKz2ab
DpBiGqBos+cgAGg6xZCF/GfKKBDrzUx1B/UTyw/+1VRKTBIjc4A7sENihBT5Oh/3xvG9Xb3A9NxC
QnqfsXEYSIuRjW8uitWK+cZXs3SwEG5gvXmE6CMcILU3xuSRLO3s+0D+WDLLxwb9XUMZ3WJI2oWy
G6OntuzP9N2HISOm0Bsg7+HfLoXBVPUe9fS3YTlWfyi/y5vt2rePo8jc0r29E/06Svm/5RvNDexa
sfgvGsXFdSOgi7P/zwbhTHkN1NtjH1eJ1MVOzz67xg4xCdRH9KrqEho3ePON8uLF57p0ZaCf0OEp
sefLGgv5Bl/LrTzUocjR4W2bPWtjS1pJXKEDhxnRb2iORrfmWmJyKH0p3YX2vLQ/WDWO0iG2oaLt
TbgQMaBguVdvjkLVBNzPKxB+NP6lips4xDIvAxaKVWVAb9G3AJWddukC2TEwc1CSc7u0iFIPDYCE
rEr7KybP+ukDA3K9imhss6iZEawISa46ymMkiz47RbaVPermPuASgQd6KHpQAm8o/y+bECpS6+mv
7tNQHVsO3VL42JwUho46V9tAAB4/VhOlZhIFGcDcxQolSwtP12JbdWsU9jFn8uohRxJEpsA/dvbv
Q4RvBcjnPih6wZANMLoKCcMzVNyibdJ/i5RY52/JYTMijSrArFZG+O232h9/Gfr5ABmhCmcJw0If
bQLT2jD3Q/zESh3gWiirMH1C51979mjOhWAZjrE4G4wuLbk+czZkaRKg2uyXmn39DDmj8MyDf0ov
zpaViblr7pEjRKKrUhSR2r7lH9dFYg+9c6bradRipWD8cLqDQ3nPAc0VJASQe1BhG7DrBPnDwwOU
niTKv1NF8sLbnxzF7xWVHAXAlHDcfvyxDXLt24TzPigEcUp8wlrdrvg2wqXcUc1Mv34+NvchBjvJ
nVIVOx55bXd1Rkp4yEjUQUNYRn8LBN4CCh/3WoCDpjaLt7bNLyqpx2q5qfBf+JpWuJTuzJJJZ7AG
jhEOoaC9OxYxJqvuoLG6XLsgsvMfO9lUkjCCvQEmnIKpxHVffiocV+Honx4bQ/zqXmFMD7s95jJ3
eF3ZqM6oTzaGUpYhhVDD33hPK2bT1aEel/JpH+178pV3s02cdB3y1E5JoNSROD2U+xS/GFvr04E5
6nfY8aMu/Yd6KEksBsFzf9MiZe8nw/3WAJYL9kJZJy7WMqBOSmMvA1r1JFgdxgmD3xuduCB+mzVm
cfNPEsRH6M02r5Nz7NivaT47+0HptTzHQXWqlNbVD9QapnbjVONBMIBDu/2jrBFUD3yUDa4SLOQr
ioK6VBoTksBcmfmp5BahlPgQ4oRnYvJEZ3OCf8zQZ6ANBBAA3a+GK62/TGhSvSNHy49f52Y+3ls9
H6pUDmy/s8tRmKZ4CDfYJqvLLchUOBh/OygS2A5cXrbs7u3ioglI+aNs99ZDXYQw2SnnHM/NE8pq
v27vIEodovvqxgza1EHroGRh0lJpybwXlUZ9hCOGSzvjg5ZYPJ4oKi5xodGwGca8oa+QadaKhYAq
+5EYHpiIY87ZJxwd93IFhBHcS5Lu1tLzCSI/ZLJrFcC8pcSY+xeFS0TWQV45E2AXUC/C/Ber+tDA
Nq6knmwS2HJ19/YsIYnVirdjl+Nu7bFNaxYaKxuXpmSHsvvIN/qxt06GgqT2CMXVMvmiiI9UfPSP
EdXE4lLvbxRnJC0s02tkVdlSJfyr4iHqKUQNLKYcruCnRSUDtOhcKvkFh+0hVWCv5ct/d7PTGP/v
WI4eoG9qynzOhBf6RVpc9tCZvOfPlXQkFHKZIzBmocFc4gaVW4GpNZRuUXHdI2K2XUDJRxqZutt7
Q7z26jmEavDhstDSnqSTreh/EYuOdLa31WehS+AUJRcpLF/BGz5vZ/e2hORgk+sBioPtJsjS7srS
24jUZDcUvxHlr7wPXuVsSA5P8ohLccPBHtpy5/CnyuUnIqODGNFt430SScux47F8OGJmyhn34Qis
NPbkraqm6pDWKSB/5DkZA/eRTSGWkjZMwFRYKK5eztQghkS0GT0VXacuIHf5JKwqb6HEVSAvT+sI
9U1/CENiX2ODkm16pxr4uf7scAi5eMvFQ76ZR1AXu57kP8rC3AgTwZ7q6/MAy6UWiY7LXa599uVw
0cXb/tSbZzBW6kaLREnv7NW1Q1ljmg2EtqAyJ2p5pCK2pXf0VUVzoS6AOvt5r2rKIuJm+XEJ3N6N
hNldqdB5l+YXx+9HleQwyueItqptyVMiQws0O63Kcb7FJQX/8BlLBCemyZI4x5twadyKYiYylTK3
Yscib2LkrIj6FNETuyjaB9i+FLZbz9rcE/4zNeBz4JLiyiXab96cEO5F55w9xjNYzHDDrGn6Wg/O
CLJ1W0hRnS3RNWvN3lj4GljC/MN7tFHhzxpyCnR3+GUrUwD0MNfogykccyboggjhQhIxKI18eyua
dsOiGx0mcH9LbCet6FF4VkxDMAKhR6M3MYy4LbfFe93F67OdnNxgUBMlQjM6jtuoi+So6Zmg7JA8
Qm+PPAhRfpLv1HdN+AqIVWVxoX50nJ4m9zZk8aQjA4zDbPZcDx7olVhtFa+ydYmuzcmEe+v82AtP
4ZGrLjZlVR/66SbqiPNxU8OPkhUEI2JL8NEvJDlcxxMv+Uyrdv+4rJ7hXnoj72rYlEyOCkVx56DI
9fVGMcOLLAcgaWGcoqqhr1sQkdWOlfuMtRy5bPMFDUqqCYyp1yM6evXYVboDD01ktRgTz4O1YQ+w
FjVMW8uthJEKGObniR74q5rulIIgPbMW4w/d/sBUK99WcZhEYXAs0BjanqWEEYd1hA7H32iEYj/E
1SUgOUK80mDF44QyoL1sN5FUgIM0fOwnRzO4LAWPInREgr6ozFRYahghs5VHfyxVKDvIYyDoywW+
KM7XqpvvGa0RcNHO9cl7/pFlkfbT3JOOJpwGrors/zieZ4sWpEzxa03Xez/kVYfd8eKSHuh6eWHH
84dAiq1JH8ct04L3eOSD4BCgqcLXNcjkMQUP4Rx2Q3zGKhKK6KHHXWtxoWCqhHDfM8lu+mcPYb8T
ovuzFaN41RWzXecDDPfwqRZujrsaVEfIOIdnT0nGHYzrL7DF59Bum6HMD30TBPwxIXI/hLgf1nll
FhFNXdFukGTnJQvp204tr8xhy403oNVN/+3LUW12LkbkxC47tQ2nsr0pmk+kBMz6xQ3hzsNVao+c
7TZwXpTV+RGGNmjKZ3FqLrhWKrvxHAFbKGo3kaxtDtbhz/qXc6n/CcmSmKEVOi6AZc8t3sRDLJWn
0HDPUTY7jpSS7HBit1a7LSOsQhdrFhE+3I/hRPse9wFs/Kn+pCYktA/x3y1q1k1Fjyl+JMt1vb27
h9uItkDPn8jTIMuOpS8ZSqt9mJU0/8trmk4l+G0aF4+J+2CcIXX4xJ1MArNCRtAWo4DmTFtowtoG
kgvIRtFe7hJ5YPsQG/fsaGtA4HT/MZ/jHNPqNC2ANmv2iJ0bv4jaBynX+I+UtpuR3oc6f/klrOZe
srV4ZDxONgpq/XMrfoFgcOGTVfPaeEe9hJ8tdiIuHEFW9soZ8WO5YkjMMU2Pg7T1BrnQrJTHOiZz
MLAeXWnYjudArBRMDHsv7d9FJTxKMn1sOYU3LWzz909ojYIs74MmohnacQ1r9610tbeVd3uTtA6t
Q5pHbXLKioJIB68Jcm2bnU0Kn5ITXzSDTvo4SO47CHdnCdIm31/haXA1qYBM1Xbo3/SWnJogMLVN
VkQKP9yuopFn7A6P6+ce5pq7yCALviDIcwgEUHptK6XlGQ4/O6GkNGzS0CyvN1ibpxoOaPzrbBdM
ytY65p1qpwHsJzI7FSKqI7knc1WGfOvhipSWn7GgUGoEgAFbcgeYXu5Ie8OlFk9FynHQHW+WX04l
jJfP39pC1R1lrk+iMEQwEqmBvfyZ4I4XpO+F/GneRxWuiSXKhDet74HlyRBD4hNwCAUzIL0XGfAN
+Chn3ShWd8GeBXhN/Gd0pHV5iZJcCCwSPupEU7rMfLExHFRjUnf8T7zgg1B/Pe9e+/dqNRrMtj5T
jDqcDAD7168HmnliwqprLkrulQ9iXRFqtOXCTQZcm5GC13x41K0yxCebJG7qbeM7wxZFgTsB50aD
zn0PnHs91fUcywT2tAqNFcmxv/dls2LZ0fm063iRFuCPEcvKDHh04Sztl4WxNbROdQcoMM8QjU3I
59VDqSvFX/qTvNOo4K/UcXL/jJFXAEx655rEiddfE303OD/Gcj1bvZWmBZ8TtOfe5hi8k3L6/OA8
kHdNp5JgIxo5ZsYOykC+ZxUkP41PxT27fSxZLHaAfP7oA8x5nS7NMpQKF6lAg/TV034Rn2NluM2E
1KhXs+Apb6OgCT0hPuPZbvVqj7pRC353cSrdHPmwhrNKaB7a2T2KQjCG4rr5Hn9EiY9/2pnpxW15
/upYhpE4r56VvdbPCx3ogK51PGB2ygftFTv65hyjnM3yau9kgkNwkKPfDuolph7z7RLKMSu5z/Yl
F0awtMk2VT/owPyAcE2wMNFUO8q4ohWkm/a3P3rRrO48iGsVp259kQDFH8BPzLgcloNAid618D5Q
G21SCht77kGjPfyn9qzyy2tLQxzzBpZkIqJHsxtHEMlBmoh7DjxpuL9sTPw6e+x9ZeeYwTr95tl8
eSxm89/iUnJMcoZGPCX9n0sW2cZgMmUH9wQ6vkk1JPc057ryJZ5m9++XqwyMxtHR8AkBpXpplgfp
g4EsyTN2+sOAas6tdSup9zQVtKh+F2x+VnnwrZUocWXLcu0DQBbyXFdlMXOwwGXoR0BOMkjh+pLg
vlStQvWkkEcsQPYeeiTlvwXwNt+xgbPPOvbcuLbOARSF2fL8gQFL4yCbDUTJj4veV0Iro6/E1Av8
SAAu/jrWASSHtOHyv03ZBqxU+zteBLvEoNH9ufRs248dwGZyhOCTtNfAURf1kHPb2r+8satmy3s7
2sivVG/ci12YFpMa7CudoJcnRgG4l5gcRBQUe08mSoAIM7hdUCr1C5K9I6l+k0nqd8LsNCX5R6VA
nSTIuAM/jgiZnk6iodgSdlFOPijgUo4S9Fsm8BLrD8Pufsg/VoOJ04J1C7EhIxVgsj5BbVcsjLZG
QS/K36uBVRHvVMJKUVps7Ersx8Bn7pkm0Ir8Uuy7KBq0klw4MxEhxQU5hpO4Qo5HsJw44DC2SJbU
8OS2athi40hfgDub0sEbn6heysbxeXKTu+ch+9Fwisnhavqm3otu7mXUXnTPznrwgjRO6wNPmH5l
WPPIq8ejb/8V+Ma0xXwOSubm/swsY39gAODHNUAGxp1oXrD5Pu0YiQ0sBbk8JZ+mUIzP3HMF7i6i
OWcLEzGgUQtFtBXEfRhBiFwTTL+XxHbXRIlKobCVSXJwyQ9OmITCxmdqmdjPmOz3fciYVEf3RY6W
FCWGiHVid3rWieRzoB4UWHzodNht1UuXTh4scjqFgRVUTerBD5/6gfe61/152gzL2M3X9QXeBkmW
jXpVEnZ/VXdWidCTzzAorTU5TxJSrszKGCLrcqULh8uNWGNlcs92HwR7sOEM3Obji+YyKmxAzHMc
UeS7dv4vHYpiJEiwGXHfO6/CaoWX6pUdDqxkd8tLswKric67E3RJz0D0iOVSebzazElXRNMmQEMF
qxo2zG+1nlEG04ukALffrb68BJpYgT/wLq1hqbycKCcjWBUvPVJ6YJLe69JNBZ+msXftK68ZT7fA
zRcUlXLyUAdcCO3c+i6iic3kGRrKQWdUqCzChlN/JwVN1LmFMfhQlFXiwFf6+c0T8HMcsddVR5I/
1Z4gnDs5ocw3wzjntSLkav66EZ5KgoeJq7z+yWn8tLE+Ozp0sq3In9gZYP8PnpJ3qgzc0CeTZ3oY
uO8AUkL/AKd5p5q4uxqQqLqvUCq4+noW/nr7gYPCP506dTuK5ylc4AbqYax3ZDDyUs0keoOF3Oqh
O099Dq5dw+95uHG8wzVOgvqy2VU19R1U74HC95EXxPVSyLNO22SsmyGIG3ZzPXnBCBEA8S4N71za
JbwfguJdf7Ii26TL2Dc+xmVn4MDNpjbil4TQTpAHrpNDNioPmZXwezGVXC/8Oa4GQrZvAy6sSCIe
TtSUvjnBBscL2dX2hiHikd/fZmtHEPIbIcviS+0AUNeL4O+a9+yCsB//YVlj4kPj3uOYldKFYFlZ
8NAiibcPAYJ9lycEx+OzEAlIXReHIzg8ht9HkzwUfhZh3oQhfs5XFQVMOp9+yrTBZVLz+ePXYCrM
srrPw+k9JSvP3jtK4wiAt5QnxE6k5bFLYGrspi6IxvnVhv+PinrGE5OAhqUNiJ5butCDfiEBFhmd
/JNd083UDMiUXUxOH5KfNtOvKqosnNtjV9qV0PPX8sFlT3Bq2Ti43cwnOLqcfuMpFVwW3HVNg9u6
Mhf4CeC1Hatkd48d5J9hXmh7OE0ZfGzFbgasRok/l88ZJs9IQg6x7tllbgDR4sY0qA7Yc5Yf/FM/
rQUyzbsyUYeEHnqF8bN4JtucpLAwPq3/xckiIZi7Tik9UvHZ38uJQtnsXu8g/NVpLMZN+H9fnlQc
NOFEZo/OpLEdbI9EB9d5orcZCLPGmFFzZdgna8k6kUDoSAJivrjZoirqRMxjFd+C0SWYkUCNZ5dW
iVwIx/4078DLLM02hMpkS956EtqGY3eaytkn6pnpU+1OGtmJvCbuajVV2u56izDX0Iv+QjsVnZXT
JtBeNbjkkhp192SBKgIWm8HBL1i4MSUjgN+JQ8Gs9rYP5dPneyyYNM+D+cUUE0NKhwLOeQyDzP9S
RCzMd6yWRbFoWS5+nnH4M4LMKAd83vhxVKciwMbcbOg0i5n8WcCK2sQFTM3KFKll4TVPtxFgtVWJ
BSKmGLZ9csg92Ym4TOtJ70PZ9J9bELMeYR3JTBL1MKvqudrENyCgSYiv9bB5XKkK611AIO/SdJKT
z5Riuq+5JedKzYjL0Dffb/8NcdcP2cgEL8+BtOcVzbXprWOADo2WmtFMlqNq+eQ/yd5baU5xWzgZ
LyrQ1Q6qZW/385JcksZkWb/9ojDaeUnHtKHjBZH6NASHGvwEu91Hs3gsYagjw2UgsEfedeyaUD3p
MSS15/36uGFlVBUPbib56ViNE/wL8yZEBWyjD9wvYpfrPNdfKBFWIvKAiEPRha+SF/++jRPdidLF
irSBxTgF5zQ9CReWOl1JSu60lT9NUvUFsy//TY2pXHo+gC0wg14tG6k/l8P3I7GcRFAAhjl0RviA
WpIqecnlhmR5FVX4EYByz72fk3v1a7uehDnAT/lMXECxPOlai2SDYH1ZShytgyPwBGDb1PuVdpzo
W18C1Fp0Ju/LwBDgMY3pThu1cN+e0Z439q+7BvmMk1/aflaDsNQWXTxK0MLJo1CO4Lu1UfdTcOOe
1E+vKGRq1JfegesYtcVBLW9zSKs/t6WymPGyy6xuULWxoI/4Z3rpBFMuesTbGtAawYJnQqUwI5j2
FfCe9innVF1jYtJKkT/SFBXrxgAoJrWrP7x9YM6qTA0HhIFHcMLEWJeOYsU3EPgWvhedlDCP5q/G
0JffS2v2jflzwsa5Y9CW/zh8LV57g7jN9IBFrb2m3vAtFOY5dXKL5d1m7r+an4y9qdEU+FSpxtot
oBW166Ijdcf2cXhy/GEaqlll+mZ1b+lLR6M4c0zT0Kh8eUBrLA7Np2FYDRdY36Q8EHJiuPmkcuwT
hYl+97VEuM3jYfAqcXyoI4B9F+/mViUL7vv+MJxbfkSk0MFI0TwxiaPs7EF2o0k+A0dh7JC07Dzu
lud/YdIYPw13OjO/Pjdb8TDkd2u81sTVLIzCoZW2wjFj7mtMorgCF2UsvryOm8ktmK4vwRyFDJW/
YsmqhzfDKb0ThugboRN3B7kan0Axr1L/BOF09cVO4xU87deAtHflrThw86/3ILzX5NW4dKKheb9T
lJ5v7gfFmXxZmz9Y2f3rX0aJl3W8RdxWABLYTmsgbmHCwLNR5YycBBeLOpR0BVa/9+wSuwv4Jomu
ReUsHi948UhbQ0uNjLXWoSWYpjdu8bNTE1BrlaWxRVwb0k5JM+yeuH9zYohkV8/TtrHPUiMRi3R3
Qgr/HGbi1nDE2yrguyZA6ZcM2mxTITK3r0pWaelA63r97/FC6d+eV0Tl8xGDNWhhFdFgviVGn8GT
Gf80XbCN1xnMc5TmaBzf8s5QwAGULdXCKTXiZR4EdKkTULKsuRNn7rt/7yGxwHG7sCp1B52vouBC
R7g1NYe8AWGv6UPhtUr7asr5js0xQaMkWoY4ElRUA+gAqz9Z6KMn39NzaJw6Lo5lqmV46sN1nZi1
bLIz7Peip0vaSVAwmgiHI1lSGY1XgX9c9Dkds9C7ydp7L4ssp29hRYmlYXbwjC/DpfAoF9XXyCxB
A1hmtXnjRPG/bYak869fFRcP2NZ2vGEssHw/Zy21eE5k5t/GH9YDPBsuAuQNSwmc1snhRmYagJMp
TnKJPa0sndR9cP2y+GlcX6nN0pz8cM/gLXDtBYcvK8FyAgVkflhSFjj9NjcAPy9wyEbcu63Sw9sR
WHhVn3rld1ZbD9qhqhzqfHy0gU0L++HY391pW3qs7Db5MWSLRywrRlnXGzt/40CKSI+rMe6vnuSy
GMTf6YxvWUJ5eTevJFvT8ks+HR0E9hdsNYUfyrSGIq+hXHOKK7riigrDW5DF+TcE70cDC3lBix5D
PNuR7xUWBimU1EZZpySXHKQsnWHywrelf9sBDCfF6Pb1lVX+u0o8CTRwpXLH84ZgWZdpQLBsWqBS
EwqRfHeHf1urwPADIqt6XZiG/ETlg8btcez+QFTTuiqZ8tCgPDoq1alPntoKTLR33zAjX6q5CG1V
2GYedqUsSoCL//Z6/QTZKF34oSB/wtdwpP4cBRkvsioCQ/0SDe8CovDJCEDxDxySxOjjZcIqyGlf
tVhwoGYpgGko0XZLOtZN6poeo6hh8JEpFFPEAanG+SXRk53OZXHEVxi5w5cKoU/PvDt2bFbCE2Zy
Jkja0+nkv3MkZ2VYAgf90X8zNjwZmtGo/F9hij9yKJJvd6LbN1eLDvvr/PxAoCLT8Dx5ueJfhsyo
mvQ1VEWCrhsDt8xv2N2eT/zH8eW5rySzdIMW1VTQelgdzUK8nO5kFNq3gKKHNRh48UcGC3UHKpRJ
793S1+aSpZCeLEFyGww5rIS2uo09vawqhTY7SBNk1A64bM8MT1XQFa/Gt6t5OxD0qP1Xxaup/h4y
IWukSpn5VtoQV28YzahEZAhgSstgcSJA0+Mmo0AFoFQq0q1cj8EC9Y+Avkcf/1TunQwm3GFKIu5e
TotVgUUNkg3Hn2uDHY0nRCvh7HZcoc0Vmi12cHTAZfqoUmEmJ8n0NuMx7f3oGxm7tJPfQjNnh1LF
8oympxp1ej4FilXp7meWG4IF3YPn6NIG/V8e0ZGLtK7vcD9PMTEsEON6QxZWbFrDT5UfK/6lqgzv
oSJnwT3gIiXeqYgBI2kC1eVPXEB/u4mE69Gl8twIj+8zkmSKZtx/nugfwdyNvmTvxBqnG/VwFn4n
yDNluuiBo08NxXphrj0LaupgbJ0is5GFlJFue55HY9oC4pp0rbOFCdqKfKYuxhxLoJEDjO15aHbU
hOlOaTeQuWAC3QleVDMcYZQxBbqQIX0wdKlnnNI3M4JsR301H4bThaS+t7U09eVv54LvUMUd0uoV
eu5MstQKHAq40tZnCkSeRJMgULRiiqviOf7Kto9tI6dNkfflXbJkwkF8r+M+JudiMZ0VKxhLJeiG
W0YsfM+U7FRgktREMqq1FersZB5Lkxr7IcZoPg7l8gU4lC+cL+e3vat5jJHZGKfGuYcZ2Gmlpldo
diwXyb04gryTtb75WYeVbMNagrgC1IlBYGozan7vkEoSqMvvA2Fe3d4ypWX5ieArUy2z3TxCKAMi
KXqSWnEdDozyUYnJD8HGqe20BWgoqMiPgrUVlZUEcncRcCOYWe1YvX5+l21DnqAdaR35p3B6LMSa
8hJNSQWQzLdwXcNH5EZ9sNBYdz3pJw8xkdebsx29bB3OUzXckYh2+CfNv4MxA7MUru0rUzj4AA43
6tkhQenbJKYaTFlVnhVKS8Lb6tXQ5KwxwHR8Zl4SeroHbXc8Ld00xv1SBoL4f3P0jjL/yMoPYAd5
rg2/NjrUNWv6UmcBgqxpSYtkyvTV5fSIGhWiLeQZ/TwQ596bPx5dOy3hRk811ByqzNYKq/n2dOHr
7aZbZHEZ8o2GTeM7On/gLc7KpQ6fvFB6zgIpUu9f4/nCFrbaZ4+ZF++R02/6AIccQYEHE6hTIXBm
Wo6TjcotBlSs+2maHljTbAZflnhT4f79p+2A8qkpEVune9/2K065m+RSjZHn84uYpoXg6E9s7vOL
AyBlKBg6J/yTGEkyAx36/Cv4xO5xyDlxzzzemHeutvDRnhylZ1cy8TgonCpg3RI4tfIwJFuES9DP
eGLc6FOYDryQ5ORgDivEaKgoW1cvxLuoCYLko+aQM8VyLEPjdT5e3nSZqPyH58ml9R/xsCqPByB+
phtPEMTsq6EXVmkBWbTXgFjgB51FHYLJp6MFmwcKKcAYMZ0Gjoft3biGIoQEzYuBjn5s1iSNHGiM
mGWLF/GftMhdZ6GWmVY5LKy6t/muQzpqzzCP1l07Ucp073kfXaLYU5UMG9fyzo7Mr5yVgORTQcjN
MGXUcnhUetmCGHlAxQitt1jszMXme54834rtO/qQfmsD2ABR0LqrgrbRMiOGL8JfH/iegYm3W50z
QGB9DWdc3Qu4sg+MBZ/ccsi+zN2NOXI+O+iCpUYLPGTxttEFoYXXI/n5dAB/ZVJKySJ4IBSKH479
9LHPH/ZO6zsY9iDF6ypr31yZXW+JlatgaoBqsGnCZa9vN0bWawttgpNWlE9ZAceP4oKjalfbCbrc
zHeYxocQrpcL3oiqAvpqnouLKHpqzzPLDM018JkzKvuumAm740lgjJVjKxy6rQfC25qp3Vv8rH9T
KlgaeO5ADWFaZuFNdZXfzRBGoMRqjYpKZA6hGWymwQQoFrMpof+LpDP2EN1Q5X4syJHI+UHqY/j9
6uAP6kn6Fn51Qc7lWI/GbWcC3R8+8PUYypKlmbvRZfaX12+OD2jnNVZmZ6w3lrMOvuhzcOcnAv7D
+v6xfn67WtYiXL7oFmUNNPKIGRFO0K0urmIaaNIe7y96ylpz/MVcXjUQnaiF3DXJkNk3VfQlp4U6
MoQGZsnIV/PvTLxHpAAF9lJQ9BZCTZYCt/KO9RPfmxPHIxVL5zKLQo8prV+llCZG308kJHmZQFBo
X2Dy+yMkLiSRjLm4ahMlfz7WpriFcr6p11UCGvSWEItT3NQhB1OJ8oBadCBcwFhrO9+veBQHRa2l
bHsrioIYA44RS8OZq0EL80rGfVQ9IzcbMGminNnVsV9x0j+w75xuEDEfTsVISaQ21rk4o420xWjq
pTtUqJGp55jt1F5utBztEU5z/Ie5nfOZLlv7FlRlrtencVgEDEGaY2hb+c4HTGQmvuL3hQm9dfhl
qbdmpHgff0SSEpdjR1F7ZDhJoXR6cTCLPrY4RY6QOOjJWd5AX3cD31q3NDKeqcNSNdlHSnIvf3mx
1mXsS1Y2e7bivGqcFJZU4gBA27pX/oeirSYeYB568+IKZvUJS0mfJBri8cvn61p+JXyUvQj17JAQ
pDJQDlKINgcpHE5NYWU5Le62iKEeupf/tVny8RKyix2Mkt5DStyOgCJ+NoTgtjAQ5eDKI2R5VYPM
1uerXFbg/XQ2N2FkCvHS8mNyNutGjHvpYZVIc67eUS6hNZfMxi7Uo+u96pYK6eRlXg13yzwMVSdJ
+vpprwIilTgGyLKaod35+/f4t+bricinv+JWH722/CgYPD4FClPQaOSoIMV/Bkren8WjW+tYO5yH
wLfNSSfk+HuhFajNSfRVTej/WvJohgnBNyXPU+ynBIhr05+rCXIAnIKX7dwRuDsxMjaSXRtNyY0S
fsU8ZAs3Zj9jdBNQ9LzckC4OjzMv12mxbOaQkQGYjfSWpDD3chw4jcOPqs3aAp9atFlTZRfFrv+G
vCC/cqnxzOa/xBN3Cw1tRuqUrdTVbgVT3Z5WzpxYu50MkrkU+I+jp3vUp8yWHd6a6n88Nn6DjuGI
ZJwEVkIUzulg02DPuZwP9Oh3t3kCXHw8smz+PNwGrCrpzUgBn5RZNyeOQgdXeEpiBGAZD6K7CNEp
IIu/usAA0oGNYX3pZLY+jbSXxQh2wR43hnOl6+Gr6uK4L3cKm9Tle2PPIC5YdZpS+lmfK1mKg3eN
O3SoIhO55dvsajAXu0NtFA5YfIYvm4Jk4taRIkuJOyO4rag67vOMBxXfy/r9EKFNMftJXnpEwcXC
H3JQdrpjrTZMYMzhPxYAMXrzI44LCuSR7W/kZeDuTL3OePQPDwBYlLlp4AQ2cqpyfMWykDVAKuJz
yfNizI75piWFNMJ+rRTBx2Z27jkQW9HsEFx+aQ5reushB1m80bGk3E8LenzzbvYD4WX46oo7y0Tw
S/Av2ADd9IRHvaG2Kxklh6VPK1FyjIhF84C7hvIA36+MHBbRa53qeFLRgLc7bZ8bAnfrYFDVcIIH
L/2UzMphIwFGSiqynMatSVYvABDWCB4M3vp+p5ujibr1A+nJjxq5hejWM+2Ln8EjQzace91NQr7f
gBmas3jXDUDZR40/6Y5nmPz6bQc2+O6qJQFahM5F55a5p23H+txzA5suI8SMNP1vsnIACRHGcn/O
bMbceIUAjxrDm9YuSk3ktpF2qFj3+8gpeY6TfvKP8DgzSwFKKR3QcVtw2MTXIg0zGsZcQsrwRpum
Gp7Wf6IEM0IVhx2BN/heh6Q6azr5z4OHGdQ72s63LvsDM6QRvWUqYsyTLkyIuiklNYzHHP+dI/u2
7F5nbS2zAXMC0AVX+MBS8G3S3bVi+mUunTbxMkNu3Hk1c8hzlSOUnFiJ4lJTqHtMRsFlbEBaOXI7
xcUsKnFF4e4+dnTZtA4xIt6hmd73ydukSKOkNK8sWud/LEzO4TAg0dnxHq/xmy80WSRWK50ey5hx
ETDFAxw3A9bUMfwU6vKAhFhghFml9xewlxqwJ4ypNoUb1BeU8Mn/gwpbV4TBCnc/J3l1Zyc1dcG9
Jje1ZTs95eiSLlLKY2Z7/XdNhK/fbsrsfElBHBK6Jh4iQ9MMRu4jddy5jvedlNUKE1NFy3vIURfN
Fw141jh2/F9r2zFlUlEfTNut+NwERTWKqQZwVE2I7bKY7MNtx7kb4kW5U29+4Fcu3rzFTsU1Ksn8
/G0J3TBVoYMm5bWCxf2NXuoAz+0Qqk8xnJ/pFg6yng8Z/b74s/Cwurek8K88qKNy/okjVcVRvzE2
lsC0AtBBw69Jt+ilqu+yV1oSb/s0LAZ/M5Jb4hCeHrNMnT3xvDdFtqDply2h5UrA55dXkoVglqfh
97OWygUo6zTG2vqazDJnpAkqaf16tH/t909LIJZug5i8itD6ceLl92m11Dkysev6KdlJ5S6XTv52
vGZgxEC5LyOX/MXqCy81LKo0ePFnYG4x7HIXLuQ24+uDANzHEcsF5h/WpIBP3UJjQpuoJFQKBTeO
rd9s/bE+faYiUubgsSpPrYvuaen0Lw4HrEKVQjboI55830VMVfGrIExlvYtwwBNz4vQg+Pmsz4/0
F4ZtXEWs1Ugo5JeWG9zzm7kPpgwbWyAsrdZiIdOkZiYM20DjBTI+TfhPwR9vnfmGSLDXZVYnQFQ4
UIJlnAjO5NuPjFsrx4Dg/o8EpjvVI6rguKa6leoL5y7IoVVIjeedVtX89nLusEXdLHOmkkT/J6Nb
7+xRkndB2DoC5YZxNaRKsNEkGkbwA7ztxIQihTZn4gq0yC23lLr9ik86ti7iFvHDMHgBCgwzpWuu
zKR/a+eUuTrKuw9jKApDjTbpeVPOGgj7t4SfhqF2Pkifv21DN3AWhU4X1ZAJAGCHxU65cJxu5oNt
gRj0OPSVL0++8gwVo7VJYLobB6wTZ/4c+OTa64sRQKEU9hqHXU2NaRf/e1u7p4iOLBwz6/SksgAH
ERSiYNdQSKl00i5rcCVDesCB0bKBUtJwLgLnFhZJRMXtB3VMZJ7m0R/iSMWNjvFNGWsT4Z0DaTjI
SgnhSR6Meszop+OP+yWP63xSwZzvZFty7mD/bT6eMc+xfstxC6uaJTESRVeI8hhVStCWczkuj+Aw
gLeRbCNpZGKsLCX1T8LNR6cNBXGSzp39qSy2XYR3DUPRjVC3x2G3Ip0PfQMPKOEdekukAflxCb4w
Djv+AbUne9XtsM2AjsizlJ5msWi8l/p1wdFG/NtHG/J3HdmSjWE2zTNq8mH87/YhFwYMcTSkmlcK
1LSrf0poCEa0lwSFisq8Lp9cSV6v/PxqdPiT/fvfqFEBATaZHvjxTIe51mgBgvyXojdCKPPNw50e
MVeqCGjszuVnV2TLZu8uI1vqpGzVa9Ap3OaQd9/RHLglJRKeR/i+YyfaR8PyryUyQ89ksYhl0NWN
WB606ZHtx9Qf6O0A/i2jGreErBUar1EAMBibfH2OIHlBs96U1yufCe6l4NXpcfFD92OCSZUBu8js
4ChXb7SSucNANF4tbUgHUpylnRYOPZmoq922w6a+cmRTBNZ1+j1AtcppS+eacc0x0qItZn34Ff2K
96hIkVRNwpsWiSZUppmj85J0KiUw9UicBPPrXmcDEN2xx5kDxVkhkrfbYUyoMq9aXV9TrIAui/pT
jntdZ8nsthkBp6grqvjNrrIvoBPcWudpZ34rATiHtoA70wpMfFUAkJZAatWMvbNEG3vu/XFe09B2
g9IUZ4A8S2fWV5qBwpZkArmXAi455gDJtj/Bb7zLMYBH8kXUF8tzALqfA+t3Hd7bM7z/YbmOb1/o
Es59IgzdjYzwjgJOeOzijyrNZPu0b9BltE60MqmL+zDBZ1gTdiTMXknoec/ZEj5Ak33CqXfe72ax
tg9jmoX1PINZzZjMJfn2Mg1Qk89q3TXe/PPntlidN1mC4TFmaLVEQpaU6NtZMI+epSa7QARL+5GW
Jt4V1a/mhhoS1kQzRFoQ7TDwl02i0JO95+6oZyGa1V8igUGqsgx2Pnet/nr8M7A5tYh436VEiqQi
O6HBVOTXSmfiMIF/r1dsbI6eVs5UwD8mXqYAPr5Orf7ZOSybAjGQJ5h6/OaDzp9F3gz79Mh/BzV+
bbh/WJmYWQezuQN/scTF4LlXdjKe97HIkgwOglCpzKzdgyvfn34B3FCLWUfOV8XRR/rvYND3wKgL
pBtNZVoHaCzxzQeH2ZEtigI2TR2dTyFEdV9NiSd4qvKhsT6YTBtCdTqRnputocna6sTGHZ7X+DcD
9jKnX6wk24GNRtqmqprDR6aC7+t8wY81Y3H59FFYEqQwoTaZvhMjYjxg7GkoEybxHQFbbXwXiUDW
9z9rhZP7zMSXNYbO4dkKgnw48EuCPA2A7EQi1MC3X0r3vZJnySCuwHOJKoFIz8va7soOBZub7qHg
vlAkqm8Kks/Zw65vSQHtITpCzoKyzBNsFy6GeM+kHJLuT8tQ0Q1PX/sjLkOS183VCxhtOIgPscDg
6MGFW33KeH0wxKm28N7L2J9qmqJ8VWWNKprRmz6fjlfdWOvmPMbmX0/6uqCLSzykdsE1Teii834D
8qieP5rNaN4dU1VASbLf3KJVnQNdEBVeekAa+o20xAkn2w7+4ReDO2ELGZoqOGbmBlLYyARCzvDd
o1PjVHogiXsnh6+uAVM9Hr7oC3YV4ygcCjahoCuZ2VSC4XAOLRwh8JOcA/FGwbOpXDk0AsjnCF7A
lXBqSdMdQXY+r5AcqIx045rIlGVHOtjd6fD1H2TailXs3s6x7j6ahY9eqZjJs0UZkqI/6k053Ekp
ubKkCAnfyAYW3zjNuqUQk51E3cd3fSE/jg5npV2JL8n4OzFabXU0Wc7BWgl4lM/F48dAX+NhIKhi
cPBIjbrW6Dy9eYDuNIcR8iqtCjEuEeVjMKCeagQ6vqLcoIhWrKjJGX7VnSWZJU9Gxn9ShpVVaaX3
HGzDpk5t6FsOlnTLFKcyRq2YV/4v0knXZFtIynHl0Mu83ZmmFPiizscon7jep/0BI30dG2ZMe5ub
6fncN6AO/8D7N3n7gOipG53BTjjhXKdbPt609gTJc+60BlY2XhAdaDtmaEd74+FWZmT1SI2qogez
rqFo4q4g0pDDFibIHDdFQWUU/Tq0v32ds+HHSpWtnhQeOL5fZOr0y/lM7pLXAD5udR4C2nyWHCOh
FSgCjBiTv7sWQY+EwL2DZw0CiRN96F6gA0loZBHQ1NRK+wdKnuLV1gqHOClQwUQs6xNwUhDUeElq
q5UGLZk01L/ra2Gq4qEY8s3hRJJSwCEjygsti5mgtt3J8qbZGP37jRvFH/v5SWsokI3/wfZ6/Vy5
aW7GPwywqgagqShnQCBhWC37yBhJZZNyMJ3SYbjhsopVmm6U6S1J0MTxiCnLTxJyurNMDSjXCL6G
9cMR6sQ5kzT83CHKxb0bdP7kzmzhVEbYUjcObPs+5Gq1p/dDJFCAGqi/T5uNR2C6iHXUSwvlXnNm
6tOatrWvr4ruNjCfDn61wa6GOPQS+8tnaG5rzwz9FAzzDOCk1q0w9KgoD8ev/Q/G51k/I+aJUhmc
d/mFnyj+lwYjq3ED73yWDdIyw4zdhVF7T9+0erzNMo8Vd97RfuJZ6G9/jj7QZRynw/+EtZ4qUxGT
nav9Srwm7iWSTR2vzdncv6Zn60faWkjy9syNsibbP3S9idDVAYrDK0O3JFokyQ0XsQXjr83ff+tW
WJfbcqnjy7sJbSFCcHdeWHEeqpCxUrVgVPS7AhH6aHJSjsvIqOeiKYBq0m2RF4X1WYMPvLXwa5E0
o2rolT9BQdiG1vF4d5TPbqATFkTPKe/fOvrjYpgGokh6uoRzG9fiM6zT7NVLhoMO0EeAEoZH9Jqg
1GVgS7SXSd6X5Avu7WgsTwBfxYyI1YTXiGPLYpJxePoryLgYSl2eP4a64e6YTL78sYnUbWvF8VUS
zf/DqOBojNDa2NX1MqIrVjgOiSAVcbcPk69Q9c/wX53UHOIV2SrPXIyNU9op/UqW15g+CSoYvW9I
EJYyWZ/IQ5q6o7BTdUlCRaPlQtRj8YHh91k3z+pVptQiEKW16NfUvEgO9sMoDISjnfhY/b46Z/wB
WgafCq93hVaeoO9iCkFotrs0SfWlypTYIeWjOPKVirRrj7hpkirJOJSqhIBsh+GMyD+yGzCQdy0u
n6lx3xnTbEYEpWltUI6gTT2a5alJapv9yN/ILkDyXWDShvCuiFPPAFxcxW65XHDYnvO8ol2S6GUW
pQFJmBHE3X7Itw/XzcMm6MCQedhiaMSQg0BYX+RR9tmmr3RcgVu7//2x+gRXtAUc6YBDUMiUA4FV
I7337iN9nw1IKThFSyWgPG70Wnj6HTheiu6/PJms/+eGsJayd1f57RQ8WWHb59n+ZM9nyG/H10Vj
HQvXSl4Zzdx/70NoSHfw3PdI7OUH3F5RjGVOBZB+ZMnaJOgb9zvdvg4A9LBTJ+b03B3Jw8iKT0ua
fXsXJFE4537fHDBGvbwsfvn72R7djeGS0lAS8l7Tt6QmtTqVeIZ5SBqis3iZy/ST+eyHoi5e0qlO
BEJJGpXBiUqBHBS4wzFmHSQD0AjwWe4OYRuS6JatM/8NgkqQn1+FMt7rMyNFDWB+jW13bGqiVl1P
ZaqhBDXCFzaHyVzioSzUfXRZiUtQ1JIBAJuu4g2VMjzcLqIvBiHd6UIK1BTt5FzQzWc3TzLAHyGk
dpqyIaduc+Wc1oAmlM2C2QoNZO444l3cQp4vYFGY+OqTCtxSrL/cnDEKGXM3YGCldlIp5At+O7ES
PUxSOI087VKlSqD75ckvvvaiQ8dvnFv51/MB0QeILX5XFdoV3gjycfMEKQ4lArVQ6s08WX4XDyh0
zBVoyGmQaJQWGDWUlx8DAK8oip0uVudXEj+CWAYSV6Hewe1NCYOBfPlEsuVr5lisF4aV+HHf9+fx
iIK92qyrXykY1GdmTVu0MlET0LXExcngUKFB9h6xB3Vreoq/LYribGIB5PXJg4dgvLmANiMW7r4V
wmGgf7mRTM0dHmB1qV3KZUmp/vISz3wbiN3cjV/imqVFUsfhAgvJpF0N4UsVEgz7xF1tWG5LBZaf
7U2xXLhP60D8jDzY8SglxLgnRM6Q+9awp3ub0Fdp6njVJnfRbdJKZClZqfsuRWMuMjvF42OmQ9nU
91W6o2wjX90L9KSzt2NBD/FO8LpCZZ+4IKqplpR8Mt7wow822pFW9zdpcT+yZcvKIrZeakz8Z8jd
wGJEFz4cnOKs9TBX8jFy64luJ8k9d28lQMLPmcODMEgJYjh+7+66VF7vdK7cmULN3CKd1eEMW6DF
vKaopCpB/sbtWAaWb9CGLj1wH9DZd8kHnfxhs/xTI+P2xtL8MqMWzLpeM7d/d2dnV0xlKOmoVv1v
/95wbv7ZyljGITy3os3TKjqY3OgPkNItkMOP8BX66ECAbL0dhtw2RZcb2O+c+axSwALmwJXR45eJ
d1Du/a6gfoatlUu4tBNAcyHMbtrpOpiDVWv962D2RIK2BOMxpTgif4tBasUITOu0lCdr3Rz2Exla
UCSaeKjkOtJQj33ObYBDAgmQHtkWtFQ3VX6hgnv6qGdZC3tJ50Y9I+yZ6rYTo2k6S2gaisuKe2Ge
X2TNgQp1/4ed59IRYbJH3sRRD7mxCcgbdNplzPU+ErUV0Us3GrzYY7Df8Gn8K4mHSYXX3Lhjk5us
2rndPXjCZ9A0Zi//hMwG0AD1h+vkh2edsRNMdkcym4bt7zQ7T0kxwO7ubdBAz86q1t8QvrBnGI5T
fvQkF1CM6PDPuRwQv4DYhKuhljrZ/Vet0GCAT5oTEw6oS3uVYu/lsm6hsxrKtesjc2ohZRHJae43
PG72rz/aSFGJhDm/FNVJYHWSfslvRVCVFOeKJ78t2pL6v8nYV0amPSl/GsJOIL6euXspClR+ZqUt
965i1/lqTOrAB/3PiI5sIquTJxPI+/WuUeqOf5WM7peX+tOOqj2wndoAo25MbGPKemEEaoUQ3PZW
GdKzIoEzsofbHFbHykWQ4SFW9Bd32Bb/UG/o+TqzopgtyFkeUtsvOugMpnBx7tQf878kwpZe8dwo
/dIIuuYcusPC7TlbdiJBTkk9tYAcYSpQHOdryRWTdn+M+ZNK3ySDgskTrV9pif2XjQlmAXvqytOL
WWDL3KUo44RDpCDtd+y5IcwXVsHZFVVmX3NZClH6NPXLwzC4znVPc74cN9vb3UIKQ9TKwET1xlIn
cpnb4FC5PXjWq5i6MJNgyp9D0TFlhjtLRbAfF4zDj4XSSM9JyeqtmgyGIyJmMNtLq0bMIWIPUBWk
E7P9EgwQg1lGDCq9+sJIEqK/Y4iOFIMoGxj2/KiHX8wNxS1Siu6sh2/kIcoDCrhYaPBPpQNjHb3A
VHkhMxHGKUX4VVaL6hoD+0QV0Zo9DUnPSYtj/ZKXfWpB8nuWmw8/c+gvUTqR6ZYqGeae1MO7bupS
HY4ZR1I9k9oUiqJTd+e8c9UKj1+pm6PsBttjvfAeSKRhaqls3ybN2UiY5mLAlXQpu1CBxgmLRzll
6hS+4KYkJNtuk+3HWN7U7R6xYwFp6EAh9ASObxSq06X/Q0YDWbzMgOE1o3TxJ/prBgRriwkR7qZa
T41PeTyisB7fcO5uBsdH6g9cXIRhrZVLub1R40LY1Rou1UhZDw99es4c9vrO0xVr9HXENZET+LdT
BwWV49ttFrPUnntQZSCxPfgiy1uKiAmla5dFAUmlkvisM/fDRsxchchDA84WoSIaqpb41BQgVRmu
WrKZhyZfawQdUqVD2n0saQroP0/suHFLZpVoRjtaQHfLSLeOfMUC2YD2WH7UXNf+/kYhY0S16SI6
dL8Yvg0O5khFHDn6FIQAr7vHuOlesWks03yUh1zFHKZ062IkC6CkhlJleuDhqDCT9y4zOaU3pVf+
sDVqo0zoRfHlUJNMc25czY3moBObsMDhUUam9UrC6efqYJdR7D6HXFf//3ky64Qg4DpMBxq/xAFt
MkZE4liX+Euedp4einl6XWLmjjUPd3wbpRVHY0NuvNcHOntZlTydZrGdZF+mbhsnCFg6+DUe9O5x
Db9MME3ekkGAssxZP1lSNejWyslVMLMNO8ARf2FyTUe6Rqcd6Tyw1V8fk4Tq0VavP+dgh/5GEzew
/aIOxul9F5URS++39V5jP1+9IQpBh/gbg57Nye5t2BOZPFY3gmge+34EOiVWxDMgosdMYyY/0miG
0O3wVdEfId6kBd8nkbrLd7MnhViQThgpJH8CLVEWqF1XDU3iIhidjwl7og1ovCvdgASZPJCUuG7u
eWvYgVrg6S2hFO94JKJ03tdSN73Ld8QJlhHG3jAZVmF+zPc74Zro7i77nLJ3oMnnW5XYB4RC0rTh
fjOaDNhTPsVi1WvBUQFhAGxyILdS/cavoTups8Xqno0+h6mvdZmkeV6R2mF4QM39HQl6i5mq1tdH
ajIZHagWOMvwSXYAQ+k4RSn1UE/cWZL4v0ts7pFqB/6M51bKJklvVJIUjhJcCJzmoK3f1pbSimpw
upbng4m8bxbs4MmJ0M/est95vA90MyhVxkN97eoBDxGpuJPP84bdeQc1nkRFin9X66DLYqYC/PoX
y3HFVQWZkBZ0ZGkKBdfkFt/zNWdDg4Ir252ilxpyAtVHBim2P+UjZOOEIgr9wepPGTn0fIxOxAaY
rpAvNLkTzOQWKhBCj6aUClYw92EexfqgqZ2FszF2RtBfGM7VC0O2Zz4AxqxlGOzEqwV0XgQCUhqB
8I6q6y+87SkkqGSxQ5Et59ueoCkh3Tmjn3/LF4RADrheGWtLoxW2ymEK/wcGWKmldCOB3etO8X0a
efI6MG6GKyuOtScJizuvQGDjDqYVNtZ2RwAdolbpWSIYUZtnpgva/Bn/gpyGwN+1UsSWtlpEizaR
+sNI9XqIZ9m4YF8hgqDMXEpobPMzzx2rMYyYD1YIYZ5tMlTV5+AV0jgY7C7Z+RBktGGhv9ysufQl
sSWEdVB46knD1rMfDmeMaUaVcD6WUI61QfEyyTwxahZKzAjp110D98TTlQKhuleYmODne/k3dJTo
6l9dpHYUDk3FAOIacB7CX2AO0QlEnuj0TWpJ6mon5xcWsTCMlDMVwDjptUP3rMDdVmCEU7NualKT
aLOvmWlG1YlMn5znmdIuIuTrVZorZsEkLq0YnDuopvw6Gz9azsEu5/sYWhFbkVJHjiKrhAVXJUwn
E4eI+LzhKHJj76DwA9ShhKWxTQznEP8Fo/2kymTn7J8D2Q03BqGSqka1R9Df3OzXYIitHJLlykrI
twLDT5lwcadou0XQVGpChisYixnwMvvNpC3zEIOanwe3+hEJCGu7pnIqPMxW6SndagrLU9Lg4fQm
tv+rR7GXJIBeVo6M8a8HxzzhfUerfizBf57iAGS2290idLwMeRdyrj9Sfsa8AF6d/yzZlimkJuwB
2x5/onOLjquwAkZo9ZMIoT4sVcNp/SVfPcXvZbjukAXJqnsMSrMvE81u8ZK71XTkuX2WTdX2+MLn
WTY9qufK493xaeIZsLPIcxp2yRGPznLe2T3lqIr8HR2k3si8roCU72ODxTcwGgw3bh14teuhzaq+
2JH4Soh+0/TLFdEhr2o+TvcEfHH2LGvhXJyNYL1nzPYVdKcHACd443xDmCpTg1+Zg42MfWVHnGIn
mcknq/ub8PwvPr/mp3UfTiYfxnfv2Ah+xRfoxH9hvDzxH4U7hW5O91WFpkPN5m0oUGjRzwYMg1Jo
T7IHU3DQwGIrjDrPpkVftXfbvDluYIxfuvEXqPf6YfWWWKi6tuaglNa9QZbIz80COLn82xNqXWd2
8yBNr8DuOOuRwwhGrvUmRdVxpt8i2IK1ixED4wV04dSrZuARX9+XnTviA7H61nXetRKtYKY91KMt
I/LUq1IrqlQrm9rlttQejHSNA87iDCzG1sJy1Lj5PfK7hz65lLCDwYiDG814hPm+kIKYa2VrbtRx
+AvjwtlWvCG+OLep26HexpQwJKNnmovms9MWKZCCcOSxjJ+8pWShd6Ar/TBrbAcQB9OYss9G9Mhn
qN2hs1yk7syzs7Ccwp6cJYZgNU1N3Uzd6ZRT802kpDA2be8EAqilPPFn4k45zelJ37JWjoJnzBXz
eEyqLJHeBt9XwX20FJHp7IScavTcbbXnNGVPcay8W4v5oxNgiwmnc07wCcZUL5BSvlgoVhLpy1sT
QNISxPnVvJz+31yGaRVGODZm9T7Jqc51qr4X0q9QRoLnuOBBTVN28U/xrBcQ/lzwTMHQ66JynJg/
cQG9ileeVcCfFIcOd2vs8a5hP3UcoEWanTJ2BOnVLSQDC2m79jtbZmv65FoldHVkNVv1Kz0q6IIN
n9hkBdpz1NWj21pBMEP/ishDg84OZsRSDixc5kSPZVk+YAs6LfEUgytTykxu3PuY9mXK4hgWltsJ
9lq6nmYLCfzGNG+1rqrAr0OYpXSpcf26WpuXuzg7mJEFF2SJA7/zb1gypOn4FKe5cB1YZDSsgiw3
qMkUl5VZkkCt3J0flM/UIatluMqYxCqego0O9bDBC/MkMcZGZntQo3lUZyATxtYrFyhYWypizy/Y
G1JeO2/J1HoYlrktGAH4+WAGf6o47riqKUBIMDbhZn4w7AgEuj1zXAYdJhgCR7/xZ+hCveKwXmtd
CVkRRjB6mRmrPqmXBdPKB0KSRLCm+/zHcJcN08Pxts4kvxzfoNe9QHKIOZFjBx+wApdz5uZSVLOg
a5HOw7Oulki67cTeWNppyX1iu6iLder/v6X143A+A2RoqHMRYb6XE1VtWpXptDVATPUwiBiC81P4
8t+PGc+2vQx8tCtrpZlzqO6nRbSDl/NxP9JJMF3vloI5JDqnlivr8zMhGiv1fwz4Y3afgjlf92a6
M2QJqtGiilvoquFEBUF+PS8Msa8r55RZzkvsi1wLzPZGTWB3JhjAhKCAWWTWH/EQJFEogRd75iy4
ols8iG6VecjXEUSn/pSgTnb/UHuNuZRw0yh6HrBHW61X0/fi/4Sd3zF2YM1LaDQKMFlj51+rwEqQ
1NWq4CYGgrnwbRlgzgfXxcx93j9lTO9knrzln0chAEsZJ+uBI3Cr3a5MizEnvHNSG3oSIL0re0+l
imFiMRR5wdozG2HMSSLYnZhmv/dyp7iC9F/eu3rLalceci9hm3E6/h012TZRxS/rSDzvq121nubO
OhCbkbtoo7IrB34Gb45a6q1aJU6pAotXqIyAUwJBna12s9YvHkeRh1UzYaDfzsDqQRx86E9MhzaW
SY3SbBAllhHrs5geTskP7X6m5LolNEtkqCvzbcpUCHBRTQUQoYNCnUmDybr2EDfQPSXVoYegJEY5
F3zf+o1owrg4A4yj+BxN4G8jfvt+sGBc80mnDbxYCw3KKchmjwBVsJL4QSdHWLoSL4ICdL9fM7Oa
6fqS0H3mUhqMGVi9fBc19fffGK3Y+dO4sWpDih9qg/pYklkY3kr9cKJdtgsS0hnjs+x9UXlraq0f
GBaeF9dQUR1NpdlZMP7yK/Fzd7Oe0AVDNVRzLz10qnHPLzmIobm7xTQm8DLUR9oEwT1iJKZllIt4
RpQdkBkq9DlEnhyf+ikYCk63TBXu5t9rhUi/niEAJwXRAknHPuTIsegAZy6tZ1jv/yDxq86VbWQY
spn0s8PEvmBVdjEEsfomM1RVzFFdiS+M6lmbvwVgIZoInxif+M05+n4PehOtt41++cc9WlgrX5+A
yx2rkMRooDd4YSK1nXp56WqnnriZnrr2oG9l0vgp8vi9Q4gMziv2NNFNH+SyiF0qWKnkUqEl/Tci
rYxjk49SNpCf9AJTKvWnHVdX5z3avseJXMB3mGo0ADz+kJDjQFjelhbSJJ120i/ZY5lot7zdZBa6
QfyAd0ewEQW5Bvv81d7vINtC+N/ayEwKxdXqTngUObCiamf7t57EuRjaxgOBk2/Kr/sBv1QSBwBX
UM9VJ5v4iRlpQCr1QB7avWaRr8w0/UQpTVlWAuhQfTkLl0zTLOYrxR0J3u+WxYBWXCXJ02NHVvtj
CtpfiLphBT6eWtvcZEGNujAsNPqjZg5V5uX0cWYcsh681152f9DV4lTV4L6DdvXS8dhlr00NVysk
FMLkmI74gSrxcSrAg+dSoYZZAK0n++V9b9mpqqqN1Lim2sSFxSET49CpuMvR41rlkbG62UJ88sr3
KIn4+6zYMWqwFbPBm23OHm4CypL4FU52/yturhNEK0QRquq55CgvTnru+GFDhh+ilHER0Y5BuK/U
p0hibaIaF0e4gEpmPgtrHy5tF5elB6yGXUkQXmvrk0ZM8mKt9+3mtgKEarj3R7a3G64od3gMKGCR
+BgySC2YolMfP1ZMHH2quKEs0jtEFHCGkIbR3bsF4SejdJK6LRl4+b7q/R+E2Pd8p+GZr4Usl8xb
iQ6KeeOKrb9ldIbzTM4kvWdUPRqs21mixuaTu76UpqNvyYegbaEdE8zNTnT0SeJraz6JI3RkYRnd
xLvXzEAXGvHfdJawtGEY2nQ8OwKBe01COJA1i/90+l/+DaSy0U3S66GA7loFm4t0gcp85lnXov8o
0TO+KHuwpP625ez5+C6BDKPCkvmjq62EPbE0G9mwesY8qbT8hyYOw4tRy+cE1DPDjtV0dlWdi8Hj
9Ka+ndDvgXvA8PM0lCSgGB4VcvtcJG3WSWoVr/oHn+f9kr4NBe8k/fXuMMitb6pDsS+/BUYkm4jx
jkvoShV2WmSOyIcB+BxQ5WftPxje12QWe4cPzEr9g5vUpj3V4DuIbcHRXFfeGdueidVxt306j1Vj
rohUf+zk02+2VGUFAqPZzsiCJ4m7HU3Vrof3aYoQK2vjlOljImhqrj8w98lOHCdHFOupkLjczAXU
N0Lw6GVD2X9m+CJyVDH/pTL6QWkqrCpTIavQ5Iy0yr3jFIFdOk1MZk3OkxmtVfWPKAR4WsB63dPN
2Cvdu5TK/U0lnpLKtZ4KCcDELu1kArREqXtKv3iQlEWeOJv0+0v36zUVOnzMyYIMyvz1auJo9jkH
KXGZkJ72Tmsnt5AeHMAE1kM8eTHGIDaG4Kw4RjHzvupG8qz/D0B3yKJV408mfA5ngWWJMZjnNtB+
MZ1phPVHNjhNz+6Ab8ZpzS/YMLz6vwTU42SrFg/lTeavy7dxkNO0/lW06olEU/0XJlsUVXeOQCS4
sIGZgI1rreTy1e19LmrlFKuxEIREI/QPYfsV2wtQ44+onpl4zrHTl2LHXlRoeoyxbxpv9GNC+kTJ
au7TO2Ry/LSvPGPZHJVf8O+lx+6oMQs+LpAws98DNKj7ogtpvUl0sRFwfxgE0tcKhMDELDUtEeFs
TP+nOu97nd2rL7zVUZ6+W/7+hJKwP98OcJVDaLY9Ftrei0qJAg5rRyiNIhAmsazvbll8la0f3yxY
qcu40IIXe5KG1L4wQRams9AOwijHPsc/CW+2+QrK6n26vqlKk/5dO0UO0dEsBmwq/bTIoIGoXsru
TVEX3R3h+IP5M+5hamPShFnXQ15xbvKf9Sx8bjqUWmnGSe1+isPuQJAhQmMLq7RDzRFnL1ww0+/H
S/d9qSlCBzreZy67RCKJpqJ4BTj/1JzxMQsHQSntaDaSjHAIRTHZ3TueprU3WjXu+tIcRYDAbKp4
kncX1kVvzkN8MfGalzhr/6ROFdBdWKWDRflXuTSQ30AsqY/r2A0C67/YR32xX7p/pn43BHlnR1ZJ
0A/DtE3diIiErqTxvAp+A+Im3ocMk7mZ4wqZoCugE0YHexOzFpGIjSvWXR9Ye4A8oN70zSnhR/LO
TwPKEVUr3PgTGoXfqRO/TvwmZk3vMlJHImR6HNdJy9zRQdmqA+jFl0+coE0vuD0BqW1PdvZ3WnDN
58jCoaFlb1V20ZQV6PG2yvnJCc/Ji94zzdkRftpnMxHN+NmoeQGok2gIdX37HGHiGqbk5EQq9cgA
sczRIxaDIEQUK8VtT8R9oj6bAnUWku0IvppEY7zsKnDAntkBSHb8dVeJPwWkHAdyO17v6yr5XdCy
qgEJwLmlxZWRNBPViWysf79o7PCvN8QVUFlhVNJ03vUZgTcJHXGfkVjeMGuJ0ioUc+wDUopr14NE
MniQJh2Yh6DsP7eD1KFp7d9c8RqkiE6r/ugdfL0n9K3Dklap8g7B5yzLBkcXDIkxrDU3spHeSLDq
HOpc2Hyb6d9edx3qntpe9BFGzsh12chh42QfyVM6rkU+sIYtDbe0cxJ+BZLY9we/Y0R98N3YiSiN
CdrJ/EyP5ONSFmj0J+Y9sEUhI0nZpodrisG18ndMvjWWWsBqXbu7lCx5fftq98JNJ2oI/vgFF2Ru
X68rP4pODNdAg+53Xw3oZpfVt4w19nLwvUskKIbZAK0W26rxAvSrCB96VXcfBefy1dm6nkeYHF/T
WvyXcPmgNUoW7escQoltv1dTpK0rV45t3SKzYNK+ID0GoJ7fTNXOHaEH+WJ6tlukdUW+5Q0TMcLr
lGRGNDi5ZMi4SD70XQW2n/W2e5FHJVv5eDQidaLCZYz+WS8SZeBnqzsxqnY0UIB8j3uJdBKDab+0
kIEQK83CRBA7e6fcowX+pl7VlVYQk9pYniC8vDAPk5F/5FUwkkJ+9OsbHZRjCEv5l4Aen/MKG9gH
SEe9PC81Egz2nfeIKmchnEgBdf0nM06sItO4prqkIpsWUONF8qFF4X3hKaC8GVgkZFI0KvNneDcU
Jx3TY2P+hP9CAQ5nGQiUtp4VfmvLnSinfRnzV6rbUdgHV8jHiCRH8iCWapRd59GzZUUS+F+A+VBH
VmzQ7tRd9sU/9ptuUS/9eoU9ABmfCPeEAL34FswDeGycsTAEM4BwVo8U31/9d9+fIzxPcykuzNne
Tthb3dTpYjGsKLJn5H4y3b4971gjD6SGiJ3VQlqbJoRF5pjF9BCWQUpj5mlFOR/Y89rRWOlIwkQi
NhddEq73hy2p/zvXcHAZ9GRUxKdkBy39jMvGSVn/srr9I52kkYzZlMKHBUy5/2PNwnavhN/63uTG
wtnVC8J9FMytGaEqJE/fa/aY8U9ymAFA8bhqxZuZI2cOyPTqEwuHdB554qI7Vl/WiAhZkVEDFtOu
1b8h7u9SdT/hXk6i/U6IPyS8ZRl7Uedw0rTeUpSxL7Az5WNrLn212ns0FxxUGraNlAXHdELLddci
bxmyyJHcgqLLefN4oyJABDQztju8zhDR0aJmY37l+vKOfhX6g+UQJxI1Y5Geb0mMMJTtMIukma63
R8Pxko9GZd30HxDOGAGUzn3pVA+AqT8GAuW3D3cbPjfLRl0K2sGsA6PkaM2XnQ+tmIfmMU1tjLAO
UrVupFwIZ+clYX06NuUIA9oDXCd5F9XuZwYhwrJ5l9nOrJ6J/LjDt6qhnseQP+BDNemW/dSnZ0gQ
0Q8vcaVXak1xR9w2oZjGntWs0xCs19AVAG9xflwRGuMBP1RxTxWgHMv6kXf2/mHAOo+F32ABKyb7
d9MgqrIkGu2wlDDvRMGHtwNzJsReN+Bz2lqugW3uKRiqdD5LmoklWCmkRHKBmqjcNHVXg4X8r3BO
bKerUFhATHvXVvT9WbSHAXnjptaB7JMfeUahCXWkgvSHmCXwksZaSA6gJ2rwwPthhCz3NQ9kuiZx
a3e6BQwxbrNlNAWlVrAEGowz6W1hjGCUn+FLOiue34e5I9eOIufSzvYsJMcYr4B+B/70AaT7fTiF
rRfeAirkZg6h9a1ZdZNx7osPlQdezejM0u+Yhg317brVSLgdfS14kPNW6ieIinbV6xQ0q0Fbz4yV
afZ22sKfbVyMipbKQ+Jotc9zxcU+KPAtoU8R6S1fnnsacLQulLVy6ZRHcjE+rq6a5/uc54qEMAdb
HS1Qf8lHLUCNm+RjJ3wusj2fy2Zqdpc1U3JoVx/sOAPJB4+H8QXE2T/n1ESNQcfB6S1Kn+iB9RdL
tZ3sGlHVzw7ZHdW9UPDGgEQ30cB62SwY5BIeiIW+P9ocKUziB/P1AJiRUUMFZNFb6npjhkaX5KsT
XjxlUFaDZI3Af4jC0APcj1aXkGkOzrlwl6EtLQcORjGQp7PWaSl7r/INTMluBVMckyp1YmaT0kEd
HG4IG7HzoJV3gtLljC/VogwvmV9wlnxBNSY1AIDj47ajvSvoB+Ppj4ADgRTxBeFGLeBcwl8IQBQ6
IekJOsNOiNYsnOZIttfclRXUEWGUC/1xlUMhmMrA492c33SS5fmbNchUoLX9C/gX4PJEc7nRXz1w
+O8uQ6AzBXYQ+XeYsViFC3y3PLsq7ZuWCVYR3p68n8IdOIv0gg2qgj5Wm2jlog98PJs/K82tuXSj
CYeRR4ZPdRJTS9qYcZbiYJteoNqxoqoauYHjaVUGHjExMOjLNDk7wZPhKQ1YR8Yr+VIzwAVaIdWn
oN41c0Kxg/Stp4UKBt8RaKWDFI53BomLrNe6fVmze0z/u3i6W6kjhHisRjCXnQavy06q0znIo7L9
gY8QEJVT6cK3mlRbxbZGwdXq1ItLANDF0yaiBSsUIGeHPez14TX3siEDF5HJY6BojhQ0fW/87aHX
kBigDXFzAq9eZb+e3ugdxHoDzq/OoSht0g8UEXq8iLzRFaX2bO78gH9FGvva5hFoL+JahygnnlMv
IsEzXnwX/crTTtXWse8U9/w9pP7sJ7ObYiv2yh2PaFBWTFz9VGIo5ZMbmlhS2xtpOC7W9A38BbLY
AdWQr1xDKPC4NCX5rP1ZJmNqi3EVNDXTCtKrLy/7FHuQUoSLfT4Qtmd4iWOagl5H2slqRkap6NlI
dRzI2ydpKQwMR4LsjQbjhZU6Deh/CBbQ6d1LWbTsRjCBlHeRU7amW94pXj6x8pqGwYmdxg95ka4A
KFTwcfdBKttdLsIhpeXfIBg5e0CeoxRMxBYzGkiW3PG7LVnhFjVU6wmZsxxKjK5647efWBE7MkUi
b7wSOoeIQh/tN1qI2aM3tT1ok1ApCWXTUulyk6+q70yrmx/5XBQzn7KxkUFJJ2xetYe1D2L/FF7t
n9z2stOUVtcbM4fysemqW3Q/r78oK4d1SJCqQSDytXp0gKwL0qg7o6J1hJAyY3sGEHHTzL9hFeQl
d0NJai++1SKCx7LO9SQzcQsZSyk72O6Di6W0fN1Ra+bNxvkmt/kBGygXj0bKgO/Q95jD9TIkkqOX
3n5Ksd+n+Ib/KDl1tsEjbrJLpUigHfiZxCI+xBy4JfK8BzElrh2M8OxKI0t5Jy4CdP3IJU5Zgq39
ulKhGJmIFfuhsve5z5pzm3ByCjhdhO9YsVDwoKA7Z8ImG7ooMXsZsCrmCsNIye8RB7Cx1QUpf77+
8HKFjCh4pQ5WJQKy2JpN+NRAROYc0xGk7LQ2GlOjdiH642LS9y2xcJ5yCZCzPP++lmmU0bm01YGk
7pS+wCkiP8AJtcUujM1csjv+JgmRLPnMiIOt4KA26+7sjelf9nQF9fwqvN3Lz4bXztnU5YPyJ+pZ
l6EArsv1mDrBVNnOTWLKiRBN3OtI0BOcNSaYw7pcTVRuiKY5hA8cDvnUDGFW5yVjMC7DFrX92M84
f2XPcMEbzpDxqXkRn31qlK6dgv7U6J2QcWNqkh2QcqlBO3b6gJzv8/51k5HIWeC1gKIhF/NmAH2Y
1NlBaBwdW6zroJu9R9Vn5E7HuaBWpAL96vTPqpP0HGRCeZINQkmOKLEkQpco96P9GBbnevcJu0W0
wqTPAKhT8gE7J+Vtp3T1KxI5sG0BYO3hE8DuV3XHBA5BocbwpHDyGulguFUOMNJrrZT6MFL78cKX
ezWK14X7qkz4hbcCkvriT5RtGQkfd5eIKtRrNqV/3rtQnjMXVT5ptGurzUVdP7KG4TTL5PrKKDDi
gE371y3HhAl7izft1IzV7H6SLH9sXkZHVTHXcfJA1kL8pTVtwnJG46o/XLQCyK9XAO2ChJ4z0DSv
zUZAokDHHv6uX+7vdIYXn63f+gB07T5GEsQWk4k5Qn7vx0BL7i4HbudyRQPR8VRmJWg4/GFPR0ws
0sjXmoR54iGkWTUaznzR5kHGw8tdcfiDhGWqBww96dk619D3hUfV5JLty4wohf97Nke2UUFF4Fl5
1rq0XXokONLQDATMeoVZk9OXAiQTc9KtjDNLgK1ZjTagE7uGqpc0MVpWZlHn7tLdk955Nn332s6Q
uLhpFIlkhTcsBhad6rAYFGcDC5kdToOlw/NhKoSmKzGOjuSHuSOu6BRF8DlF9afHlFtStBlxpnRw
AJ7BZvcfh4y0fmxBKLNV5n+7Rpz2Fw2qjCfToVYwXo6UT+Am9lAiXcbb+Vc6AYZ84lwyYMiV3zFx
fx/V7nHc8jyc06bNhcmJv9QF9JnF01X9bwNLqsVtD6lt3tslJJ1qcqwX0/B23YaAjYMA/14Mfkdh
upuxMTsD38TWSC0uGKV9Af7Hdhd6IOLeHx61oyoXd27f8Yr3A8sjlNxVDGM1QmfdeTxi06AzFPc4
rakcNpoAftg5bgwTY1TZjqxHE8n7+m7Fys5VuNYILYFgYm7MSZtZhdq2zThTi3tqXyCo6XvI8Qw7
xUWFRaeO7uY3AvcsJTLDLtelsTkp0UjCTfgCewFeOf8W5KvMj1ULYSpC5s04cFL9hJp86ypT65lB
WUm+ZQGYoDf537j2mdjpsF2V1IQaUIXuQIW8ej9dJqKvPMrE1ItLibzkrA4amauzYBs7RlvjpN9P
9U0Q1GSBB//qwgVN5FOtMZasNdkEexfTl9cz+xOqGkpJArYRfcbPHCHs6ONYBrIKCmRd07vCHtoK
VxF8g6Jew3K6lb6smkoNfE7GUGkocehappvij3rqjsJC6yyiC2FdPsm+HJB/uPBGRZ3mYq79WmQ/
GQUBmgmhzKXL1gw0MAepIA5k04w0fRi8QnL97jHG5H6uKX1+PUp09T5lRLMxmLDPcqNV3udV6VcU
1lir+1Q6S/vXecUTp+mOiX4CqOvNDO+YJeIgmmU5aiDSU99q+qkGckB7iMwBES9vgTCQvAgrPyxG
JxCdhc+rpaEGVeo79SmrKbwJuYt7M2VI8ajkyknRsslCzeiVua+c2beI2nAztMNNwyd+Q4gHvB2Y
l4C8uYSSPQ4SPgh/wXB3YdCaWd8aSBivXzGJ2nyaSwG8bPUIEBfLY+V42KWNR5YwVrYj+j1cGnji
lKjpplz3acvvvVtQDi7+IGXBx+1Bhkl66x+WX8fftLfFOXRdSZt+XsBPe/m3BEp1PnGwl3m/x4Ty
SrprZNqpMAMESaGMmEFC9ijuM3PlrwGQWdNP02VMTvidwsmaUG6cwa2ykqBLGCENfyS5/A9Pwt54
9eLH5otUrUrxJEe++HJejkY1B2EicbfI28GrNCVKdCwBk65L7/Y43pT2MkmX9LeuOX9CE8Bt0y4d
HxkmfPQLHNu0QMkLFb3Y1sw70JEJnIpK1kdJ21C9Vef3JVVxNFyYv4gl6tYonoLAFqr+ynSvoqWu
tOdiMHywwel0bCZMOfjyoTi0yWF8uAcXttA+pjGIVdOCwRiU7QMLwzXkmyHx6haas54EupLa8lqG
X3ZPzxi7jjCfQ/58b5/zh7aBlyrNIfW8jsDfu1WmY+fNsIiREo9O3px0F3ugwzX5BYKeXywMJtr8
kKDUtTznTeMszd6si71F9fgHqvaZNzjJAjpuVW6OXddYvTkKEDfJ+Y/CCnLEJ4iwFZOVk3EcLXdo
CdbpywhaxGIp7evC5Oq2VoXRV6/HPtrIpQQPLskDSum+g2mGUA9IIK5HWt/uudKqRgI/xgxiqmZ4
Rdr2vFBQ4VrVZ7IKH1HUYUKc7rHiWcJnrXSyZ3cVyNmZwvxxeoxehrYVpPBSdVLwJYR9gtvLC5xa
DN69Rg7uecaASzbkl9jcLvNrH1rujamEgOhpAVp6DHiv4rifjr+I8+1Y1cDEM6L0tEbt8cuByqbm
J2LoM8+YyLM1Ioam6sSc3svqsINpS1Q+RPrkSaTwSig/xzSATn0J3M/y+RKpoKv/jUt5P2Dv+Mbd
nVjYmFczka6xWJPW9QGmik1zCkxMF4kdRBWy31Zm1nleYmiMEABwzhYT5E5kF+Xx2Zg/lxa5LvDe
6tkqyn14xMZn1gRObYNGigHAw342rC6/JKJM7SYhdmZN2RNSFXT2rhbWFSKdl7D4PptWnRhunHsM
lKrYv1xLeT2IihakTCt1axQaZFZZTbc6zkrE9FHmPRBaD2IliQlTA52CAFcljd01nZH1/9P0vd8w
rOOIvCIIekMedkodNfcuC3ktUXVJVRdQ9iyJJkVjJCxuko7TRmJmdkHOqMJGBGmNckTwrNGN5CZk
t/+aUBvWBWAOUqdpkanSffbvmCehyvgNWhqqV8PnZVhwYDnSJd4hshdx7Ldc3YLyz4ycuzgjyrnq
aScWudzwYFk5VmB0Hsy2d+5d9kQZgT0cz7cErX0dVX3YIQN/SNrQvHs3soxD9414rnoP84V6/Ofd
ypP0IxzyF2IppF9tS3B62nMTwZ2IMKuIlhhCE1ugVRPBWEFp66qAgbgy9uktprQM5hnvdgnGBAHJ
tIamjxdQj6yl/M6mOe+iM6CfHMcYInmkva2UOWtEh+ceJU0fd6JKHQBOqgxQ6t8qTyXjMzIWMr8H
du7uKMKfFsUWhqTH8SreDv6M60X/dtoaL7sdhsVVJMDiOBaw1N7IrTb/B78/Jz6E213+7P74RUmp
qops/d4JEcqr8mqs9bCkUtRwJljqpoOeayvDXdis/4knLHO0LJzcf5YNR0XlMRRT+mTgPaqsJ5/E
48WhFQ5+34jjCorXlDgbHQNfwJltpr9B6EfesCw4zirBIb7F0Lc5imD6kWR6QvXOnSo2WbHujzsh
L5cchIiTx/ikzTd4DsIAMGcJG2Lg7zBgpfsIeS8bHYjmnM89TEIw+nMOzNTuHyYh4MC1Ubiur/2V
dVneR6t3Z7M4+EOIF9NmZu5xRdF1t+7WoDbM3A9D+buXU4KFDJ2kaBwfY+yBadqpEpYTuD5LUrHD
XlGvXBF85+vkcYQxTni3mYLaTfDCk6hqPEDgfEwT/CPynJBnnZ6ou+2ZyvRTC9BHTetMPSc4B7Hi
E1WDQ1sfEJjgX1tfbQr6XsXK8GaOR5xPKtPW50ePZ5XMhPXC/+Y1h9mowuC11s6NqObqTeqNFiiI
l4hSrgyplVU9WHc7EqWCr1SZ1To/+VaN43SxWZZMYZhO6/+LcSV2zMGVsDMul1dQblbqMFdaSBs0
7zXRuVHGZjINxE/uB4b9Ief4te6Lt3rsHaXLhk5bK/0iYBoIzFeBFRCyIMXF+4Q93lAYHN5CnW8m
Ruhl9nhzpSYYak6EXGfNMVhdxFNTmwU4jdAPnlGGeIKh+4Svz0lnjPOSV4o1V1M6EMn28JZbrLo5
hdmqlcqx++9pP1HYHw7rRPkDpw3R+AdSn2Dcuv+FZ2dlHXA2YqHC2w3ny3QOG+a1ON4mt8A6vvnt
mzlW0b3fze7xg+Yo/OSWTnRmlECQA6Xg/3NZC97cV2UYP/nxvKyo1pqoMsFCOaKuU/WO5JPKUdtE
Mh/JsFKd4ZuflmuWbghdXq9pi5TpRsMtIpO+jiQZL6xX250BFzE34nTVM7GNd6SfPdU9wX0ec8wf
QHFB/tqOXi4IU7aTIwEyT+JYa5AvzljNAvZW3z0MwlsCm/yXXM9X9AmjB0I4ec/rhN/yV+5kqZUa
wWMlPpz9876/60TPNRH8RH45GPyqhaOzxpKCfIEcFxOHsgrpwxeTbQTZELsb5h5r4fpmahwR86qm
Fu72xpP3EkMECDLuuDIIZ3ZQfuZ/ITbAEQkhVhy04oxFKCm+wqev8MvG78uEsl9HCuWfCCTzaaXs
U81lfhhJYHwO0mc0wTFmolHNO46gzBzlg33zBoqM3hvEd1hQxlZDKKJ9G56Egblx6bKXxqnp9+cJ
Bm8Z7LpmzPyu8toE0YKyGUBRpL4b+XLNrHI62rwmalO5DJHO+I5dIW5dQPXbUWFdGINT128Ub/KK
09N1gBpgusQySZbyw2NonwMrG8saSEnh/BjN7RLAok4NIhOG3BVce0+5Hxo9Mj4pQWNd7khwmSBu
MZsH6nUqQvpkE12+b71cxlT5ZNgDu6ZLGUaYtF+pyg2Ny9cXESm7qz4JY0kvHszkyPdK7CX/CX3A
BXtAyLkHzt1NfT1vuHolHKpBpuDsPFAWzD3PnfzLdaTtWb+9kmLNYJXe4RwgfWdh2xYmLZlUrL+O
B/ijKMKYiUMG1QhhngVi6adapmLBES8QPMD2KWMeX9BCyJoCIDspc/kK+lv4qkGF2+PpqdC+8BRl
5aEzLhOgorEOAaA92WGU+cpC48DNgzx7hDoq2V6EjQlowCxQrWNzObPdY6sMUbLksJXMgdc0T7zx
IxXwoInqGPhifh9TxW2NX3BWaUH9IAp62D1VD95sQxZM6gIgeutDPrdsRkfDWnvT0berHy/I1IMb
JAP5zMVDUVAj3GL0rmEqFv5SBwUjBC9OeWzoOEI98suRCfVbYT99h1qsbQ5RyJfcKMgPBsTAB5qW
6s2v24Cp2v0tDiiG0/hEyOgkbo9WDhu1Ipvo6uCJsz6evsEoN3NnvdkFH1wmvqmLdQflLMrOykkX
6MBfFBph2YXWZ4A2Lfi1sYAdjRuJPMzTowm8Q3yrM1wnA/Chs2TLLkM6frvJGhvp29wAGyBL8eYv
0W6+Ukz0ITUEighrQD4vlLRUnook4B/VMDnIPLquHubTjIzxL2Kt0CKUVZFS8Sm/10yMXQV/Frkj
KTkMaSEZAm5lP94Lo7s2f5ED1MGFZuxGq7mkghbUqCdITv1J8cH/ubjLtRRpc2in1G6Wz0pbpEkt
GXvbVIPyd4r83d8gN4a5Mo/CRVzUAqK5WNBe9eXhs0F6rol5UpYa+8C3NUJ/Fdim5xti3m1dK0ZC
0wRgKIVNOYIOG+lUfYIhbA3lwPVPTc4Ouiqtme8MSybeFZBX5iwP9+aBWY31Rvl2WhpA/OMi61O0
Qk+uCr/Uq7+BMSPq7yBI0bA4t1h3ID6f7uOJ5bqKqTcqVLXUnfVtoenWxxO0y+2NiwrUL9UOIai0
kSDIFbJSWneKKRSeEzJVM892hdAW5b8vVTWv3RLrYA++UI3hhd41T24HYwDkRKT1PB46tzlG8opz
s08jn8yKwVuPLEwhtLOZkszrl9CIO6H/ylDV+i+YDWNAWYkq9PcPmRMhWZG1JojV/V7Xe3KOUHTw
Gs4zTecLnjN3v1H9E+/TSekyz1pplXAg1qpMi1eRX2DiTvTyPZ5LtBr/xM1FE0LVlZkIodeCzD3L
/KQsa773FdyH7Svmt9N2guBorakWZLIgrpps+X2PbVCOuVdg8Y0+OeClcuQECZBAgYWSNcdVMXjt
XZPV3cO8j6BLc7BYsFajpSIcL1L9noNjDskBxX7BWa15zED2Wcs46iGVTIvc+xMOkkSyZYe5APlS
MXbUlG1GIwuH9a6i0Ur9lPUm7UAqlcS+n8j+F4oXGTnn2RhTClhR8jnb4+nCD7CMfjuUBIE4VkUY
Ieecs7BbrVYzI3CgfA1h9v80hEHv2oSW/6K8HPysb4APqkfOJnTgKAXaZamJuTNZS3FNzWNQ2lBd
dY3WPd3tobbmyZoGHtmXAvkzbn+qY0P+yFhUhyo6X9SlM6Icwc7HSE8xpw7aTy/TOsDyQM6iSNIO
vbU6OVn0ySGudMBXcn0cDOtwsQkugdZXiaVqisB4bUtxqyY5rTIiOgaFuqHyI/kw4x8tFE3hb8El
8SvnS9tqg/XIZ94iPedUEetptTlNGKR8OUACJv7x1ja4z1IsQvfPmvUDG1igjVXWJRu5juyL4v35
NoS1QBrVNkvvx4nuDcdjSIRNt5v+yTfVTvsnZrof5UFqqMy0yU5R5BH+c0womLOFL+sYhevHLFKf
7Wziv7jj3SzKSs02iZ1ILpQLS8R5YAKG7UoWknoKS1Qckn08qgoW2tCeIHMdQDgk2MJAZ/XSGG6T
qDzvKDOZLMuXh+p8iOLoVS8bsASGK8gnrM9nEnwPZ53d8dXTwjCw/h6L+7KEWX0Bog5EtqYQEE6q
2Ak+wi5T1GXhtV8vkQGyJydPeN3BWC9CxW9p7XPJQfjkLoBtOGH7Otyt0ghQigChxY1owtkQpu8L
l/L2/3SPGTIbLnwv1FJXFA4jYEIKro9qjxq66fndmNXFpmkxAthiWxqa1FyFRZLf8c7lo5qk8U2D
RNYNhoR6qg+i7h7TVqq4SaZA/OSUuvFXMNh3NG9nx9rnmBWXXoSc9vBJ68lH6w1M8xHmgGUaN3Ff
mVwZhWlG8uF8DSncZ6xcr0csTdY1pDEwFl1H4q2yGnpnNc0nJx086aM9Y6e0RRM2hKz9deY5J7zK
8/BrNqlFb9CxKZayDGZfLuJfqjZ5vXoRlDpucK1l6Zp6keyq+e3x3ShMKxAGcFEDWySUyDu4txlI
e0yOUOEUpYcb0LAv8niPg71bBnWW9H6snzgmO47ziDs0VX6NHlXdVuZVjANEhcNGBT5TSU5/AAIq
728D5qRWyAVvSrLxbpN/QljkeFQ5QpRINqYNyJ/EbrPYrDLzJ1ciy0LyPH7VlpGTdxUCboPwIFWc
RRLHS1r1Wf/w+mMUXY2MSues+Oo+3h/exZcDN5qGpmMZEFsUBW0JUJP4JlKpXgtJrCsV+oyQvmVg
PUIIOHspHN5X76sDLLeWhYUZ+p4HELgKs+UvECYH78dkBOHM7Of4W9YTwyhnRaLZ3B2kZXPwqFhs
7/VNjqjmBYKlgt1r4OKAIYJglMjmY/xHRvjTlrZWQimquyL/Y/a3R5yrPAFfjQ1uaFNYbjZzdnAZ
cj1of67KYYmbPYDVsiBiJ6QNDwVmaN6R+SOkFhNgChZ9Kmn8E6CU+7sS4Zm2Us1oQaZi3R9Dt3KP
UFJu7xyA6EM+s1iEOnyZX71Oqn7m/7MDAzRdHWtO98xf2wxjXTPIByoqgd3Vaj+RkFobDsDdzIXf
57aZvfKOWji8REqXwgQkrU1G6+WYC1YpW1L5hTj05tlglzrCC+18y3fsXmhjISfScbRG5uImho3F
DflE5nWtoZa9q1gynGJo7wO1XVR1TQD+ujDoyqotDFelo3/+AqyMna5O3GYVLOp//iqJRez43y3u
JVWPkZ+K5aglaEkhtCCxCHcologx6gAzGQUzmR4dMivuJ1TTUajBrn5UmJ6EUrnCQp9XclEfFvIA
G0o3tXYbS1bdjlTIaYL6dw+sEV14Gudh7psEV+ofVc/9gzmvCYPQMkSs9lIsDLCj8Hs4n/Mk7eWq
hXpTYC3YtyHdqVnahfnJbsHKRKjfCaxR0G+zLQCJJhEqspJhsPKA5MArwT86jrzarebit3fK8dn4
9OgSzOWPcWuVuuOjfwFm27o8ML1Nhsw+5x17SjdFzq4V2COjdU5hHHcavEsAIOt3m2mr/jF5jrQX
2js8k+MiKBGyMxNlLBu5paVR17eUdYnwWoaQsZ4ozDBA28NnAEQi1vbFxXxgPolzYMoug1xtqMiw
hhBp2X/yc21dsHJNT0+mzYqqEZpFbTkcw3jbp/fFBGZDXRu9AWRswvsE6zUiYf5ggx9WbjReE4rt
butYuw9m6uYWr3Y2Hpl7/TInUzr83Z6iGdpb60tlsiCm/DrnvYs4oh1ocxPuN7+YqpHllyB3vHHt
hrEOY5yDcYWqDK+7muMFCW3Qa5zfN4Ugn9Y4dSAG2zjwO/rAMMLUcg3RcEUYMVDlPC3NN0GxC4/r
mbs9HSJrXgoUiE1JSEBj2hbN19gCafTEJHwIWcbDyq+pRpm9TQleo4WEI/ygZS6hhatHxagqt7aD
CgqngGMYlNtHgDb56Wm2+tNTI7/fFNDjdqNAEGwNA2AtEXt0SrcW+jjKCyEgVfcjSrcIfx9wfjao
i8I+6Fz/jXzIN1nBtcNGexiLBCOs8nv826SqJB+4Fvy78xGH2JTwoJxCypZ1cknsMyqTCx0+wEll
GBR/iwB7VlBE4xJ30maAD6J0nUhaglTJ89kTHWyXSsiPsQrpnOxsPVwjNO+2qEvC/jnEsxxc37u7
CRREJbVatnpTJHu2kIY3hP2cLOX4FDA86MSlqsWGkKx8DozKDjdmi+BUGhJODFet/DYOGeJVjc9W
uwMZGIZB1k6q0owhT3QIrEf3lS1hPSXNS5x2hGfGuf9bcRELmbqyB7btdOLRnqtL2CPRHRqxDcoy
gN7gxZzYKhJbrtIz9VZSnbYQ4X024WzkmRMp6KYZtRG7j+eYtQ9XZhIy2y66dAue95BMwWaUtDVS
1Pa09GlvqTNBKCsflhWLYBBXWYpoX0UuoPxoK0GqwrPcmMJOW1IwBh/Ax84DTBzu9uoBX4iPgGCE
JAv2vDyKaSJ/ZzYtVc4J72z+1Iev0U+xI0FKAR+Pue7vxa1/SqwHEFZ6f2QN4rKwhEV6swXGrlKS
d/Fi5LA25i3NjNxdEmITiMyGTqhIcxxboEVvHq6fj8WDhn3dvQzUZ/Y/D5WHatWoNc6o7hz/YaEr
HLmneCVrqW6c+27oMAkKsTr2J5F2qpcDdVc10mtkwdyVkyw2QwI0g7A7b0fckLlNTdwr/0dIkb29
I0pcVio/Ug6/23ZJm2d1Qq78gcSo6HkVGa/r/+gsz9Fi+T4N3hQ8bQRWt9uhsU1s21GehKMHZg6Z
sY0dpIYjvDZaTeUYDi1oYraDqtkseDH+jMkBsI7B49kN5YBN+VBqsd65wKXdvwI0Ad30ZazIOqjr
qShJbBz6a73ZQ/CuDdwftg5kRk/tM/uPgQoevpocdKFRRKGgnlLivaJxVq6MD13YqOlyQ52GcWhw
6RmYdYP/dFu21RttzJ1xAdpYmrEq+WeiRDv0zZNbEN/XRekp5QKr0uzyfaZPF48Jm5aqQp4OMW5o
hcle3q4pFPXlxv11rwfZPkof6PJLioU45DcybmumzwoyhTwO8cpT9dQqQeFOcIespyMldkNQVvX4
9RllgnEdMxUdLmNuDXe6Vaiq63JIFnZBcQ4V+c1Pmtfu0KLKILpbjL7MthiXiM5Z7IsVGaexg2cT
F5t8IJxa9tTzv+6lP+6+1FkpGO+MCMcgPLrhb8ItRSGIqRv9gAgZ5TYI8k4O9/8iaUSXlmHDOIhd
T/P5CweaPUjbvbuG7hS7Vc7zXaOzd4QYu1We31U99iV1NnPk9OzJLLUFQqZwQOKsosXtHEawGtgk
5ZERmPtQN79ZB1s6QiOxh5s07deE54jAZ33MJdMceDPCg1ftwHh7+BIDhjZxKpYFiq3pYgn+eHsf
s/59z1PgCuZGimvrQ9g87E/LntYvOi8KJmvGMGQRpyRm9ZAFr0KZQSuQulIPjQ9Z40HKSp+QjxR8
itIxYoegO90SzFbQ2jQnBXCSRNZUtzvgDfsq/0gdIVGUsb4EP6ZS1T0ngqZDhsFdy5AgxVVjl8kd
INwzIQmgi3XLe3pv4OV3A3957JvMbTfq0cZ4My0VZ0wKPSTaxgNe3NUtqjH4sPN4tN+LLR73TUOh
2V+Zu5j6Q+GmaTxet3xN7ATWqs3aBfDl37/TUxce9qpCfmlZIli+g4o82YtdYr7kn4ok8aax2hXa
gt7hWL/OF6hmawZxuNtxASNDpVt/VB4CsRPczZrp8R8QL5i22oUep8/bPeRBMqLcpo3KJYZ8XaJz
HlXRTTf8sdX5YXTXjfxj5h4t9MxKGu64h8SlC10tjw7us6taVKDaPwv0kqw3nc0uRK85PJSQrm4q
ffNRTytuosm0VYrBD3E7mNVQBpAUvwU9nSuB6zJCZoV4UTr+1P7qCgx/gXa1EpBJc90cpMFWl5pi
HubJCyYFVSyy6DvhlfAw43kJu6S1Fq81uul/UMknVXE3bcSru80zbezmvv1iFcmUCkC2j2uU25c6
bgsud/1J7gMqFr7kqETiTx6kdY85saqNrYBhEoDjDUQGyjj8BE26MCbu4HE143SA8joag4DaSepT
s1YFeoKIvyDaWJY1/cfQUuoCgxRocwUxtRZIt/eRadskMv0SpuuvSPH0N/vDTOgUbk7AstOgEH3I
rmMFnIcGDA93kT2KztJGaqmJSzkDOLwzwn+2n9rrVNSk+2vQHGGx/JZd8Eyq3r33QLFCeElflNLk
UWQ31H06e4kLIUQ8ZYA+6KiWuDGdhDcyKT36QFlbnhwbJ2w16/p3KTHkV3CdjRaiE0LGt5ht5xlT
mUZ4PVRon4Je7oEFZJ0S84y7Mwmn0KSOOlykZzdD7sXW+fmNRuqbf/MCjtFG+3UKwiMR6QKZSenz
3UoE0CQHOZE69TuaN+tf1M24xB6zfVRpkN+G0pgA1RVh7gEVrsqsLKWoI+1Srpo09y6YPgezjw5R
wnZaBBvq1FjXIuzT68pT2/riL/Q9fFN9n61YN99Yya7FSNa2I//gIdS9WOVpNBr3TOmPh7PWPqk9
kOQXOMJDegetUh9HoowizWRnaVClRG60w023+1eLITxkaTy2ng4xooZln1q77He2fz3yXjVLdQW0
8aEIsu6wIsd+msS605XyocqxKkmcC2sSm5wS0gQARBqPWCF7vGqtbCYqNLiPUyO6/Gl2Xw5NyfzO
kN3xQs4oVahgG6Njw9Eg6ljBK3BgvOM5s8ZnUCL9aGGBPA+XLM4nO8ETXbiKxQ/p5m04v9pBrDAx
mYyMfOI5nTYzxhzvaUpfT2nKkOAZLBX6BS8wL0NLyeyFp/25eAAzzS3adWRy2lah2SPAsyLlrMeh
D8t6YA5BHw5r8G+sDTYrglx/qW+poQK4bIl6+Kd9WljVJIm0Z4i2wgve5xpXYiJpCpa4JzFNRDed
l/R0f0GwHBpUY1YFWrqUcLyWJv8BJsan9DP2+JRu+lxy9E1qCDzqhF7RfplNVyE4xxC7z+rYcwSf
tJbNv0/dJ5aBS4ARfBo+QvzOx73zg5M6bZ2nMToEoht/gAGtPrAW9XiY6CSepPA/n2Po7lWKIkQy
2R7bUqmvj2/Mb8dIvC8ODHE1bJ0Ddd22Eq44XPmegk9rlMMF9l4EtHJ2ThcnBk3fStSHerkr1HMr
02z5oYT9/qQdk1GSaNcmhnOvOrA12TtaorY2Pa+pVDT7M3JyVHBuwX1J70cdeQRAF4jBm5gQ4uzr
+SV6H93S/ixRwTwTJo1LM9+Z0olC+Nc8A2PXQppqnzS979lHrc7LUzMS78nqyHTwLqIeMXOBMbRS
tEZwKUO6ACKpg+mljpsrSrvCB6OPMFkt84QxcdvVefUkWm1VFopdlk2S6zSIybHKgWppqSmP0n/5
Ct/LR4Wc7nym3p7CgLCJOoy2O8A675aZ8Q/O7sgcAVbn1LQhYd4Gg8BTrangTWNSQMo5AkfZoR7H
mdAEoTO+R65/yrZYAJhLoV2cVYjXLGpMjN/U1+/U/eg9fengHxzAaU3UGp0t1rpUnkdu2FSOFe81
LM9bBYUm2zl+SmsHLtSWM9E9+fNdbORGGy3FHiD1XzXt/GVu/KHUzF26/4fG0KWucGtpA1c4zPM7
4ZroSlSySTq9uM/qAJ0fvH7KeRmbcMSKB1z+/1abwcGrADyKKO/k7TPG7kTaEeJECz6rDIQnjpnw
bJpFFx97jjX7Pq3ahYd6Ezpn2FRtz36D7CkOvHZr1BYKR41o0kjTNqAQlH67QO5LTKaLif55weZP
ece88J30NvaaYvyUGDbruMI2oLbhRT6aTN7XAan21U7IXWm8srJ+nNLvrrTyOIGjpKctClReKddY
nn74465SNmFGBpuKSmidksB7UDNRfRcfmH23MRAaung9orZztOMMqbQJMw2rzgtNjrRrPPyyA4yk
5PIHKONWH5mKNjT3e7FYsndis119pkxbK3V45WXGT0P8y8BYxh4Jla+nMXJhL5pYRCMUwJ/0cA4x
nOSFr/bZpsvnanto04AxnIP9dAkDBY/8IXptYFyplC1IWB0WOrQzEkJhYz9BeVDbHXHju1XKIjIP
TZHzL+yzWVTqCJhCNgj4BgKDU6qzrYfZlsYzwA+Zz5j0nkd+jdAkUm/KS6tlLIrBqyTwUa4SRLuk
woVpWAq7kG+e5opya6rdhNDXH0rN4DKJP+mNZprc7Ypz43Nm+vLTSdCbStGdM/eyJ8HORt77FP8j
ActRENu0Dg9U3R7Nn+MUUiLkqBj3yWLor9MlTnzI2kcv6sXUp6OgutbzBOQkPACxRFO4HuadK2ur
AiZPSCovaRQPpe8wbqwc05CEbjvzfLWr62nIUMWL9DkobXBOnPVTFVg270G2Hv9gUcMXZC90XMp7
t9YLD5SDQCztcbgpLCuCpjL9YLatEQQpHG//9wPGy8MJFgabr/JUSzbS1ubhsyFwMA6db+cR2RNc
on95MMTbi77rIB+HlPWb52ovjnsnoV3T0hq5U3xywRgaZrcyWyFkIlwchiooDHbKtvs7l+GA0Wvk
vsER8FbsoAclSthhqLqHlA/G+rXtpHuXU3sZ9lwb50ECe+1hys6sOKGhTYedIDtyKaR8y5dBTU5a
T8NI0U40JKE4e0MP3tgddT1uNn4KXXOWXBu8D9qaL2eRjKHLTjGptB6fChpe7oIx1r5bKSaNkFgs
MKVgT7LX7Egxvx70BwiWTb9tknN208kEC19Y7rEgx6xwrdepheKLvaYg3pROaIL0MrsdmsiL3RTZ
O+dATe36dvwqfFmOdEYS3LOSsl1NtGhsUxSqDLcaKE4cfX5cG1Ba43PTkb9i44mQ2QwbTXK/hETi
IZPsmeiZ46vbF/jCIKUQ59X/JaCYrsgtVRqu0ILW83Bu22murkn3zwIbayNrD3zpn8C77oTTLpQe
lBihs+BMrhGgzNWveqVrmkhkGLQSh8npJdYmhLP0kaTBQpjFf6ISeo+WWPO3zVG2nlosFUr/ycnT
TSRjbMWDxK9LumK65xyLuReoNOnkVONBQJ+E+B3RyYrnCybM/65z05yHdhDDSRrTq0b5fUs1BAso
e4j1aP8MlmuIQJvq7K0w6JWP+5uqcaS1/muZfzGId9MH5WPFyMGfKYncUP0Yg5Dwli2UN6qv96Gw
E1jZfyvfQ6sPnMjz9JdvVEpAp7fwkrncC4GkTMVEiNZMlPG3Wuj9dPAIW7FpVywxQaWw5aGnb20K
7uKT2z7OYgHAJDvbiuWMn7fIUX5P+7X9FN1a/KOukDf5aAPu5a2NzYhHbxZg1YRQK/xnc37u5xDe
pZ5aYvqLd4U+t/fxWG+eIvPhcEWeb8ssI6pFEkcU+EPLIDHwb3rFvRddUvWvGUjwUuBI7J92hUzC
Q0vJxgYzPO3gcZ2r2Q82xTuuT6ZRxcUfSqPBz8KihzNo1OIzUGFY3I6NbQh8L55UzSWmHq0mY2Oi
xhKW9fClD2GFhhSK6UBpZpQIJX909NVG4MSwx8U+Q+AYtJr+yqzj5gMtFOr+qt4mIE4/p8++xulX
/XAo0At1iaKB5Y3B6nFibSCCApPL8gP+XLK6M5RWnnEoU40wtIm8+Eb/9txVu/ueT6b/E+vcr+ae
2if3aOqxUD3U/jyIGvq5z9EeyOXuKIbMDZhKrDqNpZdLrKeG643GjlP2vNpIbUS815wJ1hJSBhrN
VOBaNfYPG9ldx7UcDc6Ff92gwSSdsaLnkTxD7CJ0FLC9hIU5bmg64QwMTDhR9YHrvQF2hx/Lrq/0
/r+HTTyojxKiJqPw42noTZyoYTNlKIaTx4DUZl2OKvRBov7r9jYgiWeSo7VTPFi7/FyuI4lQxUyZ
sLCx0XCd8ok2+gMzSwgOhv//J0DpDgKn6Itbcvh6nfsi6aAAwTriuT9/xBKIKQVquWSyruWzGFrU
GFiLeBw89vqdbK1h5xAI7RFPg0O9UyQslC6toFabKa429AuPDQHsyhVHnFwEkQwgaqkR8w/fbCmD
M1dgRdA1KJJNaLm+IrqFnj+3u/ch9ZM2y2eGdt3kinF3ZYJBZY31TtL5xetafLnHbQ9DHsTM9wWH
NtRxQHCumk46dzAi40bC8YdrJPRICSoMiek0KRvpvQ+skn4o393/HG+aNu8l4xXiWL+28Khj90aL
VlEmDQzuzwJKRdwxcxUHO9xjVLbYY7MJMd2BLYKNN1UbR47VZRd+JeRzJDI1drPVkVeAw+8w/VB9
fD1nRLP8LBEElkIOykhJbXRl8dMSOkRSQi58RDCetdAiYNEQaCEzbxwbNjsrV8XeXx6aX6nwh+y7
8mLDK2zNxg1Y/iNoJ17buoLB7VoQonGWoZcE6yyw5vhaQWvmoLPI9wbiD2PPVFNQ/qSbhzpvDFj1
4dKV146Cw1y6NSAE7bGrkRv02kyYmESnR8vF4U0MB1D93BjGZ9KN1RIpYlqDDGirvCE8SVpV9JIV
K76pGhc9wIWMjEcEoktbqIwQ+g+FAPDRCHLJt43qm629v+dL/Pt6tbCLIb3PENG5/ah3gxiSXbGH
+B8PuNUaocvgZ7UehCUU6IM1PIAKrIQbWXZI0/Dn6wgBLNuUqN6PqM3kXieJ9gYOn6ImiNMiiOM0
ie/PA4QNdskU5HrsNLy26g7oZFvs6v93dpzKhs2PNMOGv4SbfVL7hAYJBcQOkmG5JL0nESdY1ux0
aBDm/zZatuuQ4gspk1L+I0Vw+XJ3pR8wr9eoZjvIwSThCg3xa1axA7PtNqKqejMV4QkPXS5/Bc6T
ct+dx9GBJFE+psZGrOrN51cxp8Azj57q/woy3A8aooezH8WRVC3QHkMlcPGQCu3vlhq70XiXxypF
kLAoFw87mM6c6xt0VDjGT0YTXL9cDH6pDAfreUzHn3b5ii/i+RaZ9NWeU6nLtNq/IZCoCFzd/3wt
0F2pbLd2GnwOVfZaY4YSdGQ03cEfUZ/7g0OAat2MyApX9/c/rFpitq78WZMqPkY9u4Sswk9Mg8om
HfTyz2pqLJejKliyCtjtJ9sYA4XRpZe4G01xMsY2+lO/vcly2GBtXIGYsMkHTbAFP4Tja3JyY8mg
lltJrH5KYxIn4U+VxXGEyPUTPz0ITTc2uCLLt8AfofYoNRNNiwSUWobf1t5ktm5ESe/gmIja/StU
nTHRjbtfxvdtpuBWu5orw1y0lrsOVwe7RLrjS+sN3bUhG8SA7Y3VZ1iT0q1AkDZciOqzvwtXw759
RoK/w8D+14wSGjEYHgZhFKnkEAX2TsvyTORx+t5FHDqqsq7AeIb6P7iusBpl/b9Ageto5+/l6Zjt
gC2qO9Dxd54wezJOUDN+i0Y5ZhXvn7hHQf3Cv/rJRes6TOUbwQkgmKxXytaqF53hibqwMtQiaBf/
hObo+sIrtWrqMEpANptCIJSNdCW6OOBvv+dvJ3PBDBkDvOEwH1wJDA38YHBEg9WsVudk3W1dbio2
dtCkP71DfCZzJbe2sq7cmNAac8sVevvS0WOMJLt6EEaBij/0PG84zXwUPApXWkaHHHVhooOv14d3
SAh6QqRuKT4VIJOa56Zop6AeA96LW+MO5QoDwIVmJ1n3O5akK4EirAZOJFMdD4jqBQQWlqp3yE03
wO1gyI1pcC3TLp37bzkypZEs5z2CGe3GBUSJOlNBlEe2Y8VUNg56OgbUAKdknoLEydAK/+x7y5nJ
08T4/Fe2lQNsjzJrFBwOIhl2jArt2ylyzYaLSh8m9JKmrQVTzil4YIM4VNPyq7gkc032YqC8j1Hm
nui5gTXKpU+ZhG4QpOFzYDQKe7qCFtTsE3aku/k2izgbBNbaiYNOVXR1vmh/ULFvqzdUnn1pk3tA
cdIceL+qd0zEjTl4viIa4yw1bV9mLIH+w7NamO/IIY4Z6haaFF1dsRZGNQGJPqtId1z7Jtq6Mgci
XQw10gNwsJoRigggEucZv/d5g1CdMf4VeGEHrxu7O9eSKFCkyoOID1jGNqFM/UZwR8BI5LfC4EdP
ToFLFP2TLZ4dUTTi1K4aFo1kct5w9QldzWHP8XBmX0ubLK7jYU44GDKsQGh87RaANShZGuriAru8
ydumgXutQAnghz8xvUIjAHLecG2x9TsswFkfkKqVbAM8sN3rmm5fFpgsEXqukzVtZrdvAaiFAI+C
xosAxUjSAyu+zfMpSkv5LJorg/g7hWxrVvZTWscRQqXTJqJeRy7PUzsNO2t4l1FdP9YWGhwWAJFj
AIPqa/v8dGY/TrC/+nYi8W5XB4zO7/uB7pjdip372FiKMw+0BJVdBG3IicO2nYIgAinJwrt8ftdg
LVAx2OqHxn7yv0mbWzLaCQh3GhxzIit1k+1h/LrY6xFMIDpQfssnrMH+8a4Jirfo1ydc/AG6uKHC
SJlWdkql/C9zJpFF/2vr1KWXbJ4u4UYXqY8dV+ZowWuZ0P2Q8KjXyuZ7pIWUSt+DRc9qi4Bf5cS9
mi2z3jP0olKAhkRZ8zwiwHLCrKHHUxXJ0zQDgqYRc+nkatAPbQekIQVyoBI8eqe9gDTJdcGDbquE
X9mnA6c2GGGZuoE6mJmRaN//k4tixPZ4MdmJ8zqhpfgJxTLf2hVzSKrG2yhVTmwon41AWcXzNOrX
Ef5Vn8unxquQorHNeES8brIFFvVnHa5DvegMAiCQBUyZ8gHszTtmTMYvECsDWMFReMZMasVFZ3cJ
YqzUOA0watYngxgCI3L1npGP9UFecfv1sW+2kuic/DN53by24Gl/rnV8jpL+lXO5fmitvPV0t9qA
UY7/XZX9fTf1AINaOEd+TK5xrAkJkdADWc/rB+slp6CuwDiUxmHtV9E++4OFQry4Wkg10XC3HhXr
ZQ/YHV4OxJWJRAWKpIT8qyPU5jNh1JpTTqfvP7TRUPti7BIxuyRpFrTDkXU3ArUCqWR+2cWfqDuE
ZHLyVttVKYp1oSpYsiZ/QmRXBOR4RweYkgsNMxpKGREU9hJqTjv9/3YefGQYLAfTw3mTLrrabUYV
RNSPThs46bLIEyZzl2hS+TIxfY7pKUTxjmmbRySu3ssEvh8PMpfakxHds0x3B5w6VZ5Cwkv8yGnw
V+bO28YMIn+HQatJmrgARJ0SPFBzQeO5Fo1d+AwZLDFmlH/4BWJY5pcwxR2TbDdxHaH1V9N58C35
afExndFpWsnpIpUhJ0/VlE8gGs+/x9WHZ2IsUwDvkE/QxgDFlDAvgK1QMDkwGVUzdF576oAo0Ec9
clS1iKidiuMjcuz0pfP7kCLtrIWpAJ9oB/ZdrRjltrV+llDCzPqvVl/lgTOvYs2nnWnjAv+HyXTQ
fsh1G+K025M6Xq4DAg0FId5G8xxiLDBlJ10lajO5D/5bcXgFsVRe3oalpLSvkm7BYzpKivJ7piGH
LzVHWamHAxaZABalIeGS4etMln4OOzJ2eG9l84xqUTtSgmOz7ZkgDEit6uMU57XCMa0Wr7IeZ1qX
d/Anqw1jF4/GIILlSUg5gam3H6hVMLym4H6Uxuz+4H2wVjYBFwHONwuo1pgGVOZgm7/lLd6csfCi
I/E3LMID5A8EB0TOsvp/DBbSRfLwNZ6iTudOf+I136eQTXYHMrlErkqP2j2Ontv8QXBr29EmHDe+
D9BlslSkHAm03LQCAyP0YtM3vG94YbMJALiF5IyKoUWlUhtr5b4f6G99B0W+0cmU1Qprz8EBi86C
yHnkjuWtgJFK7hp2jKbNPUEaDSp1Z2lvrtw/LGO12V6htNrniaY8oeDkxICYuvzLl03LY/mU0mJN
QOiEovS3D6XlEnBL9OfL4tNvfwT/BFhWKtCMaV7ZvXBYJLqqutnDG9W/0iM6W3eNOnZjYmeoThlR
j6iYiI9gEk68NnchqVu2T71pgG6teT/hu/EpT/kLeaGjqQ6DC7Zf9LwSj9sddg6MhHrKYTpivGVb
JnEAiybkD6wfn/o8LmRPfWk3EgRHL4Q1rtMn+u4Shk15ETLbh2GzekzIh37XtXrE4YMUwJGYVmjH
eHIQLrAEQhoARBnBEdRAaSCcnYlVjpYq356gX9g5vTiDVnc2z8/PRLSb2fALG3cXGB59WTlEPccI
imleLnKnzJN7TSaPnao3nFZv2rly7ELnICuZ90y3pmoG1LB377lYECMzDZYtFYNbERpbqMjS3lw6
Q4ER+c4cn29n6Le0Rp6Rb0+sbAReWiqnALAdzFVndjaYzH4avSJv0arFftkYt03ybokhqC/I9GJZ
7vDGD9Nf35nLnKmupnQNCpDs472pA/acdOOrktLy+b0SGgZf+/OjkNF/OzpzL1NnyIZdQMLNgVwX
4zZMI8+gMKjZrx1ogmeslq4q0wuQiGRNKE1hVvQpqd31/WhaqOU18Pd4grE5Zd7fwXdHOzCOTShU
xQyjhhnGpaIrMEroyFvrclfAaCxG+pko4RfkACysFWcnfRb16q29QwjIzzpqK26K6H9M49As4OJc
Rfm54RMNxoRQSAk9l/Fyrvhp16uZIGR50c5A4NB0LZorLj3TDEZWuBeVq4PK1xEpZldupD4XxhVJ
7lvbd+nBUKFMenlX0ND3G6kNYxtGuBxFiAS1QnxdqZt4/pxZaEA3njKk49HIUSFVm769pNFHq2i5
no0AP1GtwOFAf6tYC288BhJtDLXCc8/NZ0Lt3RU+XA3b+e2lerOaKonEZoUUnNNbjsUgU+HRmwF6
F9vZ/6cFct/89936WZB9Z/+6Cy2i/DO6mDSaZI6cV5MbEm3ON9bnCXKiksKWyYuQm0jEWsnxS3vu
ohHd4LBsxr9iIIuEjG58Rm60QytN4OXK2zgqF2SlBj5gY4cA7Leo4FAHXUL/P9CsxcZImDp1FDJG
rAzbvSp2hRyaEqvCjHNS3Vpe7khYST9YbtYcD4ktw8NYcNV+7khfD/woY3Ttcn892u7GB/WYsD5g
fT1M4fni1klrUw4fFU8qLBajaqKPKkjPBGYdhEY6BCdrIVvpwU6jt9pXzlASqDhw/q9t6jj7diQx
0Sr0PKuaoWZLyW6Z8swPyTUPU4T+M9iYRo4AdtxSceZAqLS7RyqBh7hy9SlI2ha2VrjjxhzVyhts
GZ+Tro3E519OCZHWXmmQSwL4LoEJ0PKgeG0S74+NyYO5mSiJOputEHlYmNhFDTVeWDZNFjVh1slq
AvcqPi0VadDDEXyfF4pHLK5rrl7LdGFYSKPxJl8TydnK130onGKy+nWtcGHxjIeJGlBKdHZ5xsKv
Rx/1ErRj8zxnrasvFVqz7WlYaSRA4dE62ICykXsrrTKyMGFyeU3ds7F0vmnVNVBTDqU6uVhOknEV
0n1t+W5WaUsH6NLrQya4SzkAd1B2ym3U9Yv9vhBHxvIARPeIf64qiMuBbLdZYeSYmukBID21jM0p
Z7PmOn5MpOMZRjtndJBCB0aPv0r/rPJaPAGqQCSAryufMp8ORlli2ZmhXLZd3S77Sc1q1UXmrIZ4
R1G32ItZJcJ2T81jkFVc9XnIi1Mumv56QgxDyRnk8pc5mJtDUGc9ECAL7rRyfgKhS2+W43Ge/vju
NEy1nzlwfALWtBLHldNRVCykmLOuqHXYz0DtwNUA5TVP/cjb2KB83mW3YzhrXEohWNRggczLCTF2
tNcMWhyRK3yG/uDy5u0ZdephdXv9gP+xrO2q9fl7zrAeiAOPXz1U8SoiRclXMossKKmTwqRTMYJ4
+7Ap129HW4wEHgU2Ahg0UbAuOH/bQxeplsqs5WoFVY0gxEzRIWgDQE5Sm07Bs9D3OiGMbqCqX1sv
GktCkYO9Z0DPj0M5CL9KvWWjTt0feGv9jAuEGGKsJaaOQ8BJeIHczAc9L0vKjKT7f+6kmtOgtgfy
6mFurohUoGd5ysjvWM92eQdSXMbt3xcwZ1v/0tjjVFilYJGnjjBKbuvs/vJHl7AuK9UQl5EGn/yf
lUal6chILObeUjZEZevsK5olMB/ILzlFWI2cCeAFNnp3nX3jfzoz38z9OQtVt2/JZvgxq39v8Sj4
ITGEbnDav+GvilHyqe5YFRt2XnlELrOdQGoGShrBgehlWyLIZJzSoc9Db2tSkmQrpe2KIS8hJtqA
kdOHBiUHVW+YxnSX8197wpXkcZ4Mo4hdroVnSzwj4Gsj+R7Fxr1bZB1zrfD8f1GV6/X2KJtRNsdk
jhmeMLT3gJitXFt0xE5DBYzL8VVUZZSPkaPzhOQxhv8X4tOOPCpI4XfzED/8jhioGE+zljnSVH4c
jQh2zrnTJsOXBOOAM1VAquWT31r5toiZoh2dMabOsS7eQMrHofLG3sDGAAWXz5xE4CMI892kDE6Y
AK5tfzahS4MuVimEgCoXGLCgRI8T74TLQRdLCFa7RwJ7meofwBuVSxwi/NoDwI+YTQk9zOPh2RlU
Pw/oWw1sOKTKvKzzdJNYioQWbmbqupsZtbLpHfrfGhfMSqLWhOU+q/mNw98JfgCNBk8oAGyJuuOt
jSuFEI5NpaIgBUhnjmuOp6VGXJaauhmVbJnoZ1WchmKsmFjAu6K1KZ8DiwINUzgnnpxzgXpsOhkr
fH3zAeBMQk+3bk7VNbiYIoohDXreDx2zPRSCG5AmxLygKDJTP2mL8S8B8XAuVKHNOyCo1MSiGB2k
yGp+d43nbtdbGCNo5C8ncJoV2rxE3TvA5YD/GENyvJJcPrjo9qeXufJtgRU46JWxxSOZNAu+3b8V
IW+9T9m79eoEXf5MeCfJmWWPnE7TkfPvMkms8lAI5LPHhkFZme9yLWr2p7oIxMn0RpKXofZxQ5uy
quo7qC2/WiC3sbZc5HXdpSYJjraQH/pVIfxgyvsLVNgtNVKFPVCCHkkAXXEjaNio8NfSkdbUCZA+
jN71flB5gCo5hcveKfIXl87gl1qSajYKT58FMrbgA1oTS0m6i5pVM1W8opu1gFxwL2Sj97n2qO0b
pKOiZqKvq677c1o9DVkfXMHZEOH1ct/rZNEP/SY2kVOjALLGl6guj+F1ipA0yL9W8/foeOXvJY03
xFLCuWgZMbuqM4jexk50EbLh/ZKGNfvnBfYydgmR+1SxVvg3p4/80301N/CtGDU44jBemk/zrTNQ
0V6MLKvOUKJsDdU3j3e0IQajSTgpArDUeM8iY5pqXGh4UI7tgJgWbklu2+onBWlbQRpY/zPceNRL
r/IJ+DnqxSz5RENTxZATBCj5l0WHHlnBhFcAPnYsUUBcmM1IJaArzcYUa2CkRNmkVMg4Pc2fvFYF
GBSZ17OeETYSPfgb3XFDbNP7AdaU3gbNwYpBwxWtvhglOxezGVTPJiDQasjUF2nUMUmpjTZxJjRi
KNgl0dGou5BprFxixHVRdHR3qbIZTVdCSXii6tditBLZDt8O58AEAtvc3hSjcAT5qIDZj0/WmPHe
jqRBtsP65/EDRnGEG4EWk8wRM9VGLZK7vVXvi7+jKQcjf6VRwqWp8zN3fFjIBQ9GxeDDnf8sXrn2
e0uw6USa/HmwCju4qnFI4bbF8IUXHXW6V8eV4mQ+qOgoFzaj4asWff0bW+TOGuYOSbXT3d0Xh6RV
Ozz9wJ9dBDpUP9cN5s4nvtlT643Au/5tJfraKq4kpm6MbUa90O6J6paPUYFbuqBIIiNzbd6gnLu2
mhOzTZNppe7PowKLf47rrBwuCeZGrmUJhY67K4GD0PjMc/2dCxt7zE6Oe2vO5En+PT+OpuwrH+3O
n64lM+S3/HRASVMW/l5QIRHVSN/9hwf9s0znDnzkOJ8HrOf7lJT0ZoQ+6bU9H9iJJBTacfk/2Itf
clTObeZo9p9/+GN+vDt3I4mYbCFmukyzCjgE8DpEQ0fX8mSxHIHBiKQUevaQpD1r0/qELHB0GO7j
/APxNj+sneLuVjKIkpEmmFUthP3/SFi3FQvHrEvwIUbv016XVqjhQTI/ydc+Yblng+9r3B5iYY7B
C5pF+AfIN8NtE+XFOYi820u6Gh9h2D0gqqADGDepDyEdFmZtIDnkm9Jr5vzoIi1C3WDUd8UBu7Pg
19qMMulZlzAJkXfi/RIgopU7fwIFn3k6DjedcC8/RoOooyhKheFR5DkUOCKNkve6+Z46w/e+aTSc
Lw0irzFYJFIrwYKZTZxEQ42TAxXk2sQ/f0fTze/WUA0lzLVxsPubifdSsiRrt2PrDqxFvAg+Ux1i
9HTeP5Ql9c2aJYMLutKg5jhW9lnVL+L/UDNAIO843tv3FSqnQNuxjYRGrmmOc5e6ilz1Vn0D6Fyj
FJPdQrTh6AhmLmYivqcyai49y27Ftc9D+EfCN3DI3HCEc+rYQyOmwQA96Bxxu3tzcLt1JBko1hWK
DLCFnERK8aY8z5KP5l07hFUPbJ4tSgJ1vo8vj3bf/JZD2LLJ9MQoAtDeNTynBAxSdEL6hyOFwIgx
Hv+L0grj/mhHfXyUP1TcK8mIOIfu0YLSQCBer18Eyt5W8h452W19074DQxE6tkOV22RItgE4xyyV
9fyq/ORJXdmXKo+/gbMFqmAG/12lMxWQpZUhaZSZKqBSrca6wfSgWcvmBFzOpHnhweYWenPAucGj
JPPLrt8FAIGObovYlYEY3Lc1l6uu83z4pbn65m2+0N68fcAW2ia0wYxYTEb/j+os+NqmOmrbl9o4
Wd2UP1dpTFg60DO2zZhbB0Jg8HT5n7E8iEZ/0kt2ZYzDx6cIXgblpQ/ytEriFYScTl9G0pPXwK2o
SSMMAW4PU/nIsbY2ywYap23Lt8fBCXNnqNH8ThUpamFPe8qg30RuRpJE/38J4G3ZcwcTaZESdbs6
phADVRCeu96hj5197blLI9vWFpWor94q5f/lG2knt6RiyaxmwBBt6sDak+o8dYu9tWkRZ9d6wtIc
hLfYDWeXJqk5PW3x7/cE4bWqzGLmg8CUthM45wZJi6M/DUF48gN8ry+pF+XsbmNymc1uUG8iX/f1
n/aElnhUfb/5cfymw2hAPickB9nUgajzxRNelYlvcgTc4PnZCUmDIn/CeJapGgMQh+Sk0SYPm8Lo
5sFoBnqqF0+eU27V61c6bSyD+03zFi6AnS6AlbshUDBbkD4/nEw7kpSjgk5Cc4Oonmpk3wooA9ao
/xI9O3ZOmKWyifE4Kk0vSL7XyEke2ogmMVNMcGUCkKD7e1NypjUin+j7F/xK6eUbNVZizRRTGmQD
4MiYLCK3/72b0A1qlKpp7V/8sulYTp/sQzy9xfJmB6DuG5+h40kLC6VHfpFWxYRHxSjQkQdSZeXI
ZYdH6yFMMHMXy6LiieZqEuM6tNAPyv/O9uyX9uLx7vCl0WL7G4VZqiu0dFycB4IzWmWJWzKhH6it
PuKFRXYClisvEEx3HEN2c78OsTX5fHTqgHE5rr4NFMFrt6JSQSucXcW8BfaQVz+w6Q6WLd6cvWF4
6LyEgk4DbhADvLQkCkz401v2bGi+b2QV5r4zsF/diOGSV022NzkcyHSs+YcHOqngquco3OdRMCVE
2RsfjNMhQO0XGMOUhmNLUqfovNSEXASYf/zR5GBRI/34Mr8IFUUokfItnmaV2DQNpSuQ/Brt3XlJ
WG07UdPO6LxPDpOwi48dfFF2ytE8gr5TnN/co+uUgs+tOUN0YZuRkluOcjIhjpXeYObxm8mqWWyL
xZ1wz5T8iMkuXusMW4AenArwqsHNZX4QXtCC54WEtxWcvqA402wFUnrcuS4X1xMtA10vzf08SrfM
QAufYWMPIh6XacHHFAzR1V84IXPsJZ1zpSnZX1civkd11mcPLDSqlaIkpMeYBNNRwXZXV8Z1M2dJ
992ZyebL5MuSPQHrZ4PF5MnqNAc5esOwlOJyczArI7b7CsbbC/qoZBMhN8Z/Grwb6kj9iOXwNr36
sCzRvX/10sIs9e0YVk9i0xDCX/a7GyXiwD9oWXovr4Z4RubEAV8qgEjnBPr5pgk7ythz102U0S2q
eN8IrSG+qEEMM6+V6cz5UiDDHrgh6ZEqnGtzyxdFHv4kddglas/eO3iard0CrYNSHxnHS6HkCk/e
DJUY5fHLSoIerryOS54G0qQ9Jwr2bjvEUwi8VZ5UYb/VLW6MEz70T0j7spEb1CZ93IGPU0IhuLn+
0z4DghtfbuI8esQivhezfpiRICjTtsssjMV2GeXkvbg1nhhehucXjwTClDuVjtX44TeLXelWlwza
4kD/4RCCkQbj2fV/ueMCzRzfEmShB6sP/q5b0g47RMGwoMMcgRhoL/NLmofh7McZMROn0Btp9hWK
HFubZhXT8WUkfc0t6eqLx9rjEokDBW1Qv2H7MxF3psY0RQavu75T+4c90BnEC8wp0urv7gmTfx7B
oAgjlQ19k9V/O1sj/AwlSTje4BjqPhfq7C6Cwxz7fbxt5aBUmt1jbqaxRwVGQb9aY+wb0Pt0FMg1
4zcXkrw5HygQpUFn/y8UOSS4+GakENS32FC5IekgUxXnKg74xHQkPaj+BXsNOuV5TQIuYF5ifRsR
3RDO9fnP7k3EASSTZzs6ZOI4Sty4fzGGe7WK4hSvLkOmouTBbkT9gtaNm7HfgmnxfJbaoVkPy80S
/a267LKoZsUZxQF5EWryMX6WeCygdsoZt/d4zj9SOvNikZyQ+KsmCIjFCCbSK7QuXUa+gxHvinOP
2TkR5uHyd/8hI0CR6FbFlGue4e882yq/f2Q1pRZIg+m8z9lHKZ/6LH0C1VBTG2ShQTWj6l0KqCV8
xQ+ewr+zMljJ40LCnvAo5iQB0UNB0GIOAyNnELJ65I7Grx+DQ/QomZCOzuoe9Qfwg1F5i2bc//rs
5hOZVnD1la+hJzqqEuoLW/b9v976D2PpNynVSAotsOPb2S+QXaISQhZYix2RNbkyoVE8N9FUvqXH
kRWF/edEk4FC/0LTqUI2KTEapK+hFbIs3tQwWs+WMeRYbkLR/U61NlHUv4Tm2SllH4+Z11NUVu7g
6JgtshTjWNUsy/kxJmYhKLk2zDYt5gUcowOKoOd862+6kFPXcb0pVudcY0Tse0/9kwkHn2G+AeaB
ZdBepS9a33bdhy7ykaL5FS5bJAq622IaGip2gqdnNlu4FvffIOijBSXJ+zSCFRDPUYYBILciNyCn
cs19xbJc0YAtqoDgxqGE7d3bH9l7whzD4OW8FxwRUAP0DucKUODVLh+ahQvAuQ3k6f+YK57eKyBM
6mpWN/GnmIOIqiBQ//O8KRxc03PhD5QasCttDDrB/ryq6NmGWHxKrbYTtzhrc7NB6TrJP7AMnXRp
Dcz3dgtozyBo7775Vl2FrJL/YZ+rDN+kPSIKa5KuBMPvsM1ngv3jSv1S/RDDYIE76Pl1VNK0LK2D
F2KtgY3c+m0756laWhAgisJ48Ra7hahxHJ5Jgu1q3TC1kSH9ayRd8Dk34mIN467BALenuEDpWr2D
GTccnKhUOMgf7GAAenXCKXbX4lSKxpxb2WnOML8UroRqt2Qqv6spcy3nP7rcmOVQmBX/QenS6CiG
C/m7xoeFujXtR56fpab+QuCZA/Do2zhlAQ6rG+zMtxF86IFW78fy9xZTWOx0GBMGio71CvHeXZUY
XlxqR2bsTncndFWFViksAi5HocpJrigqw2oGJUpa5Oh3DNyWKbo5qamU0oNm7pxdnd6EoER4lILQ
GzABLTeNXDEBD/TIWxTK+bL0TSPfiQLOeo9WBSsibnQy6kmHErshwC601ou8E5Y6kNDy0vQ2I4Ns
nwhUfWTgLyDjuoMlXnD9FAFig4u63koxbYP7g8CZ2BUH7jZbcUVbY6IFNA0MNXCtkiCbl5S6R59J
An+HNP+Y0f8+T3/koRvnkjIsV5+ZL8bRVkgrNjy3F+xVbsPNBcdg+n5xk1dvgTCNApDNzh6/0qGr
B5lTi+SusgFr4HMWpZXFoX6XVHfFUgNdHiOODGQZSrlSzHxG2SCUQAtBhrJgZ2SD4KeksBFJ9ZS+
suGEy04oe0CndcqOzEOSULw4nLsTgp0BdV0/dWBmxqEwRB7bsEUzVUVctIdfauTrzHZ3VGWGrfj+
9BY4Hr75nSJSo2VZ1770q1nI1cObn1xLOZpqEiq+vbQWf69nPTKES1EdvxV0/r6nyICURryu5n95
qV1xpKCDy9zRAoHOGVqbT6XIho3E0YicS4D5ZtjxPDfG1cLx16DxKwTCzJ0mPwHmTATGUfuLmiQ5
LM912qSHVuirGFL7bmy3vWtBi8+eXQL6L++Nv+e8wvfPkKUh+Z/rndPObBWIf0DTWSqBq4pKed5x
SqxA+zRQtDLWU4sgnvCFQD1NWUEHBAvRiqmvlbo674kG+oBhxGPe+ugqeEx4T8Y8xFCCdiaNePVD
DJINyFOx7sKIzyUnB22kRBsxd8/wfMXZOK1RUr7sUIitItpJWUc9ZqeIU49flWqgqVoEqW0PF4PX
PqxjDx8kMgO6YDxKZ4hGBkq6ypiGTi42Rkl9Eo8oB4bKo6MuV4fvdSMoC9m0ijnjo/AYhExoZm+O
5+Pud+kqb7+Hq+nNmuwgCIB3Hm7XkEHTaKeFv9qu1Uqcr1+uirMxJL+644i3ywG1RY67LLWHuLsi
U2ddABOkHxrLq1SIzDUgZjewSdqN/MLl6BfCrS3z5UwLPhxNhFbIO10nPLggsUpiYT/W/RJNqMgs
SGI7OgsUqKqDPEL2ONo22iTzqphsB3qJ+WaK0sMAMYibige4/DOQ19tUU6y7fhf0DxlFbvbIquq4
lLS7hO6F6l3CN7MKukbRitI+vcdG+YK/8eTBq9KyFuaT+eEnuP62BeQ3jeo9y6Muihd6RylLy0yz
4B+ZPSeswYI7l+ayHWZ31uRHLBQeG5mrWMoS1GODCSZS60emNMvmEPqpfHKzff7w8orIMIku8jzu
j9RQH3o5EGndAZ/npNoaN3P2OryDXYaWGRGk2uizYLTzJy1qhuYCDeRjLQugdnYLIoWW+WmWspA/
zT0i7gfBubBYt7lvH6qK9ubjzpxqS7gcLCMGfJIUpHKUrcwDle162+tdTz71eT8fKKRuyADhCmgD
GxDkS2g8gZ9PhorbHCjcxAXKnWcc5+AfWpn4vtijdxv/8wHANWq71Tklp+0LMAH4oHGaNoxQ0z2L
JBpPfmyctxCRv3xqUvg/U4KMCeT+5YyUe5HSvWi0lOHfsOxUdEK6o8bybQsX0VSFsL3Oa+Hwv/Sy
HyM57prGCqUjutjnf00hThVlI+4rO12HWmjh55KmLKN7pdqbblHiEwXGSmeY+hzL64HvduQn1EWi
QLYNPjTaG508Unir6tfoASgcYGSbueTWgf7+Tt6afaPBx7NbKWHslacD6DAGIkEi5TFoY+9bXIg0
KNOCPoGdCz/+naYhpejZfStQV6h5Nsz5nMGkJC1PoAzxHji0T3wrt+/dBJc0cJV2sxTAScxpUGwj
MJ1eFA4OXq5pjF2K4m0MNUiPDn5WyQwKUEWRjDwotspUWP6gRW5MZitlib9Of1cCNk9DkF6q1amC
K71ceZTbER+3gvZr1gMSH7EoI500/iYts0+Bdv75voAZo0KLzKjImRSM9cy5GXi561i6NmQ8mT+o
tYcVibsfRIfX1V0zMmTM//g12pKLeOMtTscZWyrd6JLJ+D+UtMFQ06U7F4g60fR4LXSf0GGyoMCM
FnM6gKYjLK3ayvty8T3BWv6ZOHvs3DV113bGFaygg6BzT3ewppdUipO4LX/DIS5dMZ2XZ5+Ic2w8
oNezInrQ7PCGJAxfB5SObxOevOH0mquSDXMSuPeOrRSqj1WyZghMg1VlCsWTdrm8u/hN6W9ZXUYd
mZ1AVP0gnJ5nCGk0miirm+jdU/kL++AKjTDO9zv/AOlpr/U2nsTeky9IvPG83vC26q8seok3a3xD
n4u8dtKv/IP51dmn9iadBsdYFsEXVbTY03r8LB51M/K1m59AG12o52WJ4LYF59iCWa1xfD6X+CKF
COYgXRH9r+1uTXr2S2FeGU9KhJx7jHbhhaSCstHUjv3b8k9QuEpaoRyFtWDDCjuLVsVxBXdKLlLH
/OP0d5+heDHWgdi6bPIvtREkOMBVkN3qD+bSl2kI7Jjg02Ya5TTwwIQ4+8fhC2uLhdAHQHzHG29f
fLymdnDphAxNwsIs17HYR9GixOuqF6mafI465oegV7g0JOvVfD8/D+/2FOuoddubBmr1X7K9A8cS
PJIGfb7iAU24RRUu9cdyfu8hMgbabGDCS7oXq4r2qVvUB882cr/z0SPBtAoeWsPzo4ZXWbdarwB1
mWLwEO9Q1XyinU4ovmoDTCwi3w7qaqcizaRgG0NKeHOXckDbxmX0Ic9cmuu7dK05d4+Ib/9gfveL
Xr+4R24zNt32KF6V4kegFdXVmJGOpzj1tRzOolPj5b+I4vYwyJEnFiKwacI2ABVcu/84FV2ILUmM
U2qO9QbV2Et0KAX4cDvxlHvuxp78GGpTOERkjdXTLE0lmLPTn6z6GmUgYUVAGY+qC+hcUaB6CtAx
7Ve1jn8Y3dx3Ru2j9rg1hn7g5dH5DmwWsdqNlZyfkaPOYxTMBCoeNEjvGBFcpGitbnAw2eIOX5RF
VlO2nF8LOxx+6iF7UsAwK6cxSyPGmi6yrLk/rs/vUq0dosFvWZG4ZcII6RS64lrFVBryMgs8XS19
efeB/JC06VnFNdWGdWtfdnNvwVabrP26fx3aDxUeqL8Fomacv0vwWAl+VmfQCX4/JgxlXSNKo7M2
DgAXLiL1t1T6Jl4xieqJpGAJodYh5m64LwR7nrNzSJADaxl50iJx8u70P4YQX5rNWEcikA+mhZDi
11hoPlR6zbg4EpWn2ZZtX6Bexj3qeGrBjq8SrHxy8CfEmXIjNYzQEnlhE26hXOB1Pn1QXuaQS5M8
EmrdJHyKhKV3BPx2UQELcifPTmFRG1KuXIYLpiB7nIaZNbf028oxyISkSDfIFuyaCAId8DcUR+XD
jTAA/qdSutyDwF7PsJZ1LLWFqo7GmjmN/c1oEUJufAzNUBsjj8BuxM0zCZ2JcPvG7Mtm0fORj2L8
/w6uiuSHGJSSEJjGYBy5vJ+eywragQCy+syKV/12DhnnVfjr59PjHdPtwUbYZPRW7wn7cDpSg8Lc
/e9YJVhHsWvdoYRMWYDETSqsCw2nP/nSAp2ndBqb5HM2gxSPhKrkkIEsKnEZDpiP+WwHh8Z+lT9k
dk3Pepru3rfbzW7jKqSJlbgWjyiE6k+wflf92bgEGsD16a0chiukpAJCMSF7S4ndBTVMi0aihJZt
E3xUhGIq1eotPgl2nk0OqdZvAhWjeyzJQ64xqxogeMMSKe1vr8RvS2rLqyaUtYWT6/F5WqoqjP7/
eC58YejWTZF25mLE1eiYMn8eR/nOhhb98nJbq9cF+xw9+0lxLdqPCOEKWWGGFfLPA/bU2bub3x0g
GuwGHE4QDgHV2XoM/VCk1PrjPGPlNV4q4/hSY6KFL2CzsgxZle/jX87cscpW/R1uOOkWibLFIfEZ
PEq7nZAT3IsabONRdtWMvHrsTaqGii3k2hTUbG6heDrr20pkosBu1dAZOBrhu9QsEg7AlrT2Drve
lWWLsyRBzXEkpr1ovvB33wlmbJWxXwwdF6MJWrnVIPQuawvPj5pyMFxBizHG2QqEkRRa7rRbQ+Qh
b/b4oiydteLyBs0GFqjpWAQJ3sBtaPQ6aIDk1mGeOPgIJtezCpuQY3eJnHBWnXsG3zAMWYyONX/n
WeX8+9s3miCtYawjFeejHsTn/vVKbyKyzUqmxzk/2ZHm+JTfvcACz3O6C3cgQBbFh4LFqzDqlCvE
OOqZ9Vqt/m/eZJyg13aoRu0n76s2oKKmbLaTQ36gBZHQEFaYVuxEGh2jg4XUMJ/PXtCoW1Cq7aAN
iE+EDtFosxSHOqm6RnHYtP71Ohb1aUHSdEGrNdBkhOWvkynWyA14FMMTRmUPmzWDqwtQj4eVL+iF
SQcizJGyblAYrTFTxi2tsIk2qG+R6GfTkR+ccd/K/lGs3JHWmhcJC0Z6jL6KYGDxh/M7bbr7OhbG
4ctfroZdRxgZUADXzBjAZHCjQwDG8+9TX30t7i31cLFJ1CSRafGlFYiFZL5X/n/HRX4PYb+0DQ6E
3AZypX1Htscn2JJorC7/t851HQol46TKFfrqo/nYqCQ4tOlPdsokpTacCY9KexxLoJhi8gfmqFJp
kbEWiTrKzxhfXhw0V3rSoiunmVJvOoJHCKA+9uOUs9qvSHgmCC6NclCZ2uFJ5mug2cQ6sFFy8dR5
4cKZpn8eyTE5wEfDVHFOMaiq5vxp+LA4U730P+Wf90rfbIBBSkWCueAKw2LFIZviEfOrZEQQw+Zu
1sKEP9eoyU8VH6qa9/Ysj2Z7C3YFRT17EbZKVjDNuJ72tNhhWl3WiYE04GhNQmmShj0f8EzNERYq
CL1l3Pu8sjnCInb65bN29iKcOQX/eTM28ZaZsVdUPM6U+u/vT7xNgQmOTEavxh5uCUTv69cEye2b
HCZYmt2EvhJkPbNiCdSNdIAce5jhmf52P4t2tOZ3heicAKE2q+G5vhTCwxMNWpUeQi+eyiAPpzAM
18Wt86Qf3HIr9mWr+Af9TaNHnXFOx/jwOZzcN1Fkdum8CA4pvHQP5ik6kUDaTAd6H3o6IP31LpER
09v6iyFaadVtImWZnvgsHPYdyCtp0XI68TozF0ngKnhj5EoCb59l8EF6gu2A94zd572Z3wrqQEwt
Idalcxr6y+gxtLqBHN++U1szdUAkDN4Es3g8QkvQMmNOHSJERhFgf711vlpcBvkFKsMzkrzRPnh6
YrxC0zPI4YO81LUFs8LrEDFTUKg9dp31/fyCs9UrzzWIH0LevPxcGn3WHhQ3CI/I/qXoI+JMVVbD
7QkxXlO2QMBllH8t/5XDKLGTrao9d8Ye9p9zYHmniuYGe1ArlOEp4qin/i+DQg2dyeZ8n/A0ujvL
RXXvoqBhCfGO1bqnabbTyBBSnEtWa9NBgMYmQgGmzGZEx+UEWJfzplv0f2qmGq+HHa3d6Pndl1NT
nptdA1E6m676vCfZCrRNYF7Lom3MixNmvucfrPWhh+dnfUcCL8hEK69hixt70j0HW9TRj2//EyJ6
gFNzWzLr1j9eCIK9ivmwsFxpuNqYMSgIJ7fb3qaDyXK0M1LAUXMBffKXHGklaLOZPupyeD0UE2Jd
GyLxQQSJ7Y3u64+uLBLkG5WnifzamRFo6deJzVDToLSfTm5U07cFvA/Q37LGSlH1ZLIp52kfELHd
SLIikJpytEd+afJPE3aBC9eOfY1DymUloVsKic0SjgSiEgs6Nlb7+F+l0uBLRrSYUNc3DdGnFGTS
/BXkN0tVKi5qRmRINGvw2kY5JoF7AVmaJyNWhcRbNpd1wnEKl3Q/6c/hPU7rCD5h/FzkYfoweLiH
MopFuwRdiq1uNr59HpP76+MT7JDNpcxydym7bP4qw4Ljw12e3k8qD9vpSDQW/CA/vvUNyHf5HjKh
w8rI5dTh8hcw8/wWS3Aeg4Wl5Y7ZCQ47f6gvo2/iJG2WGYVe1jc7MmnjhqLFzn4GGCPO4M18zaH1
i3eMlsYVsFv+HC0WVzTHbD4A8azZLu17D/0c15nD6PFBJh5SbhSZQc9i1rKmUHndLvZn8hwPgkeO
6DJcnDYnxdobRphTujj4pc6KiNt2ZfgcCfK8U9G3gTjzUkkKPUrrmQfnu2XpRLv9SEtstfjJ619G
IHO/RxE4mm6vmN36PHL3pRd5MxTZYUj2EWK6ZkF9W+1duRDadq+VyvT3UnPoYm5+8OgLWwX8Juie
baDSWSPeXBlBOrAaJ3c+63ddRewpKpBWpSGzZQTCXKTl+z+I3t2kiEmv82SKde6yqQfFq3A4rcOX
0w9dqB4I3naR6d7o86KN3pGgopFZCzyf/nwAzetUy8MkXcteLSWZjfa0OJcxMdfsOyNgQbr3SzZH
0Hc4rfohb+LRbzHF4sFzIPKO2YxuhTGwlDOw379zPtmtOt4Is0x10T+MZd8dIni4gAIY6E/EyRtC
fDMu9Q+cNxnMcHWuJV0iG+87qjq/qe+3iddczM2eJhRD/f3990Y1cVonc6sLVDU0IMMkxRxHWzWy
SOiENW2b7PdflInywucjH3/iBwmsDMqUWkI45dXWaPSqq1LmwcWnPHU8zEMasrnV6Jm+/vwcNo+b
PMWBb1TPosXXhQuhaC4iWA3jSFKt26T/4ncAfHAZDS8NBXnQbLlSKr9h3AT4F4Hk4HncOvSqpTbi
3wVF/oUnEH6ujSpBHfxuWrjV1aefJ17w+AhYMG9Uh5VzZbBX4a2D0g9nX5RSeV1pBd9r/YVK3Wt6
hUViuXIqquL8+iY6ZYJNN8nNxgZpCxyxuNAtqv85Qt454Pq0IIREx/2ltPZW8A14L0xOBNHb/COs
meGs3lxk1SfLgVxkWgRtvOBVcAsQcip+lJo4XWQv71ppLv3WKadRo2JRbMp6NZ9+IH5awll8yyDq
NFcsBr68WuclXonAbV9eEPBEixXsmESHpO0HgyZqXp0UZLmC4CJJchlB1ZnjAo+rZav0pE8T/pfx
tSWSPTzxoh9eRPm37oApt5K+nteh93bNFmHsRaG/aaGFHdvhT3vNeb+GMPnIoTfrupYndoMpDKvn
k/jBYK/sCWQtsNpYHxU3jhL1R5xXNb3Xyl091yV+hZrePTgjudKKulS4BJ0rZQ+e0RnVK066iln4
g4B7Dlfk7N4WwIiso2I66+9RZw3jlPK9zBw3PeWB+m/oJ8c2N3tpXiRpz5u75NM9ZhTQLaoHmhY5
BF8g/jyxOZAHj/TnYLPwZEHrUBp3k+Yk1QASTFOdnFDGv8LskxYSs+9qICi6dMNmoKqHkDtGG5Wn
JE8DUwfmVTt3ceHbUMGHS714QBQ03MeDFQaY7JFvNNizrs4sgnag5BxiA5uk+6+oscH6nY5wMkCC
JJWZLFimb/iZnndTJfReg5m8wz+nI7wqe1ZlhJZZZcO4xLD1prcIr+7ETGpSOz6oirKh1g2jf16W
5Z0CSIUUZXVawZYxVX7R4GiLUB91+oYqSTc6NUVd+nKELL4KeHb+0ao0wvIakplV6vas6RXRk7cM
d1L+0NkW9mi4KkUH8N1HZnPTMivJBaQE01a53gKXrfZizlemNfSzR6R5CVBFHHdAJShwKZCh4MkV
E0SiGezZRmsWn+02plPB+9o/jSrfAZclvb/dGdMhG31GiVX7Hgi4WQtrIF9Yv6wbVB8Gw8mhQsqS
t1aNasLiDARaIEV1FlON+AJNSM9rc/RqdQRNJ+oKjGM+QSHf3g9y2+9uQlWEK7uCUlGxaKShyQEf
/JbMMZ6V6RyIOqN5F9wVAi2wcJ4F0EY/sX7xuV2fau8spuEUQoyyudreb80W3jZt9DpyyPoVrNGW
6jOrKG9Gi0UGEYwytU749HxjuZuzzjGS+TemQstdNQEtCndiQ10e/UjU3bhQRfTP1Y9AvyiM11Vz
bvC9QkJxsZHInU3XBXPCGy9HbxRoxrEbHWr2MJ6tvZVwdwFk7hOWejmRA1bUEEc/uir+MbWDJpKE
JQ8df3wmrli2MTT6G0xk1vWUpLMBm5aB/qbM7pkGiq9/P2vyKz/C64s70NJcl1wZgqRPqg3nalDW
hDQJ2KutaLbL+vejNbLTpTp6/0qOlmnKY02goNaclGIwQRQkK1T2GjQIjWXvexBmWd+9OWiyYNgh
O+RkaLAXvbwrMIYI69M1nxqKgtd6VhzXPcIQRSGGZGWkhoFQRouDjvOODYkXpZwmjnbkUmvfvXaG
gbmD2dRPG4azZfUVXyeWGQdRek7sprpnRw+geOfxAuES0vmOkiXdpZHY17xTuaJlz5UQjGaJ4y2e
qXRtTh65VPDee4wnk4LL+x4MWCk9BOAi/c/wgkXN1M//z1o5b1EmLncNrIOEnx3Mcsv7cQ1Iw1vX
Nc7t/0xhzEIhCHAnlekI/rWdI/X5hxmxBw5e+brsiatR2bv0Big0hmEsKR6GkTxKVXX8ZFL1Z7ok
F12DS+Ql42B5qwaLHXdw6lE0qSvlWm8AiXD02L83oCle3KlxhpETsMlO8CX4T586mAXjA+yPkjJI
AUUvDMTOszOE6FiN0rJVaHKS13A8diu0sc1kA1NGZcGUDDu8nlOeun0OVm7/yn5/i8cXg1UInI2m
uUJEVhvMC/o7wJ9Ba6K8ufJzyHuCZVFkgEaEusHfRmg8cWw0RFUEzBfvLJVgGm2RKXSlOvamLKwH
cWuLYdEhOj1oYd5McwS3hM9JhR7Ldpa6zRYGYmduT2v2j9m/3JLhF3z6QaS1XLZPxaQwogbwPlkn
HrhWHrAOpXU2ggHrIHuAAwCq/K6sDfFHRtpmMlWZK7pqN41R4rDD3gh3kW/jeHIYDPSZ0zWz7IRL
9PAh4LzT2U58i60vbTFx+kRRx1D2MZNLdAIQxi3JYh8OoV9UT1yatrk1oHVcA13bk2rLVdLbkI8Y
WMeDpY+SAR946pG/iQ2hlUzW9vjKN0h7Eecjy/+hEauW4edNT0YzhjdrUn5lUJdILyFLL7R3/2Rq
avEq2IxWHVhvEhttxe6AWuLJ7W+TRYrpoJzC5nYb4LMnocbY7WN6eaBTxCTsY7rJEtS2A8Mnevu1
yi/Lo+VJ3h/YZsmNyz7PDujThyH0UXRXhW0UhoAwdIDXp/fWr1YWdKEsrm7j7g16V8Y/dha6OhR2
Jccdyw159JphQCYdMG1Zs6LbNzFyB6h8dzt/uTRkfrbCHEFIpFE5IqSTKj9z13WKRxBvmB1GQeMK
BbKDPP7e+kHaiohAfP3ea29NB5Sdb1Jv8UIw5NMtBr6xhgTeCneq6+CGj3bUuwJ9hsrWyc/LAh1f
tlB0ZQdK/SCwa4NVKgj5Y3oNqaW9HENFdAGkB/GjFZ701NQozX7pKH//SdRE/nKReQPh3M9NB9q4
KE4kPD9WSH414lI3Zz/dDTvMVFJf+UT/58heeV7C9jPUDRg7fu5E05rcVwZ3rM+IDmxPDw1OY9Zc
q4reTnyBK4x8B1sq2bfsn1DXXceaLCydJ6HX9PC7mEDK+MsWALtFgwYzbp8d9qyBo73nevfKPOoZ
4HuhIJtUC8CvECnxaHHGPZeQMPeuhzICTRl72VrHbbSXHxbpORGGvE5/UP/RmBS9x0/CChW/rk6g
K/+Is/jINbJhiV0wQjvWu6g4jNGRIJgyPpJ/YwfU3I5qPaK5foUDulnkjI1l73N6xd9PQRaNHMZv
1yHopi1Pi5aQkjZ+kHjQH34kZ/L3niObzJUkIKSYIUX/pi9vQgHTZVrdJzTP9JuzzU1iY89+e5UT
zff8P1cy7n8j2aFwJzg5R550WPwZnVfDEHI56ziFGp+EIB7gbv1x0ewEJonpWA7kxNTmGIG8OWSe
ntgptrl+hQEo5OW0VhFmQSM2Ez4bhYSRTDnU3J7xgLJZKFo4nA1c4IGPJcckT0wqiuaKCUq9TSy/
D/STItLrS3gdtDhCvrX/HYqumMEBFNry9vJLKG8s3GgeeOvpX9BhEbjP0xDYTa75j5EUzlqLIdSI
7eXmRnSPznxuWIYAvW5UTSY8SeByiclbtQ/ygPPTpd7mfMfPq7YTjKv9hIk2mrYcecJrEUC8Q35T
IRaQ3Fr6A3IHgk4lIwE0aT4DZh3T1GHAyhfiGNBzue+8qjQn68uszFN66GlC2HF6qqqXFmt9mFPd
ZDm2uUrRjisMaeQY0m99w/VxvoJbYV0sMAAXk8TjRA8e8qpHGGezWqgns3hhQIq43a16AuRz8aaQ
h4PXMgo1D+5BwICpcEUye6UrN6LMXZU4SIMvB/pCtNMnj2+4Bc/8YuxV5y/wTvDR2AaEtm61Kp9N
yzSyLZQu0ORX6KPtcGNkUYvdQEj6W2rOqB/q6yj/fL0wDliRTA3nxNOHnbhxwjRIXmzGTS/IFZoz
3jlgMbMl3fwPOFr1hUMXfueUErIA6Px2AZa5qZjGJ7hYnowFZ16kZiQI5FmsPT0mE2IOWc9iqjiC
3KTXn7SThk230Qpp6OCb4sXVHZHyO+/zxxqmPu6e97POKCiRQThqXjxF+eN8h4zQ3qG6NJUpUP/+
I1FV0+F2jcmJeHmRZAu9cEilOF4kzKF5729puDBzhshOcDXNCz1ggXD6d/nndUAP3OR0YmyyOUSA
3TCBtPVBcfCgPVCSu3tOmqjfPDh2Lw0LWvEpVxfAUwE3FpVFKHzEqrjEB2TsCdnkz/R+IvnU+dzB
3mnYTK26BjoPECWi1BhobYcD/bPjy9nmUq3knvAl4MmidDbul707TMh3wT3KlNA5nsQyqx6wKNDb
lKqYVTgNUff5MHvTqqPNX3VJrEtRatL8w0MufDN/Kzi0hML5+akWsUMbGjZEF5MwvXp/dZOB7iI9
CrqUaBDkQqTBpHnyD7dNfAX2HD6HtF6Z3E8hAl9aONqkEx0NUOUiyus7mi3GDleM+IfdY8oYU1kK
2ijKAYxOUZcz5Anh4yTeyg+hz7KeRxHHzTqG6LLBhJbWag3mAqmn3bspzsv91dyPlixcvPLGyHbb
hcTI5zu84QNR6qXA53OceEM7/Z0p/7KaBVCHR9xmtnrM8wc/SJPbjf6TnId8S/IT3a9qiSpQyC/e
V3dZgar/YrwBmsT8ybPzreotC8kJdFFC6ocJ1rP/ivVbhbmk8ZWf7MoRqCwInWh2+Ot9arkZdtmc
Js+loQzBLY0OkAE1LSB338JKgfP7itFOmuw6/LMbf0oovI7zs72gBusogN9k7+0IoiwfKLWcFh9k
68kWlAr50w0mQQbB8LB0K5UJp73dcaaSnzE6vQcuwYlb2/CrsAj9uv8DnKoUScb01Mqg/UYlY1Y0
g1xa/ZKr3BQ4Qoacv6FbnD1c0FDSpKJGHgavusXfJxXTHINQ4D3nvNWTxmmk72QZ7J9rnOHbVJR1
eFlLgTgfYP3/yh2v2JFuna7KpImFWKxm+05QwG06yS8zPUFlG2Wedp78j/IK5/eQU2ff7JtYLevz
m/lPkdCRC5b8UGOPEFOLOMUhKcNhr0QewdVVBoqRGeorLN5AYARV/xOAJIQNELPwd/mkqvdPz3MG
3d88vSnWf4Wvuh1m1kssppD+CJln8f/MhAiCEd+5cXlZ4PAZv3vFxNyHgOpnZCZdYt0r9PrcYSHi
eHnB1kKQbY7AM3QxY2QDl1+anq/2TbtTXlHjiZVyjc/OolDHUFHdrWypBYOg4/6/m1BTbyw5Xhtn
VJ6ZTnESL4kcbJEd9GDNiVUBW3TSzw3ndpHyuWLyD7cdVzRrawKISfplq4LNKGraMBuoCvo6GxNi
3SLlCMXnhXm6IaufCYtmmqkqmu8Q4Zvqq8ezz+vuXBFTvFUcTCHY1pnbnTUUGXX1LO8mKUVymMrs
AFDui/Wst5IVVCmMI5KOKmKv1ODMZUjRBdon95kAfA0NfmXdxWVrpm0fpV+p8Gjf3NQHuFZbqcED
TQXMUc4tWw7z+IxAycRLKZRlvuFlwbz+XWRrzg1zFk49qavEeCq++VOHOjQDIjN1xHwahgPdel2y
i0AU56kbKUAZr8xlQyQ5888txifBp1bN0y5Wwx1yO6KDkwCcbYxxRZPuaJjqGR/G3iPW6HD16ess
u6liwYklr2mZivtrY3kZhItjCgBv9dhZPoSAQ8WUKtSnmmS8rWUHSePzhw/ebsXkXmTYwIIEsPNz
CCYSwoBItWC4cn8UfuiQtCmE7NUhA15X3LCmrSRfa1uZdpZToybGMpfTHMqo81c20GxS4wAZXGRL
DqJxUOSbXkqR698Bv94Y+KBUX5pidW1e/hE7hU1QS474IpUF/2XNiRFGbCDYtTzK2OwJa2CG2BEG
D3EajN/VAltU3/SFw5qWt7HzJo6+ApgozWWQT/CcxQq61DxEHtyq6f8V1T/eEu46c9zElQkm0YlQ
xUhjRQNYNSe9UViF7MFUDrmzNW7PV01Lc9L/CKkeXvIMmkAXtdRE1wr+YlPS09jSMJ5t8IucxWuj
+kt7Qj311zFGtXEr/xiG+hhk+mPa1W+yhM0oPsrVIQhahynucs0HvPKBqqOLvJmJ7gbbRrA82BGV
OQLWeOQ3uwyWBwFtjWrPrg9/0szX04DohxIed2UksvjwxJ2IHUDityL1B+id6Nz8ClPWxGGYptVf
2zug5Qct2gKP7HDGTpcvGnaKd+KFj70k4D+2XwnKteS8CJWouMKStQgImrtST8JMkIPZGUZEth1l
sS03+SYCQ1vCU8nJQdJ/+gwPzdUW3PV/fBg5jAxQG6wDBumg4fal4tzeumtzyUHLmvCEuYs9BOGc
F9Gy3qwO8iAnBYEZpEWd15CIqkmP8h5V2R7vZPIDtlRRy6ll7mUJeSTlslfaWxdJjxv1g1Ta0jxY
XGBHBANHTt2PBGajTK9BllKEF1quA8I03R/GRdb62630XuhSmzJ/dieMUQ5qN5FXuS5BXc+txrm0
ippLV68+KxZ9K9LqEFCeneHBcovX0jMQDP+56F+GdBg9t4cN8sRsgXdU+9uKdwwkVSELGxxo460w
Cr4g2M8IKtalXU6ngufqKP43J5NFjyzafAet4lapOz3mNake8irV8c6nOO7gi07zAQZsh+CqHDSU
C0lLHwOguqS/MY85pCbOfBmMy63XbvyNGLRmg/ae0UMZr3QmcUK6rJeM1rcAodiPOti/zGynhbBu
Ef5cXv7O6YIY2W4TuoCNhNDy8t3FFnuJp/giUNifhRkHN0g9mopSzLIwIA/2dYzPD4vudzhOeUYL
DG/6pFQp2+w/yaVxI03ZB7sFne5fIkDknrUTreF0ywY/cU8QHUsiV/br+i6N3m0YWsd+uYgP6EPd
kuru82OIJqZR5zjyLT3aGjhhawTVxPUyio3am6LowTJ3lyn+FlO1ZWkrkeRvVrzEE22GO/pNQAvL
b9Z2aycEbxUjK2FxZJBHGFBbjHYbMMGTEPKaeRuNJ3NzK3KfYSh2IzfdbPQnNmKG/qNlWZw/2i9T
WaRmbqYhVLHZDB4ghvRTGEBVuBZvKE3dL/axBx8FT+zOqoYicnZ9tWI5QdscNfpOETZiCoZ8pPWL
3nlw21NeMnQ3rno9IWwUa9SmtH4xoWi6qHkJtDYLAeO8dOTO/cI50GCIAwN7zhrBThZdQcIvm+R5
s/JLY9Y2TynpSfTfexxuVURQ3gxreqrvYx19OX11SuSP9ussw9Cdy1W0NgeB3m+U9wd3ETgq/w5L
VKr0pcYBimXYBgyRJJqypzyew4gCA+M4nBpoD5hKOrijchtlfFJu7VLkDjlRsKP6rIm9wpPduaUU
bXn5xPLdVY9WXQ3bJZtqENt4eH3TolmFYsUuFD7Em0DEyAOp3mFUZy5PeWYL1w2xGDOpyUbpKZLw
vRI9Okgg32CiykMraIu8fuMK9GZIJ1luIGV5bPezDihs25wPbFVTKTynMqrdGrteWnCBZPL6+wH5
2KQ1N6CPTvYiT/AIMPD1A6tckA8qVVvfg8r0v4xORhZAlLqw4UJZTU6VpTR0szsZCuhBoVZ9j5/B
2Bk5fY5c2GFMBIl7e1iXFq+dT6rcoyzgScM1LmAiYAL9pAn7Yish+q/g+gAF6fn+AB6iL80/uODJ
w1dC5+fbEHH8bwoXQ1ZuJhgkcbaB/yi9Ij7HM/5xYo7+Xz50l970F7uVSYbKkhqJJm7zlsYiSEi8
JmEWFv9uocrlX+ZVcnO7vrlqvUnwq8WkLxewBng5X1Xv4Yf6y0io/XO0+TMAKK7KeQ5JHQJ6CS5B
ratYXHZFnV/nNRQtJMxHfcqgKmIITJJm3JI56xkOGEuDRHL5h8vzpTEr2ydmfTQ1ozbgYOJ0yQ/Z
d3+TKQsX/mZQ96/gqYAms9u5ddokSA4rYDu0YFAYpMoTuP2NrCNAVetfGnsa4Fr/SpWQ6Dtu9x3n
sxS+TOVIZhcGRkyayvEdL/DO6rKhYus3WRCuWORFpzdBwmgmoQhIRUHC/1ki6wjCTLybSEje/kYt
36zPdAGoYOI9pnNkEqOIohjsVk1mtD/64ctnIy+lvpG1L3GURlGzBq2+Y4Ze/Z4Vr8Gzv54+QaxV
tcKgU3Q11TTNyj0zMb0qrJguMMwAeO56L+sy0a7Fzvt88rrFabtADU387SkaVk4IPRH6LCTBAUUc
3SDmGv4n8pJPlAMD2V6tUa8hV+3QNeMeyfUCoHa9TcQ4+yh5phBELRhboWgr3h7A4oRZDiH+yOP8
IHS45CnmPTz8sUARxrKLVOScKu8QU+JfI8JPU6KNEIBj9zBw8+TWS2fWpmmlwgPsY2DW33IYpTvE
66WJNZxzljllCDH0ml9rj0JPPpsq3ItcbDxXDGvOX1902R2cITpSXNx/kKPpewdhlSNqK1h2Cmce
q+UTpGEkHbv9ttVNBtt7jtnyk9hv5QXOQMohchEUiZVh55oCrXSKJeyCLlegLEQQPbf3JIX5QWw9
mEL/0CczgqWWQz8BlI5MX6t2CMPDHaa2GtjWxl7OKoJDUdxBtixKwLeZFrJaqMCsxbv2aAWeYuQa
mepnhlmzGUDQPXoBfz8yZnrWhT+qvleq70pLOj784YqFlhcyE203wMsaRCmYyQyBiRUDGH7lm9dY
7A1E9oNL/b82CKNOs6+o+fJ8kHjJSuuWTj3glTkXSdgd9Wrimhl6EMgiCKguFhW3WNI8wYPEjzhh
HAiK/2aCl4OuLeUFfkXlL5OIY/hoVLo4ga21lrBZh1sVcR/yov23ErpNBqSoWdjNcsB3E6xYqfGR
ValvtvtOipHXMecG6ifk43EfmFlWw7PnrWf4/LHxQqDqK3NrPcIulGaOPV6xaCdV3xel+EjwuWv8
r/hzO7Qo+pgkd1ZPBQsoqjQB059DjhSmR6qFGSdzHNG5SghmOH5//pyaUwC8l8hN13vOSg3lCeOx
H0DNjDS/0Q/A6KHWF58pYzGOA27pgWh0iO4U218Un2IGMn4giaEjyTl9Cil9wjfR8YWh7c9htUay
2cq3zwYCvxZF/+YLPSQ3XG9+fyLGoxmKcl9AANPmFEj8E19xoug9OCU+26T9ht2dUp4w2hywjagC
BZ2eFNseDRUu2W2OsSioNZ01wkmgWUnn+uCdap8nddCqaw2JoU7Pv2op66pFbcQ8q9qzTdRJckb4
hUeEg8yOETa2rJJ/k5p+Urfd4fpTGg7A0hkSlUWqKS/du9PfiIoKzkNNeyS6LI8YYUshkvOaGaaD
77wE2N1OC+peBKlETOoDFeZdRGJ9UMixUnyTB/T7DEZy1dtny+7ZeV+S/Qb/uiItt8OTJ4ch62ms
i8zu/HSENdkSqPrBL9n26W4OFJoMfAn1OSDveLVu4wfTG/OnimvNFVUWEnXE3kh1AKuwZgOzPyRz
mMHXVTaSa/GEGqGYFJChgqUYppJamdw1s2HY1zbUUQpcotIY7LMts++0fXs2dP/o3bwWfvS9m8I2
Eou/Usxmt09SKDs0KzyonCl4iR3sB/YzNy2OW+rVj1L8I9+w90tg3E2Vs/rMMpI9+byVD4o1hflp
NmqIqrorLHhfOANxgbdU9vijXORoO8huBqz1wfk9Qg5W8du6Pl/1elaoaK8TAQP+BH1BgP4hLst2
gzu5B3J2+LUPvVztglvFo7GwaY4ktC/21jbcuvtG7ZJHvrrlzDxs2mgLwbNEjnA1p3fOEfHCxLK9
Rrvsx76GBpo8QhLTWBX4RE6UOIFcbMMehR8RUrH04Ql/4IwBlQBubPTclXCxW/WO8kuWmuJfskBJ
oTSbAEBUkh8hDOS2h+YMd+4lvVy3Jgy+3qbbDVMRRRUX2ib6683rl/coM9Jyn+Gqw5hBcsX6W1Zo
JiQS3pBn1z6MZ4I5ycLR1Sp2UOax/MbwnPldTq96iMDC7JL8MUFwcjQs1fhEfjgCnz4XwTflsPQq
mdxabFHtscOm6pmvcsc6X9cnYZ6D7USo+2bOIZwDcKRmHz7o6NTSEzdY6lNabYQTxm8LwaI1+O7G
ntEMQf0ygjMR6jCNvE8ke+ted1odWDcPz2Ekmujdg1mAhv6nS2fzdlEqTE/iEszI1QWIcLbdTdnv
cS0AP9yfzoyV15Pd09jgsZ5Tu3QnW0jFnrtuir1RUbs/QDdnBfdIS89zhuD3nLgV3eocYgHoJJeN
UGp3Z/PwDBD5ZAv0WhP6QAaorZ52QIRALuB6uD0JZ3cR3btHG4V1Q5lJfyla54l8duI2XbcgYUxG
+L9iGRLfDNPGC5PanSGdeXZesHfxM36C9Viw/NBgTxL1q8v8r0C+G4op3CwPAnQwusjdG49I9+hb
t4dcj8+svWkfLYIrCXgL8iSaDQ/7XG0jexnXdLYePc+l0o49Q6o0B9SHmStYc/6Sm4QO0XRVW68/
YNiQsYYgxsa5uF65kKbtkMswCVx6U5LdEkZfI+cEWm3EraXzgAmtSQKylknOR9f1fkM56uM8E0sR
Wgt/k3Xj+w0BQPjn6mMHKlTMH49H9W+S3ANLHEsgRa58XnhJN9hVyWqFBig0iPySUvu/M+h1Sm6f
3xkmgnJzFhrW/Pb0OIv1xpxmpDWYof5jYIpgCPH3H1q6V2mU3GQKnWtmxzJeqc5Vv/TpW/YMczco
pnrPAQSN8gYBx/HRTBT9KK/sBt2OG7c4kxh2uyUchWjsK6O/9GuNpVCJMD2EcYdCYL6RxFcFquIQ
LZuPk0hsjLCqJAyLHvwD37EaOoUlqLvH4VwTEozoKX5IVyZA0oSGgpiZWhA567a4EQjdiceEj2qz
UNuEs8RMil0f0fUCG+w8OTRQ+kWB4OvEqRzmjd1+1vJf4+FLiyar4T0Hu5ikkBMfbvrtFeWXEpJo
D+vVjbXXX+F+Oe9eg168GUPtHlvz2SyxCGMZ26r6f5cWVhEy/CpsiKt1nQosKeeW2/GEIfEd0lZU
OdtWrl/FSfayrHuP0UBZUlbxBqjtDF46M0g82MzBGgPciPBg8jQCrcZUvYX6CIHgABpIoq969uOl
YytGmzzlUBXjtlcB8O6UNhddDrN82zuQRfw/EJc1my7sUkuBZkVE0nq6QuwJWXJijKYIvMWoMlwQ
iVGNKTgz7wzdbc9ed2o5WI2L0Khp2ed2XPl7lazdNRgd1Dxlu/SwNLNgw4sbjK9QrXifYYyHnuos
KmKG3B5c8ib8ppy2VdNsS9DWaLmTmIWHwI7RlbBEyub42+GtCryurG2UXfxAKGbcidkjZ3fQdvPw
bUtJuMnjbXyRpziUSPgTbAyxRXZ6GLV3ILSlEokdUmaBkHbZ9ecByTTZH6HyNZuloqM28hN/wZnu
PFoqlQ3YMhjgavdRc4+nVcHd1x0HA22KVdrDSOhslisJEHfyWc8PFw1UPD4BypXVx67HgaZ3bKxt
DagMTagsoa3wX47KzDPp8eYFSLRrD6ZiCvtXdZ+26KpZbH2JH4a25xaRVetW7zToZ3ehjf5cLIds
2g3quxvm1vcSLSU6z+OfDwDeyNfRnhpVX0+e11l/rQ2pUfTkvpDfdXVt0JF4M6egQGjGVutzhABG
eY5Xr4aMUCgt2/MpoZ5m7kjgvzTxgyo/eiidhX4u1aKEsdcMMeUvSn3h8pypq0sazVbM0AUIkx25
anEH368GRkVUi/LO67uevqywHx3fa9YAkU9+hvoerSWYsVlwaAoieVPbexWumDjfcY8HOtHUfWdL
j9eXQLVqJ+wFpQWnP2MIA/3EUpBH38Jyibu6ka1F1gWn/SDLNMcAOfdolpi8O9xlM5PsOThstUF4
EhWQqwvW1fmODklt7cHtl8oBzHebu1RpiyhKdojUEef55Td90eThlgnNvlMzxRI3jZNl2c8jDu0h
5+R1/IUJ5vQUqpm+XEg2MRYSMKKN6crFJVlLuy3bUgArgtgLLeFgwOyL6MCQMlgMyZsQAzbNT5Qo
aUXA/h5FZo/IRi8L5DjH03dI9sXGSDKCSlQ2fDa50Fp9HU0UxMWmYhywbHH16eBFZfjyy8AI8wo+
2wAVOMOfkNYygLBTnLHfB8ZuK73qju2a6RoUYYljjFxMYobbjtAGXj6o9uHBsZWMF9J6tO5Yfg7u
G1vtKy+c8dHGJu2VTuV9NPCx9NxEQ3u5uETLUhXML/8cBhBwFcb1vc1TVptwwtTRh98eyYtYdSyA
T7HC1DJ0udEhNgXaZEmyI911BLNhYFa3ntKWl0znoEXLaAp2grA1N0tTIlZEu8rKSXOcNG/WwJ5m
vjQQcJLlgY7kOwdeI91LGaaYiIjnGc12aY6zGzF7NdQMO2A8YfmWaJR3hunBnYGEWqNEECSkvyh7
dxHP0iF5dsWbXmM45TiD9VGTWfwRzzABPgZqM2lmX0Y82dov+3ROQvtw7IckOQguF3aSHkbX1Qbk
2WjUB3zXw4Ck3acoSspamVYxjjbeaNPqsAgjJjRTqlmkftv55cy5dLKFiUQaKsNMPxIaxSgiJg/i
J0y45DKk6f7yyb5u79y5EsKTkzZzIf5xbNYqJn4oFL64bRdYl4jwAqaxrKtYdxzKT50Y5Czcmecx
nKSMGusJGQhIyA4NPmKd+4nKui/lhgsUZIk757iyTXQsrhzv4q+xKZ+sL2fpRYToC+7gL3eInS8W
SU3WR+WtKj8AyfdinEUb6F8fQeLpTixn9GQ3aNO3BgwZoHTwERckF1aiabhJkNS0iYbKe6np+RRP
E0TgZP9P2i0rnEaeEyc3BU5QSGhTMMihe6XZwozfTkoqs4L2CNWqGu4VkbVxy0Ve1Oa20zRNVeGF
V8G0XJTcoGlN36fJ+Ygk9yLc8AhwqMFOm7R4Y2WTdrVDC/EXdMSP4EQiSQlhXWBcIuNe97Tz+g0v
Y29iqJ1kn1dMacPwwhW8xTQJhGgjMEv/cX4GhY5yhOudhApLCnP9TVpM9ecEbkW2k9uOfpDEBBGh
tQEMfDz7qDEg73nJjYjwyV7OJYUnRolrhdjZc5vIRtNTfoQ3doEsjR9V39LifVWPB2oJvviJusSD
YDL2IeFBsmZ9kZv+dHhu+BvlQwPAi7mS4qmDb2H+KP9E3kvW1lVLnXzU3Y179z8UEGJSA0lXM/Ig
WVU+lsnYTgSLsNJmXUPFmjoxf9YPVi2oqB1+edN4/+Y1wPVAkiXwnKu7Tzc/+b/QZPOC44RWpFbV
8jRwtoz3Tt9n5wnjkO13atrEh/kn6B5x8FV7exqxGqxBOZlrpiWnGhIj2CmOy0M4MqSRmtxQYPKa
2IEf55dIx8XXJy961/vQn5QzRzgAv53CPL8a8avSCrX/FFI5RiXMRxKa25K+hw3caRX7qvX1opBh
cm/xaDaAEW0gq8959KXy4oeDWcxXYZJMthK1bmgqYqInsuxCGl78ddnAN64NnY7vafWrZ9BpM6Kb
s8hsHDdv9XrDdy/mL2badNtWXgZnvlGD7T8znPMFySrqOUU2VR6sa2RDiFYM85lCY/sk+Tw9l5LN
d42O02okHVFeHPCGyQMnv+Hl4VMdVFkYedvCgadCzFpdWRh+GiTHKz8BFT056F3BDGnsX/5gXzjK
32VY1Gx0hCGKldFnRXqIgvrw3uuwsq/WlTSJ3lq2oIK5z6B5QisM/VR5xIydLz6ZNrIdYltGcs/4
T9aTNpaNt8uUmOXmbUKo2BPcfGa+s4SFG7wxrP/OUnC5K0mLKDmvT1q+3FfMyST1Gio/PcIdu+5Z
07SPze4/kFSbDpEhs28SA/F0zowPLCXYR5Y54pI1Et9DJcyXkKm9mLV8k7+CDkIUdyyRVPa9cD4P
MJefxndSgv0OIA0Yda34nEhlWTMpUv73od/qWdvJVSwVY37O+xZSNNWe9qUu45MLiGCuHPaqkyBj
majUbP8ACLWsBdYUNTyjf6idy2Knzq7h0AOkgVddoDcjbTfPGwWnakiJea9bQiu69vn/QfLLNElW
ySHbO8KPZoS3dahd1xdiSNoM/xup8gnZ+56xDgKM6gHzsHd/ccCKGrx+D1Pfz2FWa/zznTpU2dVq
KrN100PvJCWmwDpmBESxYxXPN9AM9O+1yOvIueqUCWS6EQyODFZ3nY7MLZsvgxWc8+c2ESEDy6AN
RIbDIIr9FTkXcCs982F9fdI8LiRUkIk6S+q47DXxaxPKIvKyNmdPH/VoQmPEH7GuaeJXLNR/xXky
WuGQjOtxH8b7uQPayZIfwXLXt/t5z3zQtbq4HRsYz3fv4OS0IsJ/OQMMO1DPF9F2GB+4jPCTV1YK
rafUBMXfSdX99XdbrLcb9cgUu1MurcI6jR3Gqfxw8Lbi/sRT57iusfk/+AlwNhStCVZsnfHmzTiW
UJWn+KdGPBioR9Jh6RZ6P+oX6VlZWjvuUgjRwscYUvsK/z5ZTOtrkECrxDzFF99g4cYF1D0OYvB3
Dxtdc00JDC6IUiPOi1VLFYABZz71Fp4nFChLv7sTILZChdrWhO1FhpqzPTgqtQVGpw5gqvrxw1xV
eKI4gFEuAGT5dKih57I+b7GEtQbxkjC9YwFRcoSIJdhrMEaTH2LV1w5ut72tsPiNiX0RTiOxJE/y
awp3c/9clgpGyGpXbHK5KdckrotFyaDyP0fhzOduRMo9aHxybLlj991eQe7/jF+/xc+qj1uG59UH
3pxxfNoe1JEAa9UDjJWFI+9CceQcHw1ngSPlJib9FPDpiKL8HWVocXXIHlIckv7bUyX7EbBYLgcI
M09N9h6uFliRqMCYAbS1kgHeIUC0yci8eoQKq47MhB9XFAM8W5mmK0Oz5fDY1p/zo2QO9QLlb3Zx
A8/jKLRtzxnxeC8ZikeUyXORm3Z9YOWTYPThKfdplle26TiHkFWaS+LhUcKHd2A0mZgzqdAyxDOH
iWW+gD/O58Yors1HTZQ2Fov4o/pM1j6JFNIDEvtAgJhW2VroyL5ExxTqRoBiQ83wAvmJWMyVpN70
z1vY5scHRQnbHN1J3tCk6hVTrAaJBAlj9niy4US6985RNRfh0x4oeDpAZJ5quIKlG/5qyS1PUufF
PsZXFaZaT6XLqHMX1SMbpAbH0s19mREzeUM9fJR3TVzsIQjD6S3GTigI/rhl77z2CoIpdl2qbnHR
/nwbehsKaFeMSAKxlVIwJ3b/BxWdqgnjZLNvJ8ngqztj5XW8TPu7s4G+nc8VR88fdlkeuZ6rnGRn
k74t2neOIgxfZeTktYWWnHDrykhEIo1Cc1g/IheJS2kCde/Mp3NW3x8iFZGc+sV09QGsxg1zi9Ty
rhvc4dO47uQkpwbh9is6IlaBV3Wzl9rgblDN2vrc/AhQxndrtng1OnOhxU0zSSfBo2XjhO/DZdKl
IZxHEFbskpAg8qX29W2s8HAgP8YKi3UJXff07BwloQc8XjkakytmJ8T/kTERh56FA4tldM/BvqC/
dMQtw1P5l+xqg0btT18MFPVTQ+JY3fZpsPamoCt0BjZmagmSHOarMmaWpNuwx78BQigZgf85qB7+
7jUpagmG17nuYW2Pzq6ndZR+cs11RasBcBqv2Td90gpX7orw8NmLX0Ue1pXfFtEdUQKdCbPzHpzk
o7SDgqcYuIVGUZJ0OMkfdpLjCpPwKvkVhNE5RDlGOhzZeAv6H2rlvGg2AeaR6wvlim33o9NwkOIq
cMHUnIa3q0XLDC3LtmYnUxzE7gAb/0GMIkZFGCQaPslHdCg+bz31gOLFeOeP55qru01fPOlM4fN0
ZeiqNm3uNvlBNnXq+iqYc4yWxjTbTy7awXoWSYuLCcgCGXZyd/bMgB9xNccaz+3VlbWlZcRPCiLh
dIwuzlFijxXmz1Z5OZRMM75uaVnU7l93KaomMtuBvO5sLzNfqtVHsuQRjgocU/49Uugs3gvAT4nE
mSHHEF29wyIQQKo8bSAu48+LxWw2dl/yWe7srBnd5HpMobtJMuyiysUM7jA6/V0ZN2kkUdk6due1
xD03eafXhHfU2NuUBrcZSNQYSI87jfbDHp4R2MRbcN7sI8wKTmGceUAgcPuv7tUnjmg2rzhGuadc
UnJbMjOn8A+S51MGTVcBwCKuOPSKuIA7LnwO/8FNssa1XyufBoHpWb5YrWJxKouRGcsOiFXslAXt
8ciAeTxU3n6BR7zC01zM4Y4GVTfYlSxKh7cDT7nbjt2n7WAsKYR549k6JscPBvwmlp7sT3RMMnQG
Ht6GxnQ0IONITTB+hlkVQEkVB5oKTXkVedaMQpr0p16VL607wV8igNskN3pwrzk6oh9NZMMjmYzO
Xz/+8POsLErYstS2I3Z75Dsg+6/VIyV7qVPjNeoCGnpKB2bYxUOT6pWeMJS4mNm5uTXwzDw0Et7Z
hZXcZob45kY/auMU7+x9bETr8vrwvu0x0oBUCM17X6+CfRrAcyzWUfClWPDEX2BBdFj608iA47Nf
h+8xf5Ji24tFD/vE9s27ZXJQX+X7eTi3c5kKelkCOzcsxOs934H807GQ8bWk8JpWVTVn9itRBTt9
q93ay/fi04NHKxBADk8+udr0YYgeq9E0PjDzPKy+mJGX/xDGtQm3/lAT3JwzrnE3tHSGrS3kXyUw
IU6cIeQqxdB9rjMuvFZV1Wm87FkY4JHHRTyOMD8sM2tJKrkHhclWgDlt8MKxJkHYL9IrBuE4k+lh
YXVuWXKvOrEEq20fhPeS7V7fWJF6EyyTPDlQ/+oefijybZNPauE2NkJc78350RgSvQW79sIkFL08
LZl0fXxk6qdNNLMtnicNG+Nn72nin6/xN+iDG0A1Ud4Q83JpkN+cki2jvjL0QKFSkEFypDmp4nmr
kooKKQWGU/Quk4Ta7SB0RQ52DiEOAdnAkSU+VB+X47N0HfvVxpGd3Vgd1SPSxe+dTqCR3iKl8Qe/
SinBp2c9hjjdLKrQFK20jWh18odLw0mWV0noyW2fHnUO+z1IwFaUBa717dSjt7Jk1B2X7YEH1gtd
aArAmr3hOkJmTOalz5aunn20AvcYl/u/7odqfkfIWnh9IWBrmzDx0d0kXeL69HgpUJx9DEQ9kAMT
FnXzHrjyjdOxWKgcuATo712gfbfMNXbFGjZjI0rLpylHRw2F7jo2QGheAHbrjhdSorCf9A4dy5qz
uoO+nQf/lghCzU4zAtWe4aqp+3DpGfWGthoxSv1gH7hZuUt2YKmczazzeVqcd/uzzQg/qaHB1XC9
hWZNtLPRxJTV1VN1G2mKDOwWtXSxd6Ayokvi4ZHTwkoR+ckW70vn+kpcH6ZV9VyrHrxn1HHqhBWZ
zAWuqibWXKuLA4RLjRB3Ru55FHlOPO0D9F6/5KrkLR4UFMtO0Li6ZC5m7vrojz/7MkXZ16GMYzMd
Dzn8Id+gSth04fzslPbOcrTezswGggm7ToohLbV2EI63JHQYe7uEH9oqzB6is8Pq/UGLwAMV+pV1
43mZarqqL0Z3u3nf7vNueM1uMIunrimsJHGeghlqpKGpi47aM8WCH7ynpQNYl1t2kfukNv75LfUG
fLHaLS0NI5ZPcYLvSWN2h40sKzWBfLoKD2020oPKMTuUwZgAJ+dtePLhtW/Gqu9ibmPAXKWgBaEE
Ehq/eaultntXqaN9WvAGXhTDvNeOt0wG2vxAoKA4C01/L6AlTsdL8PPtPmB07zvhN3C7MeIJpR1U
s71z3chDztw793KFyVFQDFmGT8CrO3bJwuOLxQBkUTNNhdeID/pEQfBhKMo1X+PJvnrE8vEuuVVI
Do/s8phfbHMHVQMqXY7jagkBosj4wajHzpuSqs6UdOWaJTNcX4zTTcPXR4ffEYDRGZKkv6fB7Pjn
57u4V1fX6y/4Eu7jNvukpl5/GSdYzRsZ0B7w1vuGZz0uL2ucXmTeom9jaCXBlzUKtfn4BjgzXGKY
ZwMVyEQKcIXSlhYW9Uiat+QZFLNHV27TKSDLzIShefU4P23GoaS+9qofnupycBJGqsBOfIEXC66T
hpnLi4e0BLCGgwRfmGaijp6kXPxnzEhzMEgfLBlhRxD21HrNqR0h5gCe22m4LOw6UR88qLzzpojE
3ZbmFE20kUTSVomyRwALWUoEMp5MziUs5jxU/640LNCWEsY7wyhlbebYZNN2GwojXyuC8MxBoxkg
LqAR586pp4Vfc1GxGMnlrRTu5rmIY6QTqCULzg7utSwyMM88u7Os8n3z7Erm3GMPwrcFCYE4TXoQ
ouLzwxLy05Sanfi36CYOexE++3lCEwEYebe9WsQhFjK0PYpDViwmCFw9CIBMuRBJkwLY1uQFMqaR
6DRXhyxmJUMyxfYKmYWNXHrDBHfI3a/9RI1uLEAxNU6AgPAJhKKEU1c9cY3TdNmIYv0XtG01lnAs
R+EvbXd2VuJypAGn5fK6LJbLJXjEUZwK+uPNfprbhVWM29n8jeL+sDu7RH++qjXc3nP/Rf1ydOft
d4wMmRyVjsUDdM/mEgOZKkX1cpIACtEe/onOr+cucB/rrPmwZNcZ5w46hyCw/d0fCogkJXrbrRR8
gm6yOY//Wpd04rcFNPNqKG9xkOiiuxM+QJcp2/ftjDLc0GjDiP7uSeifMvfHNMCmeu7gmgqOsOHc
dhNK8sBLjHkRde79MvKMWGPWXoumqkz+xkch5iGzaU9ujz0dyUHOa3UxLfaD1K73GNVylV3d72Bp
OGAUyxv8VTRnrc3P+iNCDYhVDXRgMNAXm1aTmt8A4tE3fzbPQAm/GLaeBNCnAGixSLOzLaLXuuCi
S/GkmGtxCtaTnJU05ngZ3vToeQRftl/Q8FNEqqib9ohf6F4D+1FBHJ8rXKE4HX+vchlrhJXUjdSN
F/mr229KS1eVrh2v1D/asKBdNGvGFYEY1tbdyv//0SpHaMY+vxn+mwIE5dHl4LdshLTBRAWhWZCA
aV1eEn+7xa2WMcE1hUMTb5V8xllGcJLQstv4FaDtIrTkwEFLGJsxrfktJ24kaZ/lShlZMPZ6/meI
jfKr3dFdOxjuI97M1evE0tVJ3Wi7jEuoAzVaHzTA2yCK6hDJTHtX4oP3Ndc2t2iHH3OLOBzI0NY3
TtwF90xW5T/CsCHEFaTLKs7TewPESyl76GL+84WgYqxANZxC05qrqJxPcHNm4TxDvbn2TMn6xEUO
x3i8Qj1+YE/YWLeMCk+hQcxjaRi7VsQoM6PyExR4aJ1W77EYWwpYX/CSUvq1U+WdNFuzXaaSYlud
Cz32YBnAstWpwvRzE9eHPzUJk0bN2gXWKXU35o/EOEKgEC4wpdeD1y47U/6xQrGC9Pe2dTEv/c/c
7GIdNsK15UXxP/fVLgnPmfSfUDWlGNmpeUPtmidDyaJlgvgNzaGwyxnurDSHSx2bCjHx2KQ1H806
UO1Oj/KYWUakLnvJ/aj6NC80jTY6Izqz3vGBIZwzQZymQqywxlC183uC0qdOQo4wDTjU22lzzQdG
NNkDQFA524U5TWIMsdGkDXv1aqK/SMVlPsij15cG++h7kOoZh00RDdO5H6RFIOIZBYwReMOmTydr
UwzqCuuU3Kg+WKD9vRyNUgKh5PDcEoQiDAxMqebl3iLygswjK8DkH8OfNZxY1U1K+ng/+MPVr71G
hVRIZgZC8WpjmPclutyMMGiX+kjL+qFQgjnLsD5fabvxszVm5yGypkE05IgQ92qVHIErgSqNLRqN
imvNPYAsPpsHKZGWEkoMnI9jC/zKF6WeBQhjx+nEN03UFYnOXJSfbv7FIpRKxOo04u54tDE4QRx0
nB26qcXEgn/g0m4p32Nf3i5a+5jlz4hRmnQGfnDk82FMaeQRZY7AUoCd38cZz13+8NBIf3lAYwIf
Wpznad8awjOQwOgI6BzKAtV8eEq9P+jXPRNBy6aJocXxuQ+w4aFoUM9JUXdPZKqP3cq/xYHnjv81
rS3cj2bnVQPwQLMOHZyjIKPg9DiwvMYSxaJ9aZH0H+Zn0LigFwcL5ecQhx/nOi6SCigEZ9dH8tZf
k42CtPNblocW9dqFcGVWX6gUQ6sSM/TY8RpGllof5rBZ/TckrAPNiUjWwJLBZ/j1jmOkVJdZR5TO
Ky+TTo10sHN9ud9BQdpnyFUGZwnYOpIraWJso3Ox7HYdXPK4a5xQT70wg9KDCdWezGfn54uUPpky
+w+OFdTY7nyk53jnUwidvORyt5vJVTRS2RRNUklc3ZLj8IEXn9kp2KckhlXt2G7ncteX+mknxuKm
M+q2rvOCBzjtL7SjJmRTtmc8V/TR0L5zWphsmvuVb63yv0CLfPO0qtC4mH27yGN0TrApIe4o8LiR
HvRGP4D3EbuBce1brzOx6hOiU6XRjBYtulL0VkRi6taNtd+9XGszphGULEFwU3EcpNx0jGtHga8c
2HY7VAO+7wP7tUfjvh4QwjDZHFI6aSZ00Y1zbhuzUXqeDV5E3ww2V9vfGCrU/xlu1pw2B5JSd0lX
nuvjRyGcrEPHr8ZQrnraXiSPG861C8qFIZkXynOjLwHdnyFR+jXUAexMu/mNWlDqiDwvEbAiyaKi
R5rswSBM3ysAR+f61Dc6xXoYApLELMV4dC0rtT9ALn9e1dcqqyW3R+CkFzAkk6uKX+e2XNUsCs1y
w7Os3j6EbjLPWzZKwnMeVUdu++YrOfYJ7pl0WzU2/9fCymNhJu3kucOyKTZfA2fBxweTGsJ7hGE9
4OiDtqp6/A+Ua11RdGrDL/g13G9eKRCpEndnFRUrDMmSMe7KXoBT14aiVSP7iJW9jLGaIrjDZpuL
ardKO7WmjpI0DFjy6UVdt0ViD2ZU4mZTMkfXLuquXgDza4jcVd88hIJEDVshnBpqtRGDOl+xfg7W
gQAMSKjbt9RPJfRqNbRJRS70wMjEG4Gx/MbMLB9TgipobLMPAeufuCOSxrrUexF+z7fde4jf4xXO
C3PvMr2mT2g/bGGWdusu7pUpvgbmJ7+7EJRMhYkPT6YVOq6p8dcTzkq010vjQFn3mUqZ7tD9nLKk
ngn2DgIIwj66giYz1bHg7C8EWmuLXP+XslSjSOgKi/SeswEwgJaGDxAPWlT8Ni0qPBu2S7BzC2qh
f8ec+yEt7PsLjNfFJDvSLFix1juCf9t0N+uALQR21sflF2PUwDyP3SsLRcLs00xhPmZlErm02Im1
J6dqg5cE4m6f3zpFjmXGzox2/2mt2liKqM4uhyVQmMQG/XTCdWNfvldRUJhRrascGGWBZSgrpRAB
ujlbGYzySj1pfxeODLJf1aMtEyk8xihAetveXlSFJACJbsjcpnUWeNqC5GNeLSktBGht0s82T0Pz
/IELgcDGj9fMVK7gHvZX37kaZMnJVixkFv+7MIGUqXti1OLLtgWSS22lgHmiUCXioJlD5vZ4dPBg
h15VsmxH1FZnySu6Wb9jkpb6E3jPYW7eHveNK3RWcaqr2efTrzTGGvl0s7vszDICJytnrlvlkD32
UqjQjzBjU+w5H/761o1HvLNmFAw6V07o9eBodCqu1zqA6SuMcwFVt3oetZ8ZxlW5SFt6NXsmA3R6
c0DeAsbP3U0LS/5lIZb7dp/TdkB3rUzOb+dX+mz+9YXI73ytEOs3ngO2bAe8sR0tmfHTmfHbYKz4
8UTXBy8KEPoqIfqxI24RZt6Y9Jp6ij+JP7SUTAj7nY2LWq1rBIJqDmrETMz7ES5wiFRyr93A0+N8
panN88dlLoXIgZGfEU/X5W4DCjVuk0/xJfTbJSLUkmBt0Iq9Xj3L2cBJV3zWGK9sg6drQM4wl+F5
z97YJOraWrNmGUPh0yBbM8/MQR9nUDpWOczd+FcCM/xqAwTjpoVbIWTyPuXtL9/hBNhXOaqUqFcw
AFhxypcNTdAUqc/pISVty47Pnv3Y5mxnQjAYo729VmYKfoNBqCDT8vm/GPP+R+liKhgTdNE/4LsU
IpkrSBFOuSgCNqUEcTL5cM6S44Yy1t1u+3fU98SveZVvIPyrCq/2YXy7n42h4TIx53NnJj+9PsVQ
8ip72Z2mgYTi2ykSxq+aPSc9U3ZE2k9+8L9sUFOpFsX7Qo01XK0bIug14HXwGC0EonlPzBOTMWz0
wEAMB02Vk65XDAStOnKJiESM7FWVV7Zasfzr9h3HUWrv7V+3BZkUwFB4Wj+RL4XK6DPoNDlqnuU4
eyDkiP9t/bBTmWHWXIdKm7ngdohBJm42uBl1r+MpcptjjVmrgdYUmsh98mN8fdhc7yDjP5wSzduo
IkI6XLMnSC/9o3LinXnFayYL89yRRvk2cBgIJwuGqzrkaPx9s7jhfMOZoDoZxrNfv8mhyiXCBJ1y
/erbSGmHfNW9ouXn3xdhfP+CjXtAoKMm41Vr1IXzG0AMN6gPq4sJTyd6Ultv5p/r8e68U0pWLvMh
wGeUIXsbVxvvfzwrAI7mFz6ZYkd8FUZ28zSy61Te96zJXcsWCt9ViieTfmB7nJbc8TIiqRHB9SFs
LXMuC4Sa89vyn7g+H7Aq6AByY5W1XDLqS94jJTktRdf1zVgZDPe9gBx1IdKBat0fBSfJUpeGMeMr
jt5PH+XET3gWtuINJappYWUOjOLutNlU9IqH7vZy/YKDig4IH2dBSdfVN002wO33U4BjwY6XTj8u
XOuF8c/Sb0nMQuAlGznf2DIljBwknw64vEFJ6f7tt0Ci05VISX/1utakVyMjZRyDp7jFNijmLqR+
LABW/7cYa7Avhmux9fZ0rQ6xxHnZRs8Q/jekmc0R1rfeE2VHAnfEcmXTkIefcpC0X0u8orusTfKQ
a5fqYUr8VIp63MRgRjtK2dNcvfBVXk5xovgYX3D9/bmCQ48+JTeSYBKnjImlC+3dnAjTFLlq8Kbt
hpsPGcalXMoftvdAYwsaqKoFSaeFAewqGiBPcmU7bTnjS0GeVZh/2lV1IeQz8iQCF/iDt9IKmkIb
nUVIJQkEsz93pRuaezCNKFdhVWfr5HKXIP8D01XIzOacBetSq4kCf9qa2XKRdhDewt3v8tzrJ48y
6KYsMOGMnq3Oh8/0zHGsUF2iYe9tZNUnGCdUAy6niwH+/XbhMUjx1ZdnKX1wRJTnZL7l+4WncH/i
kgxrQZMkMVkJDj3ZrbVxgauqzg0LR2n2DYB75BSfE5lrNFfM8mmtMic8IngY8D24GTs8a+DD7bCg
4Y50u46KkA0RDFyGEu76UcnzCC+ojS5Ylnb7EM8gAjr4KgLrPYiFvzy0+efAg1Wg2UZBB7xKaz17
q1WFR3/OFUn460Ba9HdjcNRn1BMyI596VC0e18R7xToytvZ705AXIYM3bVhQaneAkirHoWf19Kcz
CoSARckTIf/yVcqPcsCqbkxPLsup9xXE5jRuWSUdddu3x9+JEiOdCAdvaMyiKVMmQvyEP+deMU3I
+SLme1y+2j5BYe1BmEmfdqT8LGTeFCrM4Y/8+Pp5ES7zf72L3TxNNkWuUCm5YpD1caQ9l8UEsYTx
VS0OQvW3HTNSK+V8WzYE1kJ/vWJmIpn7IlAGzfMAuJhYfaa9L1XUrO/04bw/01uUydMyRiblgR7R
6uQHxOj1lepWV6e5hIzAVbWlFsA5UevTZv3K2IrPBkMNJt2MOYtI1hPshZPi/A2DjFU5vB+QEhjM
5RrKrSPFcmi07BiFzUAraTwQ10QqOf+ATI/qMSKuOg7AvjxLpczzbf+lCy2oZcvqO6BHb2GN7T3/
oBT8Ma2dYd+CZc0WOIHJafF7pbSOxBtuOfKEjFnmFEymD23Rm4lo6eZyCkqTbiuP2jbdVdq4+fBg
BmtRiuulqpq8qKJ7DFXy8PPm3aV5NCahcjfjqjUbzO4kG6d4DBcUoUSmWbCUMXmm6q0OwVgZvrgn
tJ7qmwt60d8J/Ht3r1Iu7HURIBvw4gPoGk4VrkN2CrsfSu8CMUuOjW94T4W0QNAVvLQ1O+Msg64r
Z4koD9ThYgMt0TMhPfGeVlJBxYHRDoOCnNvmLGb2kYl/3rzcTIGRWWlhEE1L2i0WpmY9BZH7DgAu
FRse+X621Vb0P+OdIiy2i7luR9oC9WB2Vpm+9Mn9v19PI0ECA8gGIXTvpRsUFjeXk2TgL+N9LKFV
JtNw/jtlyg3jk2ze/cu8oYIZgktAFc3ytUAxiM9UDdq73rcq+5/BRH8cAbS3rkX2/mAf3ud6Jran
G83dH02Ea23sNG+zArpBv7Y7qH88Fks3OSzVOC05Rzs7K6YX6fTCC8CDuEzvfuJHUFXTFjOGOOic
cpFRwJ6V4OYEaByGMx/NNP201Pvdyet82gsprRQMo6j4ICNNJwaSiLt+Vmy7df9EAFDXi4zvfj8I
cyhVKXoMhVv5PVJmmmRIrfPRQoOVGcJzjMgT51oC+iyJTcxrpCTUYnetdSW/+c+vRlZs2rbEFTYT
E81GF7t0c+X0x6zZBr7U/qExPYURk31DYvdHU6NqV15kaxra0RIs5ZVn7kN9O9bLT5VKYzG7wTOP
2dU8nlk6CYLc/AACGBPR3ha8mDuK5eq9kSFr9PkPM/oGVsNKsZT8tSzQttv7vAppuoav0B2CVa4X
PXXxK2x0RyqJLLUHpU1wqGiXiZ5X+IpB+e1m8nCGuqykghdP205wyHHU/f+H523TfrA1v7HhJ5fM
RXb+NMwNbzCFzETFTWrs4j0XEpJKTNUpxpOQLrvyUqKY/sUnZBFBsbhNkTNAdKQ936YTGz7GAIyY
r1lHbAr7G4j//TrbRBTpN37swuL/TTsm3KpApClmSrO2UqHDBwrwfGY6oZ05W8JzMWSpdxo/9yaj
s1l2CucDoRTifQSEfwCsbRnXHA0mq0+wzVGicnM57zLVMn5ERzHcu4o4M0uuzX0V+ego5O3yo7pn
rfO7mGDsworwn1ImEjcMvB3kuVTgIay3J496DFInUHpxb84xWIEI0gW2kARVTj6FkR5/wqirN1qH
6gZhcDyrkUlMPC2RYOZuSOFVyYtqA6uxi6NSejNmRNQdlr2RuteiG8x/KcXPvuiuZiLJVScFQ6Vz
P4AYQtF//oa1UASzVarqrxi/v//YdrR6siAY+bkKHcFKuM6sH4F2JjvBnpHbJAKBJEWEPZz5O2em
OABVPgA86QwQd4jXJ5gRMnuG3Wzw+YpAEz8M69RYVY/HUL/UpxOGGPaeqXdW7mf7jNzUa/Bmigkb
swbYB6IeIRvNWJnph6qeBXX0+xzBDAMdCOH9Ab0ChXJ495VXWWQuweyW1wrExs/ZfmzFOk3a/kPb
llkjIh8DbNsYHBaM4BqoNqYpGrIX3UoIKMC/jZF5Qx9hTaRJ3fEr3KCyQmIHZdtWP0ZgglIcE2eo
v/YGeWc5821Ll7v8KmQw4wmpNO/HNG+5D5k39fxWm36+b0yVGVTYS6Wn3uVACwlRicuO91DLP/iq
TywNQyzB6qzEozptHmTafCgCZAyshlTu97v2Qv6KHkVl4ZUqsuwnVeF3kWBgU5LRKJaY+QL+Bn/7
iKGoGOcTgZlXQ3VUQdYZkEUSMr2YwEPkR83ib6l0CxP5r9rYTVP3RksiRJUtrQ/Oj7zuU94SMVpH
JG1XXUV0kr8kJMPsa2BW1bHwkRzVhC8MslAwaC09AoBq2pdlxf+neXzfyiQxaMbGO19OPN653t/R
B6tEKtdlBZpcDc4F+pmGVicmPlT8I+ugRwDfmwrcJc6ylWx5DfWd6ycEOqLdiqfZ9KxQ4mNOn943
2Yy+WcFV7h5kX8Kg5mkOUmDGIhcAeJ0H1wf0ChXBO5CI6ZgRLq9gl0fstiOPmOPMCp4PgEcSSgPs
U9wqM02tJ+RHDPvcTr2pI4JfR5mq6R6q2UkGB4qjg4Mjg/L8ajUuXqZV9x49dNoD+F/xOJhJmvMm
J49Sz2zw+zAgoi5nZUUNGG5nPRnQLPnd+2pTgsBPPYF3VdY4aXa7qatRso/k00JW679nW9VJOSHy
NsFyHreNVPU64asGmOrcscP6L5PI2Gx0x4QDAZwx/d/k7qoywmKzpR9Fcs31jZRX/CGswRlJ5koM
a5hbQGd9onlVwL0l7O1HtPiFR0/oWOEfNSiSDTGiYoMNL+9JdMLIISx+v9aKiWLXF+OxiFz0b9B5
ieDm+qPhJG2AEIhpbrA9x8oROesMLg0LR5ChJl7J0PyJpP4XxcpcSrQTlpU6dk0R2dB2DJQA1hIo
T5YGc9AGHs7hE1sVhhn/MbksYqPOzF58jOVnHqJoy39HMNRc8GCfumdbR+S7rCVSmakvaTqrHv0f
kxOXKazimAbjwMgeuWm6hTr4IjfZgH/iI0shCTZo64yq/Ks5I6a2ecuu48W4itDsnAesMsEAc3oL
jg0ThCfSiSGjKlDrMnXeM9jeeWu8LC3X6ect1BGJGrFt/ysGqHAqcozO+dyGNl6oR/CArGEYGIuu
ZI1pP0ugPK4wdgAChdFRVVwPj1a4cHf/1bTyD2pJzpNKcfL0CAesEZIaIr1bJJ1exd0XqEs4pZ3O
aZ2lBh74Zeb55VkirgqPMfA7ijCy/kti3z8XW/N7P+ICHhOrJl5Xdcjc7fRRYsD3/jY0DdfY0dhW
Ye0UBh4R28KZpq156FaAVqIY5XD72lNMCMnAUOQs2Se6+HgBxhCsZH+Jpyg0OTPOdSmnq2NvJUMg
N11DmDzulz5B+5RCgsC+rAL2rvLmyU8Ff1AMOSJn7lSbjjUrhr/MEvnwVm9F2s5fVVqYzLgx1EWL
1lMdFuitqhm7O0oqTZw10hsJuZ8iCGTrtC3cAr2HCsfr1+rtwebPlTLb2OlZTSH4hVaqRwcnZzUO
k6XIOlvZi7c4SP5qDDJF8GblYAvKH49+shA5UzRyxN2Sch3HDucm//CHqDL8N7bUNw+Wb9sfeJR7
jBMs+TgSt0XE/YPua1rWPQzJtzf3LwC9ZSc0eLfS9Gp9zfdLEnWWrt/TvAgnrPLBwN+Kt7XGUZGq
SnI19qaUa12YyvLSSHHi1F33JGZMeRzqBnZPN14Rk1eYHmI1VmOsbR1ocadYACi6DhEFATcjeAQ2
JGVkhmGMwo452QVk9UU18ifztMtyExnGvzkKbtYAuwr+fhWWA3GICi0kSP1aqPIV/kBdTW1OvdwI
P34tGfujdM1xIBYLIL5PxhpNfJllOX7P3WNiToJ++hlWGbYJHfdYKfgDuGxy5IKs1FDiBS2opm4E
Toyb20R+09S8asQ/gDPApazxNzfjn+PPp3bRvLOwPnrZn+AOdfYxUTEAJIfuys5XBEVYGnu/e0hy
0AnMmTaPLF+VOVeg0HHqu/B5rT8gS+VIPV98Cd8qOf2hfdh2ALe/Zo9+93ny15Tym0RkBgr+NCQO
ebFV+krZEbITZWFg+J87+dPUp5bEpbwX5FVk1w/B3ORsU3qHeeQ6Sig5n1TNf7CRKLQHycCOwrrZ
kMmUeg8MQ/OtIiJbDehrT+qkA6MOpPJcYiJuBVa6I95fmpgjuf6ZcGoMW0/OI6pEHA2xqKBvBm8B
syNwSBK61oy+HOoM4bTZm8I0pZwMc0CxLWU/SxOI9kPi+nHwDnAa6ywkW44Ct+ytgBnXFtje5NdR
KnPiR8nk/649S1iBM1GMP1JJ/WiA6uWNS0nSDQ3ddM8rYNpm6xS60M7lLAUSWBkhfhloUDpt+U7+
vE/yMGtSJXOKI7JWzWO1rHlGDEMj5l0DNCkhZMiDnqpWPz0Es2h+ctzAYSq6NuSEwZDqF64UyO53
uz+0wy/zIqEPdYTVNFhwgBZcA1kO6tNwQwwYyuX/09zanf6wqy40P4cz0d96xJ5xBVEGG7vLoEXs
1e9pWUSLAT0QicmgoG4125m+0eZVkJRm5R7Z+Di7aUKkaHgus6PBqNspQxLdE/XA09IwD04rmgHQ
m0HWxSGPX3kcyGMTQfR9bP1xQ2D5mPxxgu0Vpb9E6oZ0Qw8eyNzATOKvK5+47UxjMIrDKdsAeBpA
q7n2FILjtHkf7QnV3vysjzqsmPyD7t9ciDTBt71S0zC3wFSuemG2yacXqB83DCqn3woDHrKdHZKt
upBv3L0oGP4AC1m5JEAXqOlCJWRm7VHpzEUDU42TFgBiHRQM7hYrjHmsBtNu77KQzGrSDqZleosn
Pd4nDsaDAP0f8GfYm9YlGSA51gGjCRYy3/UUjj/RBB4yGJdqM+HcTK8gu2TBwZyREDJGBRZwI7HG
6mIFzBqWj9zg+DAIGXbzN/9S7nkmt4mHMmZSecl61PJRhjREpXlgyLJKtCrie+7Aqa22jpas0444
T1YeOYdEFvaUQcozlnjEicWjq29Buwwont1nirwyGCcPBM+2fEK45EdznWgWzAdFRgaEAM8MpX5J
cbqso6cdg0EGJdWUfEj5qNOjFj9y/+U4Q5009hhSSGjkDvhJIMIuFkHD6dF95fGjsK++StGhETlD
NwxZthuq6/u3tRqHkirkgkolx3xbJdNBVvvInn+GhETZAdoWkkvn4XAjgkAs11fIztcBacdWG88E
Ua2Kz/2v8TbgMcj3UcVXA3YcpXwOuPmpNHvaelIZhwyfNle7eJgXAfPt1RbaoYfMmKykCRS4wZ27
HTYMki99UG3CJ0xsTUBsAfUX3QdwNEikv1M6X3+OhOFHBWvEtqqZoKFaIFoWDRRPHA7EamXiP0tP
JhMuekr4o9X6Zbzo1dhQDJcBX13+qawLqaWmnVHJE0daSa6O5CYFj/iJyY5qA7LAziEolZ/+xPTF
xcXzSFWwvGxh+6oe0/dT5tsMcodk9pPEMCk1CjYd0AoNZOkkrVnzrrWDOgBHiLbT/dGVgoBYKAuO
ZWXIQqEZMFj6DKhF5w8meDnOH0I9k6KVWPoDIKqkWnUjH5UV+HWsu/LgBqyzeFo45fWuVmqaEG35
26AlyGsVjD0cPg3PuziSMP6Zt1cfAOgH6IjeodssAJuoYsr87+9MpliPICNHtWWlw6KInA62wna2
4zp2UBO+vjzIgTPqv4jLyD4OgORAv/6t/gWa55D7Es94wZrki4uqbT76eqT2WX+ADSb0GBOPvVTC
hA74cvHu3XiMF/pyuP5s3wUhOX/IkClCrY1d2YwXhpaJWes8OUSsL2HI5scP49Xy0kdZSK+XARh7
ZSfrQ7RWV6+xDV6Zpp05BRMqK5HH9YUnq5stxFvmOZqjOjJUm+burfn6qkYBzRUlIe1KB7JcpF2K
zGo6mEBVupnTsqG9cclgKIXGZkJxizFpIsojES6xeBSA5/cHbcNedKQQE/J1Qi1eCDV0WwvfVOW0
nZm4eNKHGvROCR+sCp4L6dtB5B2LjF+SmwsZ98eTWRejxHg4YGRYbCbIh1/Ef+orQbVXo5HnQ2DS
QmnBTDKEjQBXMOPJyhy9abQep+5x2jslq/eiWQKKbulbusDGbEHdiEi8evaTvBjDTxhy3xUo4HAy
pOI4isSjbgLydqTeso3KhprgyqN80kW5D0/xtCsPQKAkvlkWzsuqRnJAosVicR0kABp1IzF5LOWe
liy45F1wxZTlCeuygzVT2joWCBrO3n83tz+AG+t4nqnMxu/RUgsOGIVcOKhaC3JlEAZL+s6uAJHy
66UClZGzCECX8YlXCraTv4odtUpLPaOqQe6xy6s0T4jfQNHjmyp6PB+a9rTz4TR1345TqBHOTMFJ
L0qBuncdWGe0ZUxig/jWEt220LXHj5s/EngYKEII5YEQxf9sL2AkjJurcjuEKG9iHhIlesPNGN4v
T37N5p3sM8Gpe+IJZxPbKfxZSiLs+qRVRUALQpqjqcySwRn3v5YbOneywF1/M5cpGeXaf6RaVLet
Khumkwr8mXkOFTpwCnGDnxLbgpTEz/kmS+cW106gP2EOganBFnxx0z75GQAu5ijzIkmcWz1Sttj5
ZdjH3IE9QfXKoamxrfhrz6DdfcBr/5tkPzv8y7bN//E1ZYzmFPNJ4UNZ9lS0QWG57CLYRjl9zIhn
65HHwhX4MoLrl1bOt6aAia6cCMjHoMZIwMZv08g4Pkeyx2zQI045+tzj2flFzNfLNnjqhn4GmR38
e4wbx10z+/cUzNISNIR3kvFFwbicHs7/b+VhRN/jvmU8nmpEuqDZHj60PhboSrjezmAMpeHPLUMX
37dFWPl4mda4lY7XmrCeY77YN7GPUUWvzwDbGdH5pAfj7WrwvSGTfwErWrnFBa1joX6csEGNBpBs
tjPXiPJ8J1PjMCTZ2PXrE8rKCpAjijadBuTriO8X381mvmwDT1Tg38aQ6DhX5Ic0p2YEZ8tprniU
hXx/pGtu6xWn4stC87ssZESTZHx8Iq2316h3/3aoan+OTpqTnlXylzNnpU9vnEXgccNrG7FlxRqP
nY/61hwegSQ3ThtIu5ivT3fMFkFLmq3qQCC9S8VeQnjx9ip3BJC81IhK6UPgjFGYIGtwUN8bKCaw
/Fx2k/8Yjq1lTfmcerkq29lsHqeHY1j1uf39/TvTRELiun7IEHVS6ihY1ekUzBqxNMlB1zDiDyCc
HJvHy30+5hMDGNAHnTPhAaUQRDL58+epHRFe8W3UT5jdOpWqqdYbATP6mE0jj3URoEPWoQNmJrJv
/8325o3mOMGBuV7/qCe8sMhtcFw5Qr193DVNjIvUI5oEExiggTy8U1wc+RJf/QYtzytdFyPgCIxA
6ITwwRizsP6UelccMD+f2CDPoUCkrpNKNgcQkzDNI+Ul0fK4b1YjM/UOA+Sf5gFIxO8aHafScbCz
6ED3jH34BfxON0kaLiezcBnag99fnqSnxESd8g8VEySt7nDWMvnpoLMniAw846dmv+F9O6SMyHnQ
AZmBlO6qZWUPFAzJimNn0NIsc3+cZjNGIKU/fBXKxz45K4X6guYZ41y3kM93lsnYFmlk5XUYF3US
b5gU2sG8Oj23q5hIXOp+06QpPXE1kCIpFRyC25WBuHnw/AAqdcJX367VV1P+s3XYJ1Ss4STq3Bhl
ev1rfDBne6Jr2gafkhbgDBlFD/p0cVF7fYyZqY8kMSvSId0E4nVAnmUGRDFUfKnN63shCQEmRZKa
w8jlmh3UIPRH8sk4cQ5SYBwCeCd/Uz1MCFMW4tbaKydM8i1VT5HzpA1naDRLcEiDw8yNALnzvOzC
03nojyighAqeVtWuosa+AQkdvPBqoI/ijod6vHWU2tojhYkwhGyU7VDhUzTLLjni38BVGscTdz44
JhUwHO2hchUGu0brdME2j3sJu9LH2TF44S42JLFlklmvdhErBQqqHCAtvPsgr4s40J/7sX2Wayg5
MA/VlgLcMydur1lazfSLGBI0LhodPweHCSW5ISYMfF2ctazcdscXilKSbnL0JnKTjknepTM617/b
3TjmanJAJhnIDI2ENZLdVGl0dT40OdQCbhQzg0PrtmV+IC1hlQcGYpmss9d1HWjHyKZXvLyw5aLV
tpFMzjc+1z6eiPF821gQMvIQlYol2gKL6uVufiMuVLB7i5oplsghqchjPrlKZ9C7VgOXY1UEfiYj
bi41+lfl90Qot1leVWtfl2YBKiKxgqZmIJRcBlEtDJU0llSNRWh7bEk+F1FGTYJ2ky8UDZCszkqC
EXkuZACQc82r/oYwtetIwz3HRD19Qdfrx0WJXSfT41dmLrNKvPJHxe5GOrH8r70lxSOePdQUTEZA
X7XuvAyPzB7BzFSey6P9yXZVveYAgE2hEazRjODullrsUNTDKhcXJ1UybsQqOU7lDOlzeqryJogf
lxtrVdEE25nbF5GqIPcONE56aEeIOQ+xhDdH1gMZPfdqDEmDuw8ioHGPxZk2Qqwrogidn6K1XlG9
EGsIGhiV44sGgT5jAn2xRFCmfBA8dj2FdTuHpiONbjymg1tyd/qKVsQLr7ZYF41jhzN3UPxki2Rh
bcAfCBmep7srToxgi3mcWHkv+Ec41hYphxYcaWy4aZBrQT6SNjX53iOIvy+ub6+iOxwi114anoS+
pAYXU5mFoIRe704VZvgNMi+6GZau6MgJYmKSg1r3TF4gE6eMvo2hyin9o/bJYNacOO0O5J2GHYl5
mna5y9mIB46gA8LnGdj+hykVAU0BYJN21JzchIOvRpWVEsCHQP3jMroVGHAKgzhltroxINvNvbBI
Zc5rxy3DSzkXCPxmy+wqHNR7wHK8NQUjHtC+B/HX0VFTzBZxB7KaImeyg9v6UUi4/NEY6h1GdX5W
Vc6lO6oQa0UG6DCeL8a7b0W7sVdd7cHyAKE72Sk+pzFCfvunY/9XJzBEykUvb3E3Z89GYs5qFSZ/
yeihBY5mzu3BlKsr4/M9MCikuPKjcAc6ablVFQczUqW+mqLLza+pxQXiWlegf1qq8SBitgJU3D6F
c18eeuWseSkTi8Hz6BnZQg3idnG7dg1vqO02KaftvROZ8cemNTLuV3tbI6D2jl3R8MNJObhiZ87Z
2Pde8SQFWQvv+lxQdU0ULzhXGgZd6S2lGo/OEDDQ9qQd3z2RvuNnuM7X/ICIZPU057QDaInINGrD
e0OpbYRO4sBc/O0foLxEqLGMBI6lW3viT3aySWKLv1VDpapZ6cCkj0voebsOcai+P/ICM8nt91Lo
Hw3H5yYWh2KnlmVG6vcA8nc7YqZbuHQYiH0+BYtnZkipHdzrRB/Y9cUuvusKih83SA3O8yJVKEBT
nRywRbGDslkpUlz2KUcj1gcDp9HbK8dSOpgT9EdgepJiWn4Gtgfk4b002mIZD5Fs6VAQCvXpKBJa
giCkMmZnJ8AXX6Y7Bt+XJbSurjHeXaj9TtNgtptDfQNbs0Tztadwz7sSJBbYp4Y7Xr2fBAgUSBjs
DnX4CNA7saAQKgKkm67h4eOA+I4cL2a9n1htBP0ZXNiS7bph2XHAUGmoq8G1+oUKX3okgfv0YUEn
TXxHhGS7HTbn8JNmpyWxLweEdKhH4c8DebeJ4RmchbYbebUyGH8YZyRMtqggXn6dxpdPL91RK+qs
M21IPu4BVriPnOczbiv9wSOZM4+lNiEIJpvXe8iFXuWsEWBV0V54wIiXpTYD8uxO7rmPIq6HpDjv
ShbllC6y4sX2YXqaTzcmdXSjAF/LkLTPloXv3IJAVFwAcZ3+R2keq+7xcbt/pgLD8glAi7NoP9Vq
TY2PhJOr9oooBrtZsCKBpdKqSY2/zYvWK9JA5lacUt24adrN+Pepqk8eSBe800S0/Aat7VjbeMd4
GMugPnvMeITUjpQJhoP9mREwhdTMAtzcA6pgpuFhcgzZ9FdEofcmxiaRPRV6xNondwoWwzQhm5Tt
ccwCpMaUZK8T9dElLpOv9ANeXGpYvExIcQ7h7m3n7gUp9HzvGs2Pcq5AmnFUWOxAVyvmhNhckL7e
V48VHuikSWru+ys/ngdoZbroq2+eJFZrWkyWtKtA+ipaOIJviM8iM4I8b7DurrLS58DRKxvaVEWM
YDOJWySXRvO34E7cJzL3A/9pK56XWfWvf+bsdaKBfc+0/1WnDtK2BSIhuCAO245C8D1U/yfTmyMn
mxrOU+us1pfA3T0rTSO3Urbw4nUvu+n3wNMgl25sG7IX1bd7L6oCzDAalcUkfCMQBtzNQUxgHDuB
jbrROmqcyYeHCtxx3ol4ZpepuBdKQCzcLBt3h6MgUHBrvM+fL7oeP3nRNMM5n9Muy9UfHa9oaBLZ
Q6OJaXJaoSae2Sjcdn0j0VRT1OtKuDL6QVy70cMZxSpX9i9bbIMf40DzleXweGIWpsn5tO2vq0vK
/u5kvBaBh5EYzhFpKS/Au+gX/6wxQExbTLbvDf/CqutNPOS0eLNScqb+QN3P0/315XxjIuhLQLmh
vAhSLb93eAbYr7PudMTqcjVGZUrt9qgYBQl0Sqzx+do3rYCvgld6bWKslpiZoQ3H9jahKypPM3aa
GcsZCWkuXeoLiMxe2xV6ARYSQabBB/BTAbQ8v71iGGiRMox6MByI85IxCqSZ6fEH1qAfqyK+5/vy
tIYR81uvSWDtnMlODxOP5zZWuGc8Y6q/56bO6OWJvszLxzbJRvPbXGGTQlWymdpRxcPBUUOrxL5f
FPilt/isvCw+AGsACL9cdvd9PsN/UJ1DA/IkySgurLOBYXjWA3bInJa8X6Jpc1k3BpFZCjKoyPwo
/HA+3y8NJAgUzL9vq1nRLF9xj1P5uU7BDrS8LFrvgxkDx50lvXgEsj8VImYcoOEP/kPGb/EyPmgx
o181QKDkxPuRUpnB9Pe+K/vHmYK2FM+LA6LcVYFNYs/FDiqZVAA14HJ0fCKZAgkhK/jm5wZ5KzXA
OYeMXhhgCiRcxNB497FxbedNMKhmG+xI8fjhj55SZBciXbmdt+U9uk8b2/pr8JvbQPtNWjbgy5KJ
xh5LBZ5CWIHJJCX4dnoFUS0xzUBrvYn3lUE+U3lzE5IE/sN0Ds0Dy0UHUzmcMxhUtw648l2Bv+Wp
dbBtm4qMS8u4qN3CSX+iwEedPXCbUa88utQXWuPenc3XVySQHcHq8eJylYRleeUOIrdD/jufwtwI
geGDBaGkchVEkql/4ae+Z/lAcjbah9vbZGHjL/ux/X8wB3wnQvTYzf/JGD5+SGG6SiO2IQrjeTXU
iOVWhCLTcb9E8Z9wVT1QE9fYmIb5KeJvAHcTYFAA2y/FywuEk4tRwBwu3QgF5nf56fjmtjJGJ/YW
p/ZUwanUzN29p9lFFDukcYlI2jpd+lAusMHGMngSb1cbL80xzmkwgWDiKiWITE9CN1ZhoLDfHDZt
59Gqe8YCjytXajtUlejbK8LitYRAXzXgZuf7yRodIW0Y7JgZwa+NBILLyh9rDziQK653aiew+G2P
03CPKR/lZhto/8ntTbXfwyPXfM3U6FRItM37XdOOUAgfvH+b9ycfQi4nOvN+QzOhcxr2wUolWlqr
l43hJwCGWuXsAxWuXGn3AtZegF5GvBeaMCJPzuvnlP69iIzNzriLCgid00FAG58BSCa7PI10Oy5q
PFvYsYfKMVR5m17zza0Zc9hJzNHigJh7RDK09SCoO6/0C0I8U07lZLhPNyBGDoyD1GndseIQrPqP
m8T85lIrOSZWTuW1vOciO6ZcYnghOapFuLPQCBm1GPgJXTLeLRPoMhmrmxugw4bHKZwgCGgY8X+6
4CNLzMIfvoN31BoGXXsZTFF5o23cmK7BAsemi0b0V0/JXTVa6SyxYL+DviZ7xGcpkjyVhHS5YulN
E8nyQmpp0B12w3mlMHaaXmpnO/M/cxXu50aXZMp8/wDM39jNhkyyM/2zJnaVVvacUnFAwxNd+TDS
phWtLPIfOpfXl0cOYTaAAHIvROc6V/ecN87c1okPCYsH4860CHBTyrQvOIiKZ6Bz01hIlfVWpgFt
fKlGF1Jx3PODa92przya5zLL3UxJh3/gSLDA9cnEBBKvck0mWRNlpziYh7idRn6GCKtVwrg/4sK5
iyS6ujm83hFp+3BBHZV6oMLOC5Vyjs2tKHB6efP72wwnP2LYz9HKY+5D94Naroil//Kd6p0J2Nyn
rdbqfbOUMMhcaFry0SbuH6tKYoJ4kFNETsYzYiX+QsyD2jO85Xoi5GtcdgvNqO9WfV/EgVi+mBBC
WdU2xZ2YoRzq8F+YmOOcQmHadDYaN+Q6eB3NU75/KKuG3ed/gRLf1tOY7rw7nCXhugPKRUgQz7S/
tNa7ud1OKpUEBbOAV3i6wwpsn6teJBzr3QTe/BzqJPs5fDF+QetnN5Yq2+Odf7zvluI9yq6mZWfK
SonrFhgAlcsgY9GiQjUFxWzNbqkIJc+ed2VbJlKddTe+WBDsh/NzoAs8Yg9uuTzXs7uDakPDrIHE
5xUOeH6V6wEnsFjsqYt6cF8Ft/4cPiGIi6ZLQ5vxYfOoqjEs3tPAiWftjCG7EUSbj0Q4WBGlhDbu
4xabf7tHLrWj36Lk1UwUjbtr2e+d/ujC73iz6T/tYIOefXbMIQ/8wHLJ7thja87QXAnJ9Aa61Q2K
6GpN78vDQRXYf5S2TBoI9hbvoHFo0HaxUHADGzJYj43qxkbr3soccKMata+huPokpYmR2CsroWIQ
DBwP4AX3o39SupRzo/KVjfnHb6KKRICuvZR6mZMaDRQRi1OMXdQtuZ8SOkWBra2D9K2J7tXZGErf
NSMRAD+dxG9VUHEj6R5mXy37wmbQ2IjmeaL6pVchByoOL/uola/+rkNg82Yv+kOQMeHErpKlqGBn
+fNWoecIb8UoFrB+LjXgL2OSjvRPgrzItqOQOIFUAKzNd71LigmCt2xWc1GmsAOwU2oLZ2p/xwWI
l3SWLT0+eJNxcrllvhQTHEEYProOhLoQTJEg9ud03+0gDIDUT8Y3ZD0ySazx4RVyUC/MzDXNfiZV
BUb0WekeJgVhyuQPnLtgJGWUZ2dUyT6VY+b52ogenzGn4aZsv4khfyJ19XKN6rZceHcLrALLHtJM
R19fmBIEHgZL110lqx7PdZgl9jW6EvE2bm0UqdBsjtmXbHeUdR3qwpi9w4YsgrvnNcwosqQ0F5G0
oLwQFh1lPPzcY06tvbh61BJSDxWudNuYaDX20yY7KLzEZ6WPyCgidMIc9tw3ZdWVUmQi7eKhYkP6
R2aCTvyFY+hbYW0zEh0bsmvONxWSzbVoOReT+rlyC5Qn/luIg+z1lHXc4Q1h/zdoIFYZ7DkkpMpJ
vvQclCZRbOT7rf9V8/JsLW2LwYTt+rsB1u/5WabDDBp0PzEvSAPyUC4+I8UyDZuOVjuzdzr55F+O
oY9QUEt2YDoNHz8iWjwkQk0nM26Uxj7QpWzvEIWo+luXu7tcTc5oApUfrxLKBS7/mYyk1CjFiLQ+
T3G4pNeYT8gL3spN4/EHERL4DdlY4O/KqaEVv6vcaDFy0HgLTFnZg7f8K1PrxNRCpUcCNM6GZRBb
es30JD4rfkeBesG8FWqUt26tStm3FpWlEprGGPy2ddKSk3BQE5Q7AsotpNRT8nFHZhjbBeTAb87M
tclAiwDptoeQHo1B85yUGvpJA4aAxuOlVg7tjCpDHTg8RDFUcW+lkF1KpLquYTA2DboQiL8QePXm
8N0niFj2c8BMz9aSmbxqLRYWD1F3+fzgOvaadEnlB/gzX8z3ZqvPBGNMsYJ7uZm0jrv4dIJMOxCZ
N9MKuxGaI47bgYn1AeXs8FsIpEwVT8GyKBu0OpQpozUh+1VPrMGNRnOzHhhaA9OTDWDpMD6CfsLb
ryzxv1IeF4uoSbeVsu4yMvQGXKfkIl3e3jjvDVHw+umINx2GAydF7riqxHFq3dlYfg5DxSsxdzfN
Snemxf+OMPyzuhxA/39vJBwUN4pzXGblxaCvjirvZQnXC/Bpq7UFnYpP1DvNObxe8MRaXI808TYC
8nCeahH6yeI5Dn3D6Ne2hsuhkVHjy1yuvfcSVbiP5eTCSebHwrnNGq5HfsK2u9K0opReqp+FU/XQ
QapbVezdfk2xxtD8sXOdCPLPox47PMQaEmWt6kAWILD67VqckvDDZVF4TGMG2/sFrq6Fo5wcU0gZ
l8tHPGRauLuNUyPuyZexh4Loife6n0FIKj7CJebmrI0mX4YNzScjQbLyO9e6wBALdGCoNW1WN0ki
8wmhaypFUnYpP94UN9iMLogR/EvqbFZhanUm8Pstr+n5SgOd7gOM+rqW7AoSm7AXP8771T+FARHs
xDvPigvVBXkszoghIH2up7hDwI3j7jrPHhWIwlY0RTk+8Se/DEvyT/X+Yr6Mepr8Xn4jJTZURD0A
pjFT1xKSzlC5CGr67mLJLZ3mQnAnM/EYHmfhXEsmcAWPdknj80kppBeMIWzbSRXgwC9m0Y4mRjb7
s7OpAHO1/MMKI+RckXcPsPRIuWrZ5KJ174hp4flTjpNw1XH73rgRy7PRRe6Z1TmTqlOH44yrm3I0
GX0QLJ/krLo+EuA1J5ccWHZhqQ3QNqaecVEmCYYcGIhbVmNWh8ofXN4HHu04Vb32IHA63K4NUsiX
MrK7NpMMQqhsoO+2rqY7HTlgyRN+f9mmCyZBMF0w6lKOUf0GsCkmO9eGRpghD8wLs1Ok+94qnq3A
Hy/3MTjl9eSSb+ohc0pEPl+ioCBak0as/A+hlRdv+1XxaZvZT2VDQUwDjFeuttlQ5BS16Nv1s9zj
+s1QlXJ5W8cq2UzaukWr+y/PupRwE6LDvRVYM7NZbI1P347iJrkVc2G9DDClJUa25qFYqtbvSJVZ
QuJATT5czz+2qWp4slkNndOiNfjFEdlgLj1j6Z5Qp6qypIqgwAWLTSXbYHxex/n8Ky6EnBvUuics
dQg4fVN7/ahj5GSf+GQDd/Mr6+UReLqxtXe6CwTydXRO9GAFbGPkNbkIs2/qTiYHt3RH1V9GU1K/
9OrNj+ZcnYF3vbt1gTdsXC4zYb/laiA8JhVkuXdNuAD+/9q/7tRKWs9+fYjjND3CLK/jIwD0LqBG
zvZTRDec7OUyXY2HwTE+fTVOsYu074fNdhRrVI3AEXRk5hc2d65sPHH6fM1SSKnzFAUL8UNgPGmx
f7iBUpajLJjw0/VwEuWiJFoHGjtXNj3y6HNoJ//qr8QHzhDrCA1hl/7aeUG0dSj2q60s61cUmpA0
qamIESSq1f/nG60OW/GuZIPSh1aVILqyGxBlKIWyKFu3akPoXFxO5qQqt5m9tGZ1/PfJErRY/Dxd
wNAWHXs/Ia1ePwdvf4XTJUf+r3fbOTCQzv6UTLEmrPwhTZzFr8B7BFqC0g61k4GEwdNIW3+Wkq1/
JUULh4npv4oFAAbsEgyEmgrd8YaR3KAonjA3ro9s80+CREgRygq2CSrus005caMd5VqP2s+ydwcw
OYMJ4iSiv/sSD/I0KYoMUXCrW7gv7SS73M58Hoz/okStRDHvN4GR2MWl9Y8OmdkaExVhleIwDlkr
NgluJG97yafkHVPVhc8jyI2YZX+2X4J4QM1P/39B6i4X37Lj9PAgbAr3quRD0pwx1FTNNaG0Vlt3
MJIcJe1dJLsJKjqoQR02woQnwtcGNERrtFxxBqGXNOTYQUuZFOLdNPz4Z9NgXG1Ot0CVVc0KYjAv
ZORVMzUoZw37XbpTyBFxoNQ+N8HBQMREu2JLUl3BR+Bt8gqwe0nZzdAHryWNMQCeCXiMg6FG/5nS
WlqcePhu3FeatRfBayOr2wSqDPKTcrk7K9CSUPLMEReS2r1NMsoKD6JfYX7++bBkBZpYsdMbt382
A1iTkGE/X+ekN5ZS0it5qcyAs9j7HUgoyVHYZffZjMqLWne8lFEGGJ94BE2+h1xKtZG+QFapB61O
FPvKH7KEsUMOmQgpC1pagWkg5xqW7MnXVHFiE65Vk8kLfspwfDagn17JRdw8/N5RmH+PVtQ9x9KU
2cH+Ebuu+FWSaObccDCvxTHQrZESgjen5WS9OaVuGliiY1aH/fNmPKN7CZpkGjYEoXgQUSC8VPNI
0ZBe4M5TiEkjMgdGkIJuLFMXJnGJoHpTRGegTsVi7dE0Uj3OdTDGRthlsBVf8tNnsGUwTWL83gYN
XV8tfd38EMJHA+apvUwYhi1VHjj4SqcF0TASH0T7BMyDS6q0O5zeaODJLXC4mKrC4x51ccOysUZS
6iQx+yEqGzK7rzuufPWkvGqbbG0H3SyiuGTu4BgVWUoiOiKztna34gbOjvliFDWGFVHTQuDZom8h
a3DCcQBromAMrFUSJsIlxifcgh76dUbjgnx6xgfdumz7J4lVK+LoQTbk8E757JQy+6e8QxuFnkjt
deQ456RoGYK6wg8DaIkQmqNiLG5qsowvo1lqRRV9lgwyLO/r0/yyR48qEbHbZnJMXnrAjhr6h54D
BdmGygPMkdA2aTR8wUjI4M1IxA6qey3ntmM9mtM9aCUyVsPFLSymXVUNhfOkuYSwjW/TzCrBjRuc
vui4rFC3+nlKSBo2OiYVlS8slg35nfOVZhoyvodoZHST04aYySFe53Agz4rmDbQagJjwcCK07pZA
rOhd48jFnpWdfunIIkSzO9a4WK7PxdmBKoutlXKASX9YoDsGGSV/HrXs4aYoNVVavbAL0tRt+miG
gCGeRkwsgH55eFMO1GnnoZsD5wVARWgqMVwdOnGfSOtvv31OxRTzZPrES5r5H1t7vP8SxCGdUxwS
kaxSvdbvt5t7Hrl7SdZAwcEcQlxN1g6GarCDax1ww20mFsHhgnmgYdxBIGoVWzVEjxf4gb6AHvvP
WUJEvn54Pw7NjUgK9+fQziNMevHg9D56xpQycvxNEqmXs4U2qnuLDLocftkg0VGrNOduWoIW6KsX
HRIDyzlPpN6aqFm39f0cDxLeYvOlPmrOqvHL+WEEYDRrAv1iguRsXdOCaBxS5azThP/XiCpxMN1i
ZTWFmasIDZzYL3XAcrTsRvJjUThlgcI6fR+FwBCsyRX2d0MVoDeX5fjSwjHRP6FlwLSBIsuPPQs1
YIYevtNTDMFufpelaarAGMBXNUno48Vb01/PsrRfuDKRDEfEed/u5xfSMPbiPBeJjWLeo5XjYCZI
XzdzjCCmo9UGYlxI52I1swKIe5837ugRSzLadZ8fnz9VIVd4rwE7kw3ZqTevR83vm3z/FCvzZVKc
4hcFioVUrs0JMuPZ6ypGjz6L1/U9G5qV/uDVMhmlBN+aOojbqueHCwi0DsPT65GSK2TUxT5r8goa
fq7xreyGqRuswUcxwAyi5Jn2y2yIhMG1tScTpRKYNX0DIMgRw1aAhMxA9el+Rsy6diY3L0ZT5693
GU83th5k7Wlbp2MtI1IjHSvuQAILV3EpD3/NTDl6/PzeMVt1hM+VG1BYnpusHBq0UJvdegjxPFfh
Z9ld70HdNU58OD31ye+dhmylPzrAXYVIMX2c3fZ7hlEgc4tpxVLNTEIOsMeS88Bd+9fUnBGkD0Ys
6DshnqeqoAXq5pa5CcNeHuABYFqpEcB0pXQPi14W5vpOKPYXvqgwqUbg1J9w1F80mRQpiXEp8575
Jiytcbzv1Qil8uO/szpUTrxowE8Arv1RCiG6CCmWu5YXgu3vAUJtAl93T+9+JW9NTg8nR0MhnNbc
GznTadphRMDdX5fN9AgadbgSD7dkKepUC/YTJd39gSrUDNOhKKgoBpwP8rMJq2ldQfAp+358Ki6B
nuBgW1xDgGb5yLjoD/3FEglLp+bttN/sllx4HZxG00qte/ksCLfWup0UkQ7I+JLsVXggqWwBBQO3
fEq4/iTT6ECicuppBo8zMfffVCbscAddijiMdjLzdF03tjT/jweNKe2kYT0UuLKpH63GzQ/f0n7q
nM8dQ4EMzvK5YHiSjEQECj+c34u6GCM+LCs0au9CSlaeUwiL7/Gwy1oiH1e2NNHFGRWEkPX2uXwV
DJFyVfb8AL79wQhqCawqaqMEJmCsFAXOMF6du1AWJBMvmdOAxXXXvmzvID5AphVQ8M4LRSAcIBrW
Mzyv4lLTyHsrDMlVP+5649CnyFr64oPAo5Jnim4yZ7X2qgc24qE7qfDnmql2VidRaTmHk1guzVhN
YZ7NRmHlMMVgIUjnFkofe7Xz17BQtX9AmnqQG16ubCUXtVcqI2hTb4ltQgUFDufOUzpnKj/XwdEL
y7Yp07eep/362d4e0Yo7QRK+Hf4m25pppDSeBXBrnHIQBvubV51ciSxNT1cridGeIYCOhdrnczLP
Y2PZyzquQJ5rSKtmn0+1eQ85s9KZHdfnFAsdhMjAfWpQMIVgFrTqtq/SdZWGfBOWVbcb7VqhDwXG
D93faCk9zT6vUqJSkAeMMP7tUobKNulSZd/DSxH5stKbZBMGa1oB/CxRTymt1RthdpLlPKQbjYLc
GHk6jkNW+LYLyxxcORCkO9DjR3vMBdqD4QBHvXK0KGJdGWFFj7YkvZaEh2ErNaY6Fypa/kS9zYSo
I8SQyIfo5jC6tdnRd585En2hRgM59zThvuA6UsH0Y1ax7lmAnx8UhJ6M9oc3/1BgjqAZ4wb/dw5c
dlUJzMdZp3wJu8nyc/t0wc6PgmHm/BYenSPrWvEieK8PaKu/2ztvzLeR0zJXQPkrZOie6mTTOYzs
GPWu7HvUqgZS3duWJf3CUHjT07p8Ymhu8hzHLYfMqBlDy9yTCgf/Tfx6KZoeD5vmcTNdKQeyw5SR
9uuWtTLpr3LzCW1UWDmlRQ8lt0zF93JkjwgU2GuPd/rtP8LhLHrNy+uCknZhnO52gdD/vXWAtvyA
SgMXJOB1+M5kZZjC9RuWVj+vYe/fb1xxI0UsSOrsXgFUcFUtTcppVBKUho63qH5Wy7IVPP9hVtIN
Herkvs5/4HBBI4Mcz5Fizvi8RCxd/mE3uSUpqBFvXxBgf/SrPa0tdPJNdRTUGpsdgVaMyRYIItWR
ZJxk6WMOXw1Gac69/ZuOqChx+DKCTiRgVRZO3d6b2PbJGvNpuGM7WFNEG4G16+hGDOSv8P1K65V8
bGYIE7fRSGubf1a6CeqvadC/TK5rw4GUyWlQ7RQHD7QWHZmv+GEn/lQKNst5dv49u+k92XwtOFEB
LaGMqCf5uRCyyGG2NAdCs5yZn3Xu9RdAG3qqA4DLjLagJP0O9ytrqnxfitvW+7BM/C0T52UvSoM9
JoYy5isi81yniWU1o0YQG45oPdxpzKYfjK5c8mrJ126LRsxii7wTxSzDUvYo1Q+3KIJUzOaQJjdz
aeSKULswqLLMvicb9TKQ1BKlEeviHGWQs6BH7IJfL4YneNF+9dE+GYEdSbi5hLqBoNUvnMF1XtxQ
g8Soaw5yB7gkOtw+uq9yAbHwZqUCs+RJeoeEnao5sQF5OOr/6NEp3voi5xQ3UKzHV4IjJ/gZL+20
KSkjGCt/5cb1trYSap5trAY5MjCkTMxaCri6lwF3GTsKHxLpd6UDEuma67isD9Tf4eluLZjpnKEu
SyRg9PMgCWrXh6rRdVF5ZXVEEjmoamsCuKBzC+a9miLACFCHHadtSF31f9cf6SlihkHr9NNKd15M
kpVEgJZ21GrrR7n8ildTB33+6vwD1tWVq+h91c5RafcIN2qRovHHEgkSADkLj3x0G/FVjlXrx0fk
4WZw6N7DrGC7aJL71T/hrlA+g0WK/Am/zCv6FTVbclfBQ26S2mbhfDCJpL5bF5DhCB8O6zPANAZc
svAm7PmxB9vp3dRVx8QMyFVRllb7wOdbaVIqZ0VyhduZkPaGNX/z5pn2Farvt+iApwuSeasNXx8s
Rahe0rfOmtviLRpRYDqeGhA++eD2iGhsv3LDVPNb+/oJwRAKcF3TH9/rRq8s1GGzBnXdN3oHJpW6
tjxAmCmxWs96gM8xlM2euW3Cxuo+S9WlBMGRvK09L/EVH3WJ9Bgkz+3T+b8INBkE9I+f/ATn+RYs
uHkfMqlH1f6u9wRNkqrTFFBh3otLqJ4qHFks4cQ/1005t46pmuB6cPU8dRodxKPteuhNh6JQ78zF
dBWOUS2FtjBeloSHNz6oWCjIt8odVSt9KArwIyfTXxF3aB6H1OQNlDB5RILvLMLnGQFySuvA7Ud8
u9pKDJABeq37++SPjZ/XgiL7HKH2cKKYaXGDMBDYzuG+KhKpnCit92/yjkhc32spWDnHH3dOkNjO
6Tm+ToKL+iNcIraIdw8SutMBdXb1LzosfiVifWrx9xUE7qtcHOHBduK86KXLsQBagcrqxf1Axq4Q
6I/dwYyrKnqeG+bHVPA5k8wbqyXIyzjE+mUu218H+JAYEannJPfstTWyC3EbBAPr4dY2XBxmF0w2
ibHgtzdP+zyKeehUQNgd3kPDooTc5Yc+oqeZhZa1BfrWVeZLH62ITH0Pw5WR9nJ4mZ3xRvouv3pf
9SsX1+rZwgkPDu9uNwr5ED3yGsZwYE7Rl0407mV6Vq4fpaAI7fIK7mEaqbhticrDefQAZG19tEdE
T2J0nCOA+BB92eD6WNSeq31LUyPMApnGl06Ldc0HuVa3XAYCPsJ/1+FMgdj9jlXkPWoQRfOQ+ecw
pmaf0StqVPddBO3+S28YVS7XS+pcb1uWfA9UUxm7/zgO11pIL1lFUw/KTOGQbVBFoef+iZQnlGyN
jQ29Hz3iDJmTcsQR+zAQL/QeS5/GnMUO3LovtfvfXH9b/Ck81DG9t/UNe4sRGEZd17OtVTE4QBv9
gdMYoWF7cGDUZq+/7di1Q94ukQggzKdst55DQwhPoQox8UI8lVKxWZG58lQbTQWv822nNxJV8TgR
3Iq2Yxn4f8l5OJ5rVk26WlbbalfiAv7455EgrOLuIm7P736v2RxayDsmwefbEnodm7CyQUMP/Auc
9nGvAdPXYskbWRlPbpLKovUWom/pw+ddMrSu0TZyowumP6C2SZQl+cQuWYpBrDFJuoUlPj9fydSq
IiuTUqoU8cjfm32ctxVsA+OcET7GRSBlrDcfeaIMwX1yTCMRTsf0/DfAMjcmawcDtNXz40NVcDYd
j+GrCNwDPUpEQRrXLwFbxp4pxiOQYMnv3H4hlxAC6os/EOvzVu1hf8yQ6ler3cFtbIMITCUFdnKe
TxcgsnbaL2LkcyjRc34ljCg6OZhtMux9/mugyC2xRJw4l+QffJs+s6KveFS7KW76DdFGE4FupNvl
5tqpqed62SZ7zkdGypjJtKDpFu3klU/aoOzKpdnIzV0OU3X+hM6kwZExrC5Dm92GEl/HTnDVT8ce
VgMtvu/B5kdDLSc7oCMgnn/uoy79dn44HZSeTxYa5V+BTCvcjYSC9m9vbUSN0Uos6fP66Yu+d/Jz
Z3sb1tk7F6wYP/+llOPZjGf4XcIef9bQ1sJw0fiFbTXnLjdrGFEznZumt5B4vOVnI2c/8TXQ5G0p
NlbwycDVJ/6xOW3g3Mnc5AsjbuTB+INDbfZPfkrpb016UJ53rHhr5aZIacIby0FdEihB38MvHLXZ
idc07V+2hJMPMEUey3N61AJ9rq5uKRUeEMvF+SofkdrJFx4I1DK8++w6vEFprdDo0QsK8blNQzCf
aoDiuPTDgQLsQr2DiigHLt4LUCqM/G4Q2iKagRZfinI6SXgqD/kfR9EfYlW9/arb6Vs1mMxu2oIw
mVF2Vpl/UwdYW2UQAbV3Dwt8Bk6rwe2mxzoHjd/8JIbX4VI+hf1FTnWDHpiKDU77g+dEz/GBFwE+
cyaWmhSXj9+VbjQy/RlLLhfr1RYSfpRWco2Zb3jjNKs89+L6doyrr3hd3930585v/mKIraxZCiLc
KWQ2JdaCRFWHtOUj+WdTVd7LEWVkvUbPh3RKnxC4772fj3gk6uqkktFOq9CfUVqsEyRBJ7wJQkV8
brD/7E2EsR2Q0QHtZmmgjHtbmACwCfPrmM2X4/T1xizoBdv1KoJvAmMroiPwdPPAy6xotXz7BXCt
QmNCa9fzEx/acACpVnCax5JXyLHqkEeyNNLX//eWrXxkpR3heOecgPwg+xgi8IDF5pBT/nZ4+BcX
Befj5hXFnEcTtAwHfVEwO9jLXNfwlAFmnVXQ8Ix4FAN6UnvAD3H6m6Fs4eQcgTOppak/pu7JhPCE
cD1rk5/LupP+3UYaoDI/OiNyWaaWd7kMtOSzHsl5rqZc1AFNY2PFew0KGvfOeWXqb49A1TdC1dIn
qzBal53hTcLHndmSr/V54SJ+yzLAoSQ61qh5bVO6OxwPdhpCoivh7CgdubWnRJDDpJdeGKVf9wPv
8Jw9M5wwaRerqm9+tgyhQF9Rgfio+xMLV1MbBCITWc0DexuZF/npwRpQ7mRwLaP3FsLnjvwX97PC
nDKw/751FreZLSELmyr18HK+VmxleTBriYYDdzgIdmOavHgiBHMuX8fqOxOtEfkBa6ErjYb72JiS
d46o/jWep7JF57gYWdhMSvB/XoivTwBAsDZf6SwxqWSo/qA7VkbyXE51wkS7xvMn0W0iPeyvygUt
3tJlG2nqD/la8Q+D9fO3iiSvZvzY8gbKFxtHKDCB2w+9J3rjkG515EFFXHTcu2HxeNgtCINMuqIT
cQSFbeCCV7SAOstNqJv4ySpgeCBMo7HSyhnk90wYwbe8OvWTapc68j/PAS0R3ECP1UclaBcHI9zy
DtvfE9jySb21cAhONcX2bL2PnmtoHkLIPMc1VuF6PgO20fkXRlxo5iw8REf3Oy9pG53T3EWWBlpV
3ggKrD1a9mPFQPaUzCu+qxsOpuQ+FJ/BkAa0/BtFc5D8MK17DgoLzrYbMzNxiDwCKHKEAAz49uWw
nMBVrLGcJzIgYckrv15gMsP+RtV9VdI7CQQCcSO/HdGs4RKY/40rjAEvo8GrQrWYKCP/fcz3lz7t
2Rr7G+D29GPz/wtBA7Phed2o/ov/rF6hSolMPOajE8t0yblDjScEp+TYHocTe5H0FgowT4ck2hP6
8IdCsY2f5SMv61oRlgWiWUCNBapJgZLMxghasVvhAVUCvnyXf0q0m+y0wEaok8i+Wa87jP4Jbsd2
30rmV2rk49h7bFpLED5riBqrWD8wZfSlalqNhg/knHtMAqZhyTdQEf/fJPEJ6HEMppr/3C/bolz1
diyl2NrSJrUctzTvHSGf208/sVXImuhv/IjwwlUjXPf/KocH12O9hxIMWaAy/NGRfyPajVuiMt7Q
Hm6desnYq97nY/0AmPdCaek/FpVEe0mbIOpH/0seDi9uv5sGVehtNimwv/CAraJnZG6l46au1Q/0
sjhRPq0jgCMHKK0fhg6WcRw+IHgHsQlK1GlnrigZoVuNa07lfSU+r2v1og4jbKBCJwHmFDl/v76/
0qcy9fnFFblZRnVjEtkCMwLWWBCwNd9o+kjstVGZAqEunaZ4kQf6GCezj/ZF57JrxhMbUrjzuZnh
E4IPgcv2UDUVnzBDxCtuzcL8Ec7bjv0S6Bu3cxIzDc/4HIGAEy7dcr6LSD8G7Ra9Hk64ETsPowTe
4ZfeFj6XAtssliO5xGe/TqGboZRort7/0DcaqwLT/JJpRqWbH/mdyGAsNXntcmN+CGSGOpGFDflM
y7Ic7IJEtn+X4hz+BGRSQj6+hZNJJycSDjP+EPwtL4wOTeOCEURI80Ac6epFXa7wGMfOAbatIlVY
LZIFbGKbEJOH8kRE+S5S75tekJTLJc9Dy7BtaD3rRcKwobWzjjuJhzA47Xg/+0hh3c97oS3uCbv6
O0uggKJsoTDVTIGCB+7r+RRl/QvQX2JkxLxHgFBPOEIku8ZxIQjVZvk+2KViLb+6c/QJcawgD4ek
LNbCaFN82b52Nhe8gdy3QTXbMm6YErzkzec0+N3+KLsxZXttjsY9MfEue8Q8q+6DIzPD49jPwrkW
5nt2pZqRgXQxU4B1CoYTTT6CewdXISxe4vqfsF6d8gzZhAlczV3lwzhqaTs5x/hgPtC5SIZcDzbk
Vcv08rAsaA4vl2wJZSGrSmwuZAvhYNmigKxQGBtCxi+eElC6O+CSJdDcs3+IBk23lotmkzbv1ots
+yOq/U0StZnrehq3KI0AvNyDVp/i7yOHqS0rAXXsobiwob2wRhF/jECLQ1FgnHccLgajOfApsdib
I5/8zJ1Dgb48dZAaRECD/hSeYY/kbiwLnUT4f1SZ1gCeLSM7ehnF554KHV53cfNeh6X/Pir5Wjvf
qxBCu0/mhFYqIhSMV4XBtOTstSIoepxTF6eUWAHZ2FMKg8SerwJSm5BHtlYuB1GW9fOo4cKJPckU
z/ty5hJXCfZkcg+8nfXmNsQTSpxYMHK1kjsblsoOg8diHm0NBWLn4JX0Sor3/Alv2ewYlyqR67ip
LDJ+eavhMCXFtatJlmcQFVbEH42npvCUgnCEGZWM/psd2Nywj2isiAkkrw9TLnj/rMcMEqdc20Hn
h73TgR9u8ax91RAFG0+aL2kX3wss2iZXwcX4wRnvMugixfw8yyeAzfO85IaZujd4SQw0ZvLoUlzg
tKIX5ll0iaeOo1RSdp3bp1MrIl2+UZDjzEKv87T9BvaYodkkB00NJz2E9B+BmBDakSXkXXb8HvlQ
pp1H2rKH/hyV8AWGL5ABXbMheYpiiuBRY91OE4Z8IU2fT1UUrp5aUKP2fnkH8Cg+dYNPVGv/QpA3
k9yvGbeBOM7/BOZ1elofu7oLIOob/yTrhA2sUUvIlY27zeKX3watIRfhR3f3v9q9ubNvKm8jV5Yg
Pl1Th/9fD98D222hy/ay/6i1WBV956cvg952LKT8nMd2JdBAn88J3KPNlx4KeL4T34hGmF1kc4Hl
2gAFSI4bIyGG9oLD4IqmnjuWjxuTgGXbs6Lu0Xner3cv5r8szpP0Dh754r8ZZdOKjTAWE3WhzfUe
LFFowLWen8xNlv1bmLj24rwHLzkzz5vwLbdj1NzszfAqCo+HUqcHELF3UOR6fvW4OI2wx0Hbsky9
Z/oXuqpvtotgUY43+caraHIEgYcCkQiI6/9k0Ud7RcA1lGOwrQKHy1vOpz95yfN5ETw4+CrV960I
SnpC/YD9K+9PwnTnNBg/Kc9TFvsdX86KSyKkh9UlXD219fsbF1ukpUBFWivFNE/jiT7VwAI+3VCV
EV/HS1vqeAnkIeGniBS/UMv3Y/68oi6u5dDn/jYdKlaGHWPU9O3n19Vt47HIPeLZ028zHv2GKLTW
sf70XrOQ8+m2K8sGxQmNi1+i55qdijuT3uTZJONG2TQS3RIQQO1UKsZyRZkwJEhmjWsZXIijflQl
0AryjXVbxd8J79vmYVu3nb2+ObkYQ0VAeVagY427K8YOwuq60FJ+vHUoYF1XRACHfXs4mh9eA6u/
vNkNYUt6IDmMpKm9xPMfqzenjozTph0NulVuxmnqTqSAw5y73Gl2J9SxqqzXJ4BCdLtq3Jfij5+J
OkBD2lpyOAVFBsAXDr5iegMBaI1QokOJSCf6HymLCt3c/AmHU/hP6S9fAK+rPG9fxIvf2pKOVzex
vrDozxPIQ+fJoty1wlT6EWPrvv6O0hgOxSVKC18UNNO/UuIGrYI/FNXOahNBNuoYYz8Zl7jkQhvJ
NvsxU0/bKu5UXVLDN+wAK8UVfEgkSOSFrJf3xfNn3lcVf4rF3tM8J8WXYr4FQsBgDxoD1kVSytj9
BeiebOHVBacKmZYKs2v7jNKA6/y/jg0KBYQSS+lqPjOHJ3AlTWDj1v5bW1ZRiFsT79rl8/0/tCll
Azm3gCn2Z9wPpt88iMQ7HAFhYZXQKRTYyDwUis2YbtIch+9KoJv7+3LtkMlwMWURS//kVHov+mz1
HvG1xjdwqsTj9IDyyAkkJlD8MQNBd1ARFu/uonSYyeNBmoZFiLf19sQpb72r8cFoyUSxUwsHVEyo
S7Kb69XTq120o/BbgHyMBRaKtb2iDmLYIvSIo2cXnKMDYR0yOO1B1aRsCsgF9V7b5ZpMhioxruXt
FMeLqvGft/khB7P86cQimDXHyDBI1EG5obEG9jTnbwKSxSR1NjgoW5Fyl6TrZhs0tuDywVWZQLOa
8bexBb8t35pybea0ZEe+IR37PaRutpqDHZu3DrkOybuJM3HbVwgi+Rg53SUrJ8ODYJQQfxOwpkYf
HF9t+XPzYZiV0Y8UUQ/oOdLc0/QbOivRYZB9aqqI5r/3dq0jUQBmIybtS6E5R8k9V6adeJon+Xs9
WZbFL92U5VC44kS030jtXoRUgvqeJpw8NfgrcihdGP+rvvec9eKj/b2t3W78Iy59mAAYcYwZdvsw
makvm2QN9Ex78TQee+ia6K9lfBBTBSukWe9JfIhutAx/nfjLxjra3o7xbyxB3LEET3wkKtb2olVB
4AW3nwR5yMq2zqmLDGYyF1bdhQy0c/cvZ2QpWZkRVRI+nHsmjUSqU2nnfPz6vj+nBgDBgXYogT+y
9zy7BGHheSU/fu5ZYkykiTvmt/E58Z1hWHhewIJjQdCaBsa7Hqj9+Tx6KfgpuCepmEgaFqxlQ4fF
UU9QVI7YabgZg52YLa4odFkb06Tpdl5xJfbp81RIreQXR5EcMu0boB7O3L1Htf+V9eNOKPTbRMkI
KUbA83KXMQzwj7pC7Mi8hU8HuC36uIAEgS6H33/khrtqRwIfjL5hH+xfKyQSqiyxFN+R1MV8qRlh
sbSIP4Ne/CvHmcZJo+FNNj1BEZ3ixv4YXazWE1tGrkWCSxLIRiNzxZBstjYPzF9DwJQ9eDzBnJAu
SdqqETj98tlGkziPTwauR+vma+KNNR2bTnMplnqbnM+TfP0bkEe2KHaWhnmYkGMBIJrjc/QMOmeG
uaWsk7St9IAzqCH8WVWCY5bhQxDiBLXx6oWE3YlD9+oagZ7akZfsdZaJlIIGhNILmhDEhxgMAUUl
eyWVeBnV1a4x3D+FWkCBBUK8Z+O71xsgUa5b7vb6eLXazJed9FNqESqYfVzlZ2i97USpJ+Br/eaM
aeeQn3kdeF3L9rQIGdxFLbmVnI+xDhkuk8sTOrzlAVWFbcjjVBoM7iLJQBtfegSuZuo3RG1NaUTX
xROPwOYuS0ba1CEqM0GorxSRvKem/dZ5fs7EBHItRt9xG+DXbUYpCHfIOWe/yN1ah1xKbK/xnKex
dJMalxFGVy00y5+SvNMjakaetIMSeTcWuYfVHsOv8lRdw/6XRndlZAY1hCeGLc7uVaClHfDk9/aG
gDIfv4871pUXIjTkxVcBENBttvDg/Gl1OOYyR5wdhObJlUrsxPKBZ4zItMpJ0szfvl7lt+Ecu3Xv
7QXEKjH965XjANSLVJQDxWVo/CF6S2s5yCPyM1ZbUacWJ3T9965JZW4qTZaIbRlhq9WIRaS5Sicb
3lCc6BEQhx3GXWnWDr56r0WgekdiYR+Tl7K7QVQcrMMQbhyyZjjRdyX48kmRvpwuOHgRywGWcwxL
ChJd6oWQAAri5WrAs6tdNVRNDBo58iOHGWgNVmxkJC8lK1B7KNzfL0+kpRi2o3HhJZ3/ogTPNxBE
CPCZHjokcpD7Nqu+kQWKUceE8EiXTmRydijup8NDvWuGGH/BHoyFrQacDI+AaAOvGO6iXcfxCRLQ
NKNfzzyxGOCotQffXNe3695sVz5ndI0L5pnG3TsQZccAUcJCOXCkn9LkqdilBoZHwKd6FK0HoLpv
YHh9F9Dz5bHXSeu771ZKhai8+YmMXoEVFLxdsFUAVg8oRH8trBXK63vO93GMvMmuWG1cgX/yM3sU
JJbmwg12UDAW8uGBDldyNeFDBSTYEAOXtyr0VJoPH8yN28sNtzGzGnNh883WyezTqSX48wnV1Nuj
vQi4pRfZBLVyX65QdNHB7EQuw3fvKV+ku8qmQ6dUI/4iQq3U+IJ9Re99a4eaTI37sE7q5VE5LtAa
Pfrp8tY/9T2X0YI0U9K/eNpF0bmDRu31MzPdbIr23buKOnr+ZZHK4tWcPtAc398m+sGXq3IJnr+L
Vh495cd8b3V6xxmjes5I0tuWfRWmcumeagtzoy/wKP3gVaro5rRnO9p738mcXStFrOWJzTwCSHsw
7zsfehfBxiEKAe5NpCcDI6VxZetCzD/27T6RviAt80nrCPa7AIP1IBygSsrON7kHLeG8/nTNfoH+
zZioQAqmF2bpasyKd5PhtZWhGAT6fegBOQefHhhdYMEeFIONPX9TM7/QNOJNmFoziz8crV6PpAD5
gO9xlYtYRUqRhKMvctic20iJssVNqxjegomPvHnScLDPywpJP5tdn14gnf4iIp/xN/5uMVfhjI8k
PIXD/BvPmstK7rKPW95Bdl9HRfPzPtazxvkeamM+X8E3k/JgLH5spghdDF7c//I6bB8tPctPtbHf
Bo6y+tE1aUrekgvZv+Ifn5kSla+y0Hg6aWnsFMvw/92RgaYmWcga99XHvhLW7Lk1RKSJ9NxALq29
LJL67V46KQ0VZpOw2y5aXcs6+faDJsq3mpHLKuwywgb5gt864XNekZ0XQRmkOMuqbmzOwb4SxbqK
iROJiCes56tq1E5Zo0/MqeEKFviiEFX9su1E7IajOf8sdVyD7uSn0Nebc47qgGoElppZLpc464f9
yk7F3qMsgO5ECQEnpPtnKLNkCSAfUPkkfzCDwOOYvIVxD8JEvbrK+L8CBlEmGT7qU1LFLxS1nYIN
6ebDUfRc2yCu45nnuyziZ1XFsR/HDhTbpCzvw5q9NkBXQLUXfnV2VINKLMbktCPXHuZxFRaRcRaL
CJ00zexsL1twM1dHrsxh0N9IYPuAtpyu7JKhWFUqpozc3dTD+OFpwf3Ih7wItIsrX34kZ3wba4OI
d5S53Cp2kAf0769JjhnVpC+IR2TIBJb0QmBP+EeBciki9JkiJ7rclINOedBV7rB1YnpRGSzb99dA
qVO0Bs1rJHCuIk3/7uILoFblSrDvPc7qR0+SzuK61SJy23Ynxm0UuIdsgCAETJXIEtPXXGQ2N2Gh
zri6K9ex1iueb+WqujcPTlQ1wjtbU+XKgdN6rxt11ysC44BrM9l9qv6tnH2gDIP9qOIirCM8vKmO
ST/FMpHC+bcPG5h077DimqZTQCKU3nCErPsfcAP5+PO2ORfY4G59lawrjUHYreZCinbYXy0aSitG
FSJelNKAVsPLMa/xm6/doC7keYA2hdhxc4+JoNLeypwjc89dGyRMxFW3lf8vTu7cJXZcKM1zHvIR
XgtVqrmN0l4p0F7+ugdKVCFzda2fKBIeFxVmFOGeXyZLttTjswNA0L2cPP+iBsvm8Q1093jYZLub
i/7V0tIX0UvPUOhY2/4PkgCWA+8TqVdh2mJCo4Z9/lem5oKdaM3NzAptwh/zHSzMnVh3bvIzuzv/
y8Bo7/gexW1VXYRGB2MfmUByZo65OyDJrbWmIWsmWS3NNlRvDphdeWNEgP+I5q3li0NRXGb0tlwr
U+cW+WV7/ogyHSFKcLBkYsfL4hC6VFMYhBWpR3OJlI3Ehmm8bOmOyngInd6LduccpINzngu3yO8C
h0yTws6/MhOn87NKEUk4iwyTzcHomjAeeZ1wyqIsbK8RnEl5AIj7JbJxhLACv/ePU9drxUqoyS9z
c9I4b3OY0Y+Mk+lI/5HCrQdSTWcLF3xSzB1FbWvQETXSm+VSeP9FWRszXvsCgk21ir0d93GSKq6v
wzMGEg3G800+PhFpkrk2Y11DUqPAcv3muehtaLGUC0t/7yd5jxNH61ye5uL71e5zM6YFnpysGkwn
8bup7NwxHzZqx9lHbf9EABRlCATCRpTr6wWmYZ/2SAh8ENw56sBqkdS69r7Tk9OB2zZY5vhUl/V3
6LoyloXCvTsOViFvruZ5la4gRhXRYF8U5yvF8iA56EgWFOTe7l9B7ESTBV3hHim+1MKnOMD/p7LO
Wt2WtXC4UylDywjcw+noh2hJjgz+9oHNh1ldpkBNEdQL3W20eQyeGNUtI6pFHfYqy13DRtwVSEC7
mV/BHB4wVKNKhhou19RO6yA+rcd4JCADfHFfTVbU0pdvO/Q7nQ2aPw9ap8Mfnp0B+yYc3nmTor6j
zKKgSKOKSR5WKfizKSGAoYfSjThicOHxFpDke830oJjq+tkL1NA+xQIp/iysddC6/qzCRIfgOEW6
lRfwA6yDWDuO3IaCxC7YrbXVnXiN4Aze7174QJMeVfAd85ldylzCXl/jMJbSlm5BYGvGNL4+UG5O
b1Bdrt9bJnaEqHKCXGrPw9W1hnwkNI5i9LY0n8Q+/ATIQoFXnJAlEXO5DS2IaxRbQBoj1xaqPPeK
w296btZr1WjOW6/UgMwMps48merxYkbtQrsjMLDTAF+vllqJluO7BfrWxTtBqWRBZ2chJASf7AJG
KDEPcJx+pyoLXPqAK/jNdICXiOKhBjKiM8ykI5DC+4ZYNxwfdIurly5gPaIJ+eJirTxXvfIkNB8/
j8lfB8np4+5sUQm5iW+p/ph5i+2ZczVYyjakiWjUUquPmiLzlgUNGT5uh9y/bqX7h5JlY+gSSrNO
NLkq+n9qNzl/fVLmqMmAR0Vb6M1LnePohfcAQ7hKNxp4fXwadPGmXbyUNJwvcJ94fcOV1kGRlTv9
MX2PS6md5OU+nyjxVIy99umsGP3Zf2/5YqjGVXS64FSJOXCCz/xlzktaH5+H/mqsP6qtngKUhgXT
BejCwp8t+b3RarspzwX//KO2NKLy3jNzFMbOVaJ70kUp3yCU/+o8DXr00v74CFSo9NjArqEFQhxl
0PmraLvq4GBThqVvyErtsGXSlxl+va0Ea/NzUnmxwmcNgT+6xKfC9dfKf7WyCXX8GUT50XZUvPu6
98jCk0Kkg9pc8rVsvJoASWyTVUMkZuYf5wV/PYh7uW8gXiZaoCmDfu3nob7Ll+UrXMbtERvcCRuM
V2t1Mv/21/bqW52o9apnLAVgW8+IPWH57K1sAWQPfkSQm23rDQ+F49WPEAmQUqRvvBbAmkATw2t+
GqovNog+Pv/0vJfQ7RJFv54qjSr/zdyZCqEUqZh4mwUB2/5/gRhGGtLfJfAqzYkA5mLPmWx8zOaL
LJRDvIlZgyWaLPvXVzIi1BR+4KRZ+ViFwIzgkFBNj/VEViJVxcxsRLxwIHTgplZbNhJfUbHA6cOf
SEXE5apryW0YQ5ZQQcPDnnacQlvxdrjzzMv9Pq5Ns1549X69b4nRiBhZs90C8590GlPgsCRjPSOg
/J9y4aGLf99hnirNQp5cQeNpCL8uF+DagJaT4qeDCBeursn3lspFGIEB4+zCem/zcBGFLmHsCgc3
8JROSFnS0XyZAmOITHSCmGOZno1HXCxJgbQk1joH5lVUjBBDh5agZCPHwcC4AtyeLiLmjH/HxDon
sO3y9hGXixyw5T2gJYF90eB7/OqOuE8HJfDSTG1y1injQmqUiSSVGXRg/GTNxoGBHellzpkZSntL
PSNYDw3V4Kjw8IvLdT5uj4VdYUP9EQal6A21wcS/DwSZqCNr6I1xnxYQ9XyHSb6CMr6TL2J+n19F
7ZCIs7Ss8duGkzRNhx6hubwr2OVIPtUnfz7UCoIoRkUNlGqGQVZCXuLaCrgPjQ56ZQbstcvgnJhO
Vmmzz3r7+5B3WGue+MtTmS/T2kE96ChFTqmtfKSeGTIAivttpDX90C6oaAItUwJclDwaReiMufHK
04oYxOihVp6KfqKb2uw5GpTYTgIGxM0p8co5T7wDQmSWF58D2MI0v41Q7aEeSxZWDse2XjeJrQG5
iql/mtG4ci3LHgsSZ3DYjJs/q7pil7wv5USWfy6LiYp0ps8B7SJAn3i9OfTTJDB1DvY4SXJkVmWP
pjiplB2FNYlp6LPU9DTJuRiwx9JQ65KJKiFWgIJW8/RBvXnU+IyVRFZHzo9R6FqeXAEy292Z34dZ
DaDGcwm4FDwcs/MJjaZ7KoUuarYKGkCf2bQiLnFg+AHuNMNQYZdJG3HsHQA23BGvuuSyYCyYN+fA
lzz+QPyq6ewud/JR7eiwk6rgpPClS+6npgqfjg9epUtglc5nFMtvkfvi+IEntvnib/PR8w77/hOG
OLtw8N3IHpe81BOT+QLZE9bLCEIBoT5Dpzw69dTdqVSZXXZy29vNyhqa5SWMlZrwnEfZdSIuTzMF
INfCeHbUFY9KaBbryhR4/X1lgavmDqt1KJEILgmTKk9uK/O8u6qyeKf1iGpuwlupaiuCgoQj4hfD
cE42nRF3uDrIWkFJxOx6ZQdIC8WjptvQn22Tq7nwoQ1m9ZRTJFBSjwLEI3BMlNZYJbgHIl8FQC9R
9ViaMI0DVSJhQ9VZOURRFndy01aig2DylNYUi9KfH566XkPHHwuP1q2aB8E9BblKzXquCttDauq+
10e+ZxwsUi5EixZd6qoA8FJcuRXXOVrds+ucdMoUP/T63uZ/5QsVFOxOPW0Tr0DhJL/uU0T0RWsp
exOAto6ljSXP3XPiQ0uj24VhjtRtQ3h2MGQFVyxnhkLvBjjeWkmD+1Cev8m27wB0gTkBzD5NBWNU
UjNxU3X16Mmw1bYWwTfbJmSXeJEubLnlNsKhS6GYmDWx6fOMOhNGkSdW/YeT/hgWCdLTESygYrUT
wCe6z9qxRDEQCHiKMB+/5cBfdL+doV9C1QAUQzhjgpto6bXG6ix+WGqDugVMooT+/ceWrMYW1Vpm
ucy2H4VxpYMNB+RJgh4JWtQqQevIzVRu3mcu0UIXwONwuxbk7ENkYEVRbLhAjKb0W0ZySoSZR+TM
bWneDGlEmnEsmzY+b9Q+J7H5fOlYRVPYMg9JAox//hQWbmjo6MqlMB7IGc/37uGiPPmTYauGf5sM
0N++VHrRlwanBZx9rnuZuLj36D4BgmWeGYVB4gXglCwYuFVG1YQYAjAF4vVTao/3b3AOszYFn09s
kj47YiPrVak0qQ1fdtoOjNMIsqt93IhgNtQGN0m/wkFD+Oq8D2Qt82p0FLo2O1AsqVEpcAyYzUy9
zSsdKi4+jyGlry1/JzA+fdSLOF8cH9cVQpi6DX9MSPv3+Z+jmq/AmfVirC9FiWhcSnlQF5qO/mRY
EiGqAhdN+f460SSBgSNOH5GIZdeG+Ec2NGwiY5Uuw/mIgQDDPearF27I69u6+Od5QGJMITvHsRpw
2prqG/pUNyx5AwdQpNgk2MtcZstj+FzbQGn8cu0wlovkDAj8zcRFrKB4BVq27b2yLLm7r/ubQGaO
k4FWrrgkk8AVQlGoLea+C1VPoLGOS67elCVjGKUShsKY4lG//+upHnhgwGk+lH6UGuUb7HWM4ljP
eW2Lln175vcUoQ2ozBdhDcTASP3NnW6wY2x57hPmbGII/KZYosoOFzCC2VTRuxi1waE7QcWFOmxU
LLZu+Y4lcQhalmWReWD2tBCrAh7541VPp58xQD88JIyNsBld9KbXGaNQxrDkHTrL+WKdHgNJuw+c
RdKxRuKtbT879q1JQ6syiIuE74d1KNZ682YCPNzVPK0DuCBOW6DGueF6K611t3TGtuvXPiezW1Km
k7224s6YH7wZASwnXiVAFazlxoXQyD9zQchZZG2dZqilzRKAPIJcQJVnZDvMaLghriohGyyc0EDD
un2J/d6g232ZMFsnw274efR+n2hgENntrMb6mMtuzs3iGggxUlfbIxy2gx0DsWotZLEasLQlpOxe
mMhIJceo+Smw3CDeHdjtlQd1WbvYDmk+nGejguw6wllb1vG3S2bgBuXpGHOPcBzHKM4NdYu851QX
lxD5VsksHsrLcO0KWj7ZHnpBAbpG36rGQosfybxnkUhb32ZnvOMMOeM3FqBmOhDSvJ67j48qwdv0
cBCWbE+4xHea8aZLZ7oT9kht462kGo159fCKZjtlTCWcC5HFmKD9CqyPO+u06vg0X8yt9h/kkp5f
5M+jfvnRTDy/DVwR9AHpTQB8Y1K4gc/zbpMppSdXo/7yZ6dAfJdVUHeNExxJ/gqEk6uTEiApeyil
puvNc5/G6e5bPhjv+5k+1dJ5DnwrDGykDwbrZsTbHMSKn98dbRctelthmoURNfN+Rj77FA25Y9ck
UP5cmoWE6m6F8AO70Ch+WScQtgW+adwyJBgtd1RoQRDCTD6pZesiKIp4YL/HWFEBVCvTyEcz5/o4
RHlbFIws30mLjb/PiFF7Kjq/aYDPrWzqj7LO70qqDdpw2iwquPuCOlSdjyN2PcKLYXFSCzLPYopT
wO+GCvqZ+3/pMFPfFJys50GmLjKDTbhfy8hr8rklCZzFUIdAbfKFNaycM/jA2Q5OE1bExj99VNlj
ooRn0MPlS3NsPBOvFKskH96V2nc2DB9lj7h2rXTiydFuneZqJI9f+8M8qytWJsOj50pStzcWj/eP
M4q5zzEh90CcnedxHuhX/ViRS0qBN1saVxmn5uLx/9PHa1+lo44XTT4POLRFi0tvDpD1/vBVuDOT
Rl+U1SLKCLN58fMAGSHHbuRvSQA3zFcZrCanjfaVoeecwMw/nzhGSUi4hQM4squZ6UFM6wlwlIO8
qtqdwSXbmJLI0OYTWFq8e3Tqa/L3n7tk900JOuldIKy1leLxo3fr8VLBAJrektXdrW7LsRuWLDZm
FNdSc0oCcD55+K7zNrNTuUWKtRV6Yfp/9Y1M8SqfQfQLh75+LM7nNf6f7RkX1nXw5CGpkd0G+tR8
ZH9MC5fnsNsZiyx2YIOYYaZfnl9F5i9KMILKIobUH37pFwBwNv6iBlwHWtP+tBmX/u0Ij8UHafMI
tfUXemNEVbLQDa9/RQlVkHNQaozVewHvX5xpRjAbGWBx/mZOb2DjxuTke1fmIe96ui2JyjdU8age
ExxIBZWfNyEQQpfunR9Tw5/NrO0RDFQgUAQfQQOC8RrybllSZ55yVlwGMvbMusPeSx+a3UPFU5lQ
3XeOkpXxm79amI5TTqR7CQAsiNE2uAfuuFc4peUYj9aWGFXIS3eoRtF62HrKONN0WJkuRY73+uGr
EpfZnphxPpY00CMhc1qPe6VWrJw5qPfhHKqumEqYq6kIqTJ40YMmkDlXYDppC4jfULsDRMvA21dg
vvPthjd/IWihEk1kfAsdg3wv1Kxdhm+rr8qMd91yL+1FCyqMMwQQjGljJzwEmQSZVaVW6CrVwqpG
R3pPzXThHrabpQGIwYEJ2htNrsLcF+v2tpinSk2/ZCg4pTwWZMBRa5hO4RvomWT1WBxCvN86zrEX
DkU7fcorWVIk2uRzrlCMaBnJXp5TGMxDdkYpYZmxaI3KkD3Twd8c6QkG+YnjYX6rh3M/AB620tXd
Jzd2TV/hZE85rrjXnCiamWAV37dLj1CVcf4CiB12np1CEuXZXaeEaumQqOvsTrqWwLL5l9p7j0l8
dchfsUwXSXNlcDcsGI/M6/z2HZ+Y5Q40gQdqpG/TEr0gu5y1NZ5iwYE/V+iMfbdzVZJ+eifYwkXr
PGA0NMxlvKpbBSbscX6ap7U5ClSGepIzJ+ibx25R3dgsWml0SpNF2yreIDNGXyGG6HSmwFAB5UF7
HgSwZOmPCaLLkz6ryxOeH7iZBsFDWfoM4+3aLb/+XBtvgACMA53tR+9A3DXGdVRFRRRZL9DbcB4w
r3bQJFovbIoyJMvtwcqDqk4mdLNPM46IrY7MkM/726hEeo2Lespvr8RPOn8GWJHrIcQnEveH0+9c
qOCCrcDm8RR2fU0N2XQcuwmvIz5QnBzalqL6tB9Rka94qjrByN6lJR9GMQvdi4zXiNJoCFHkK/Yd
q2MT1fzAuGFe6aFrVtUQgBzbsl431xviRYkYI+SmJy48Nns07WW9CtHuqwYlfGS2nlmQ2tAuAdaj
knNq2WWyUwLowG2JlWR2D17/qCVjWdgX8kKB0hxbuirVYq94zE86wLFQYcTgNJcUmyogNiN+JsQP
YavMfkq1QjvTIaXOeDpWZm3UGNvihGlyPtEKqiJedluhCjH1Vc8v33YMKFGgR/38E1OXGB50WF0l
wxiTbLng74mPPla7KPE4EpL25/THHKZ/2UmR+7g6xsN1HAxMjELcroEaJc7tlEHU7vww93OdE7TP
M2Aw2YlZSMd+x90HIUm0UC7ta9Hix+Q7mIeAzU49x3ZhQEg039XepcTAwjNNuTKrsbzAvkrTHQvB
R85E5Ot9I7FRLtZouz0aNxAlom8zDEX1SeO/VlZhHmFSmLXYyJUbcgS3tyGhLu5uh6zObu4beIXO
AteABuHalOUA8nAqiys3MKaSFFEg9JiHHJghfHEF0UiahzlgVTkmEmk1joHvKO0Ums3d5aI5zdYQ
elwPeZdm6t/SNi9IdTGJ337vTpI3zXhhm1MEcmlTfkI60SZiO2RENpya1oGslp0h6B8uLcurMhmX
Erc1xSJf1J47b59uJ4FpiXcoSm7/P9C+nOVa2fV3AOZn9TthtK9q9V1tLjskAXb2Y5243g3Ijse7
juOFh1NM6ufGvsX7hAGHiA0YHzHhNUmx+hZjidesoMxNs6P3Ro+KimOsZm7ipUvnwdvroEx1Z4kN
671q0NLOcl8x6KyF/NnKdLx9OT7T8f5N3Yo0o3rHUOp2AB5PM/ZVXbRiWYDh2T92wRt1kY8nnmOF
/TG4UphB+tPig15OHnGG8tExiNdIiiG+VuxnB9ZqHo5sV7k3actY4fWwAFPVkKI3IW9CQQy/34/s
jy96vut2evCNG4+0a/9zzYN+WeKKsS4IyMyp6LEJwxPyRnxHL6CbtR4HY44mgt1yDUb4PIm8pmbg
wAIiUu4s0qoe5ml40wAmKRcIz0wrW0k80KGrS2LhsgAiwY5IJQUEvicdnBHBN6ALpUwWTaw2dE7Q
BoVrn0m9W2uMKzI0je4qgvPiqceXNRdRIu/4GdYNnacfaqAU54TWKPbOVFxh0RVTI2pEd6+C/TTb
yyRzY6yDhHk9otfTmJXmL4N1OckqYTDUBs9bfToysqBPpTA46QvCXviTy+9WsZ95yITXCDIBPGR5
kj0sfxAeRUYnld/Ou2EfiMHw2TDDs2e30fX+//PeCD23mqjKxZ2LXl9YaFHDsUMRAKIB+VBW0mll
hl+VFuVmYHunB1hyQJ4dpgZGZQymO3ox70nFepDfi2zlC6mp+xIcreMJvtRG/oKclYUDDki+se3e
WN+IC7fq12yC4y1ezWr7auxmukaeZvIUhIKssUAFcjxQruobwqxFEoKwIGDrkftmAGbV0cZvizCq
skqZ/Oslx5nhrneuCn/Zo73DX/gizAfeHioAwa1TjF5gJUBF2BxJHbKpEouO4Iu3dXKAsOrJOpP4
2fAXJ+4OJrdrCJ2I6nVgMivOLkBf7CmnWi9c5eCtf4VSywCOl6cWU9rg1KV8JFykX4isbFOzNIBZ
lAEfTSTfRhpw86ilK273VeCrSV98x5jQul3UGORIHciiTyHPuQbWkK3rz9CqUosyTh0ti1jTha6G
0vTqDRyozStlUOvUiY9dDSmOwpZbLtJVecmQKfP5VeLhjEfYyTUngwHo7bsEiuBWvLosi90Qbors
G9GKs1jpsE098eJtsz9nT28+ALfTeXe1llx05QRM3GVQMTbEYn9auBWsslfdhoICSjDvm9DYjeUk
32RX7s5768s2WWAQ9ZRKTV2YN0FeT+9xkYAIBNp7Z1IJIbDBH/SEZ4zHmfsMmFf/mrvEPtuWdiEl
ewgH/hsC3XkKuzBcSJuiDy/lsAPzojOGmZz7WjJ88L4Im87ZdJg848gcmhyQDxzmekH0nu7CquKQ
1PmO9N4ItS4XDDV4ooWvSasMXNxOUacUwAp6q/UoEDu0qKVPQbwSMd3fnf7l0oPocEO+LTwnwTVT
1YCeQ8VwKPFtxxM5OdO1yIUpVYdcnJg0uPq1zpekJ/9VdSaX8kYnHW3Z4oNiVfwgWOxvvmYakOdN
V8mQcNB4wJD1JpJT5W7nGHykEmifl9MjZe6o3YS0WiTk6G6nJQ2549RhNyqnSCDM5RKsysPrg+4Y
YsedniqcIyiiDOehXYXBW2pquJ4/QLP03J84cIqpR0UMkySSJVhf0fxb4Dc776t/2n83wLhr267b
4Do7Ch/VHrkuV3X45uzjZ2dqu7GJoyYUlW2tH7FdIDtrCtDXcISGCHAufT+XYEyrxT3uukqElXDG
MRHXDM4JjV6EKVOkdM8C5dXMigazJbclB0/rwFpy7534Z9PSV1rFxLwaVzefnY0s6Nj9zgBTlfDc
W/u/jlfVVG+EB9pcEmGujrll4zH2L06VX5LbjeeuDm67KQS6C9kvrHLQlK6chWW6vygKfKksjeOR
tKli/uVGCMiuyFuSs3l7TZZlFF1M8z6x37Rgs2qu2+B4LXZQDAHE2SJII4vit4u9UFSDoeFtJOAz
YQdP+NxBaqgY702BHzRCYM6oP0GEaVjmUGovuc0UyHMWVnKvXabfshn9kHKIAsmQh16CHE2DIGx5
M8INS8tWW6V8ClB7soYCz/HZMAJIW4Zhs9hBnBeM9y53OXLbMn4rCAT5qWOb2VULy7loIOb/cK8R
T1jAHJevLKTuAjIJghaTF2CX5DQ1KamdnccxnmhrOnUo7N5LwRJacxRZQNHwU7XbgjfyP4G39rzs
8V9PtfyGec7cs9nhZvOP/XPO2jX2eeA0J7hcsBveXp7Mbcl7BeF8irGbPvDhRPfVxf4FsXkQTvgg
EQW5FAuiuqWImB0q0wTijclW13pj3dGOKzYc5OSj9PjKJiPSsR2xWuwQDE2O5hswwtMUiAjnWP+q
OunP2K8eHAiNY4sO2XzwEU60cvj+FZjSfJWOrQXuI8h0KKit3GyOwLC5XYjIAmgMs/IJdE5ZqPc4
ehiFPo5Hg/FirX+FGvMkznHOLK+IKL2zUvenVLPGlhP7uHxGt9j7SE24KxmuFxjdmoIAqQho1sGl
T0kRKix8ZD87gaw1KeN/9pTgBQ9t01ww3QICkGvbfVyLWNSY5GLEW+tV6D+cdS0KOBoZv28Ku0Qn
JkO7stBKHXM7HoLlLfdzyriPkExc69yV49kffpruM+1cC6hyLPIJnl7Y5GD/ZHKlH8wbF3YKJ5Ju
xL6UbclWCl4cssVS89+1C5QSHlWAhmGN3teVbULVyvaP3DVqUEpgUXH1IJPCmFvrRqCfclBpIWv7
f0itJ5kIhkq9J2Yr2jOkt3FKJEh1L2yJmVVe4Eayh5J33uFrv8PUG9UudijTUAWiM2EPcimN5Alm
9xxCUaee6Gn4ob1nCO8h2IDjXZRiIYNv2ZrI1CfaoUSbm1NLW/ddcgOHnU+XVboqutveaTsgqKcs
rnNJueABBBc1kkminj5OE9gNhwJcg2ukIqazyrMSxr/eQYL9kGLJcxYw72apirGDrNW5Enhm9lbe
KRSWwaUHDoX5qvJVzeI5AYO0jUX5cyMLo4Yw/0JwSbhN7uJp0UqrBVC1skJwJ0s25/3N9JysUICK
UHAywkkUu+rvOisw87kXc85cNLKcSDL1qfG55mXF4pz56Ut9KZT6iciFHdUpTSrnl0sQ5bVWf7tO
Yp/3zEL31zaXXAy0LSU2duX+Pf3gidZ0zwqLwkP5ASqBYTMVWHm5NzQQTJXiDBkeR2zUC9j9kteV
Ewxs8w4GZ5Q8b5wshk5YWqxaXhM4bqic7e5Eg3CjPGyrV5s/x9Vqpp3Y1AtTzd75wnnWrmailVnw
hID51+scBm5Z1K5jakkICbTwXxdB8gX0uoEYrTd6k0fLbU+BUCAsvi5evbqbseEMmuOkbqC3wR4o
i48lDf/i67f8zjsAta8zppVWdDGhGNnuU/ewFkUrHXx3B/pettVQZozpiYxB/eDs3SZyYEZmiQLr
IZLntd+2NXIClfw4/wrT+rQkHuoTAf9bxsHi8zJRBm4qah2uDEgLkaYL2oSAuuQgcrFBtfTmWxwF
IqA253sARtSx5Jl4KG2pi16sEtaLqVtN+WEbK0lR2sXd8TlVC0S2VLIIghTJtpa6389ugfHG4Ldq
6UPFwGJw4lj662oxBLmCbSKSMaprlvJHRa/NrMYd2PmPBKbPYI2Y+J+sKPNT6ecX11+fNX6Oigg8
niL637aFCPRSBlsNrfgFddrVKVxW5tbvcvNRIdaT0+wwal9bUDMQUmxokYnAaGLfNR7hn8MebT/l
4ML9WEP0EGEhjRgdUuBvnr/Z6uAwGYWTTuVhBvBiOZIT3Tt7q8k9oNPNsTBQo7IrA5kv2loF3gjB
Mvygj+yN1e/FbCezx/nr6GPFKVIPpnLiVt8jvjdT8VIABaM6RUes5btIhmDal25I7RtEUxbMhGQ5
DVh4P0KLmXG9Xq88kniUbljdINZU1xiW+imsT8jD008JbE5Op/V5YxZjVmKEOwxguqs72HLFh5Sb
vWpXs0auKCNPAzL2lPM95PxwV0lqn9jtJWAy+p0gaQq1kX/aDQ5HotDNTqwyfpQUDJQHo9HDPj66
83uyZIiU4STQONPIZ6lwuL7FBKnOUX4GsZNCdtjTbR/93YwWELWGK16VCGuAImLmnZ/RkQ3apOEs
8wDjl9wNnDpEr15MyG243IBtpbW1ix+wQ8z9HGIT1cs6wEiHWcrWG+PO3+/jkUgn4NLnpPc/zxfA
nRA/1mbzfhBWlaPEGZNdohjtHpuk7jYYknL1nCIWK9wq/cHjXL1N4XxSElFRpucSYxoPqa5xTZhB
hE6SRl6nTau9m321VnH8CYKJaQcl1cqbQLzPoCh1Mtxasjc96rsB4cJ9cACuK1iK9l37Qb35ryV0
EedmFFJvvzcSakaLcMVE9HEGmez9K7bNIPd4lTxDoGwOSvgauJ+tCWLMEoLJ7L1q/dijchrA8CmS
ut8HAwy0muC561OgebRu6Z9Y/Ei0J61ZPsxe5fmOLv8hvHBbacWfCceZtpYJktdxH/lhQYUKaTU0
41GiNwQ08negSOXwvUKRuvv3YfScKs7sUjr6YRQ7zehVGop8M9l2X7zyGLdz5mc8cfv0ji+H7RVS
mGmR9Do1zysTPHo8D7L5O1nn5mKFLNZMsAPRV5t1iROF+jNDtXuKcFfQUSM74Nb6FYrm7ARGhqmy
FpWlx6W/Raawlnootd9RYP5lAEFLMlKww/0yQDHWXtO0zNG3I/EEfqXNYBEmtrJkMHtLq7YIp9PE
IBAz79D7o3ZhdBtN+AExBWcmPp7v4NeWNb0WdOGgVbnwT+/4+hvSSFSaHroBtvAFemV1UMKeIbM4
B/3Juc1tNVUOKcwflD25OwwlqY+kVoamGoR8H2i7c6TAPyFzpnPQv8ynaOgaRzt8aWv0OhMBrOex
qfKj9FjGjRg3x1uQ23zKd4NhW0Wfp1gwIvrctbRDzrPMr4a7m0d/Dj5StrAzn6nt4PW38Sl2wj+V
7jDZJUqKthPZs7PoHE4q20T6YMHNdUCmWD6Z5FLc3GEKgco4W6AOz6mcXk6j3kwzuX6JCDwtJ8dc
EPn2L7EKq6Yx+X/2x+prXErzhBoZ9rv6+1LZ4qxs0LJACFOi3evpliieXkcH/zwq7U9GeAcGWpDM
PfWy/tIy0vwyihNPJM16NlSuFNGz9E9+ztNrOByUTsoGyjbx3DiKH453DOWINf1MJODVq8rSXduJ
xOnCFIGsWD5B/EG9OvTDSr4fLptSA804kNIPs+p0lKdU1mOmQeAVjY6w7iqVE3d/VLtnsEJ6BILZ
FrW9ZY/bi8eH0XhteIzmTbhUV/yN9Dvxcie2lu6dwA+GX5VlMQ7XHpAOJULqEH724yNkBNOSz6VO
cYA3ew+ckcNNNiztU+hCzRb7Q6LcO+p/OkW9qXKqGCD3MF3wf2CBZRWx2fHKQda20EsCXjLFx1sX
8xM6WK/BOi4o2BWEryyd3UbtZ6n2VC9ytzMqex97DQ9N1RtzcwE21VNnCnpPHl396vu0AWUTi3eC
SI5Z6lPQtQliSPMKbHLxwaeI5GtyK7TKNZPYTPh8Tebx+7QPHDqM+IXwmsFYHLPOSzSmOeH+/osQ
0bvOLxdBKtOgVLT94Sn8xH4JwkpjYJUDFAXZZx666pRniTWKkArUPxsUBOKv9UGacs0GnuGJpsOK
Uss3yE+qJ2Kl1yPB3jykRkHFhRfyhLP5Io78b3UV0D6pqyiWDrsLb8K/OvvJd9L9vIaIBL4AD7Ii
zwA+UER23R6FeP9f8WdO+tZWExTOEnz44N4NBUxgmbmGELG1L2I+frwjmYxiZza6ufxcsWZmQuJx
oqQ/JGVbyhj04ShGHFCJQ6w4GvD+WTRSLNcpM2xDCWPTZMQ7vQVAZJ/9AVoUMZ38RIBnqY1dXx4w
CmrRX9GOeJO/Cl9xmsvrHCfSX831pih5GYfWsIB75z85Cyxne04BiFiEJ6qVerE5adN0gSrJk0tE
HTcnGNdv2yFJYbPff7zOWmkO/TbeMLpObvdL7neh9w0yrsL+k06UTlfSHPRje1dHUpCYrMxKSxiw
3/8d7j0iMSwPWTEWNizzDL4/yP0dCELQBf59IFNgvS823TtK+nGkcMH2Sg3jE1J2VlekTkoldUmC
N/TvxvzLb5ta+RX8S8K1tjJE63RXaelmYawc711pkvLjBU7e96zvzOFdxzR5b7hswH2I463C8yoj
8l+3FyYo8XMiSU9gssuKG9/x+caB4JmIPwtgteyuG1eq3Suo2yDvr1IhxV1MfSQFnSrAeHAPetM0
cD7m6g9Szo22/ZKTxT5Mhr0yG8v88fJtTmIEXsaYrM30QxVgE7gZ6P66ap0e0FCOWGLo8vVsP8oK
of/dP+HCeNW+7OLp/N5Lzu+De6PmrRJYfYAkH8Zen57UKfoN6xpTf4VvE66KCToxD92ch6kK7uBO
Vg/C42Wfa/1Wzl+PGW2Mr8g1A2BcxnPXTbdPBaAFO/7bHxf4OKi2kKp7APBAxuQyHjpdHvwZgaZt
o9I4eug/G6MHtLBOW9WEJ5MAoZ7LNbY63nfXnVYoOm5N67RepJ8VTlqGLZ3XOgBwUkXNWKZ+4RFb
vJ32Bipqv+nmHZBPlZ/Yxko3oAMMcaUeAmPpnzz7MwXOLdiOczzsvwEylcCwslWo6AbDvMjbYQYz
9Lz43t8Pq2KU6QBeofvtWu0JXXnly7w1zI3+H8Nm1N83ayezoL/Ner70p4wexv2BdE2vE7kUzlI+
Dkw1iCKD7o6n6imr/Fd3/2S82XTurB0mxQFBf/pHnRJSvp/iHL9MBihkM5TsoYEu33/daApAfFIw
F2DPPQEepo4wIEYE85Cwb5rGfECu4otbwEvkIuEHjezLi5KYnJZ3YLv6hgpZfo8FdE3sWTT2v7l9
yU+5FEaoDfhOwcvXz0AMUymHi68geaPT7WgJ2VEcHDjsdAZJcxEEiidDaiN7DcU/u0X0FLBK5lwa
pR4Hbz0z+kzvfpcT6YGuMT3NH/J0Dw3XLPtavpNydQbg8X/VFMopct9RfIg9mj+ShjYlc5d6Iw9w
ReevgP6XsRN6H/pUS0dx9jGoS2MWQJSql0WLjKY0QuSgqz5DuuP2Gw1+CqzxnnKUClhDQ9Y1jT3H
FZv8Fr0IpeOoyeQAxO9IihxBw6EVEmsAPFEuN5OrpZmrLG/GSKwGkQFMdhDTf33GReJr+m2QUdHo
ISAY9LAQbhy1IMRtV2Q3tnjSqYt0g68JGdQRV5YghhO+3082+3DBXf9mBKcmTwoOfu048XeygoIW
faEpto+zvb/Iu6rtt8AlzVbvkItuYHCd7lh+yIul7vROhtOG+LMf1PjlPoI+w7qDbFMze2qM/XmD
pcQdbPpu+VtmyNOQFEn1HHMxaLa5In9n9YflleanD0+yZ5osRd4lm+LPPUTBa9bmrjMeFW1Rz50l
RSGWmEcSLq5rBUDxLVlF0VJiF0z32JQQo5hjAB9Jd21FP/+SZ9N+yFNTGJ6+QnzdTKSo4FCaxjYx
q0qUoT7O6+XDDH/8NH0qUosN7NCcd0A8amzznLrR7FiTsMJ8tm8CH11k8+Uh5JuQXwOoKZmaTF5B
ak5WbEJx0RQkmWTSFuPW/SyRBkXEGy2CTJ46p3fiUT2VOnWDaQHdluwzXzXQpO0C4OfoQhC8mAlX
JGP/JJuLnkhsmvxPO4HBkgbF3g7P1RyyNHoCPZxxFL2JjNBGqSwlfT9YX2XwHhOSlZ+ac+FLnw5k
vO1Jv4dfQn0eVAIdmjXQdF+IxLuOKIV67Lh6McOZBqxibo7uFrlusr38GJwVuFBP+axIaXfmlIGp
+7iTBsJnBldMhfXTpWJkaqkwW9UUNewF2u2Y4W5pbZyRwLlRflav8jTQ650bacVSJZloxyFgMLA5
0WX4UZ2h+wxdult51uvPw0e0aToYAFskKmgumI4ILVJoijeEgo85sVj2GJi2Lygvf5jabRLmWVzP
AmfQbCnsLMZst/7b8Y7L7VVpyVGcv68UBWNqmNSeUSfeMHDAn/owm3z2x62VPmOdlUEMu6MTfFKe
Ju39A6g1CCqxgr3c/EcLHtw6JgJbl5s0Xv3A0DkG6T+pAOaVkGuEQpY51emAKXiBCG7/MnBKbx84
p/wr5fNVn1Dy1AAxOSU6rAfWYr3icStBbOwsu+Ia4yLvb8gf3KVOxLnKsUcWPfoPFK536qvba8uD
PJbzGDboKAw+IlLOcwZJIdFQWU6n5aqlq2f1h65FsgP+t03J1PulHDotiK9YsfVdmOvY6hUyMKSU
duvnxUp+a4egSEk09LqnQBBrf2PAjXKWJnXCPzVZDGjP0wE58xvvnCOeqAtsC3gmDz+fCXPv2Otr
sq72HWR3+VmDXsyJk9JnkfvTfXZM/abkwsi1hzfRML8eVCbqngEIDdy6zKgXImGQ57wL/UtwCKZd
rKZ6HfUxFnlrPJ6BECkfqSpeUCgGofo0RQfOTFjFCwmEdk9jwRG2GKPAEPr9+m+qYkUsKYo5+YeV
3zByaeLm/PjDEEHT7kIHvrpYXYmVg8o8KknSTiN+N1PwfmhYdr4ecIlXdRJ6jytAZTUjVV4zczWT
21758yac4D4O8iaFSZlPjPq7p0N9f1Wx191WWRswKORJQZD/uiwp0M8alfmC48xb0PuF8l+6RDSl
c9sqN6NJuujETOgOkf1CJenxvT0T4+4Yq6jTGYlN/YetN7+EIkr481iLMQIKhIob41Ie+icCXbCE
2ZuQvaMguNuMh5tiGX7RBI0MRMZIBGZ5FCjOlpFr/XAKIbWu33+D8cXHJckPzvEusy6+QyWh2qc/
hYQNdVIzGTeoVPcPp2m4G/yrnArPRwGUQqSbPAUA+Nc8CcjD1MiJ88TeQanAJKY4LiNEEwAIYQI1
/R6WwR3k+vZhuS1c8qDUG6Vhy1CcHMDkipqyr4+CtIunL6mj/p2dRrtBekw1hKgrFFIW6mxj7Iz4
DAYA2E8W9DPkP3pIflH25lY4MpzDzQkozsmfxlLeFRfSX5kpLvpaRZ/MWp+treYOlCf9IcM1kNZz
9zyN55SAGjZLcKBQJTooqxAT3domqr9NfDqbAYIyxHRUd1ImkvRGTBZLADBj7aoGkAhlAUnQgagr
D8yJPXHnen+ozIHHSsF3S/p6/4TzrU5xSicV6kwyQDk9dhxVlhlpW0GjyHBXWRJ53E6jTDpVC7IT
OCGoTGULZ3pnqbh4xVNbK2CnVXAFG7NMZ4yrbsdP96wfLVr121iJS+PF76H4oydapp8P1ldZZRqS
4DFc/J2JbD91xyaJC9wblfdjHOGDWVJlt9QIOY1czKOfZCL/axP4GpUDKy1f53D8r6WGdnRvm5EV
Jxw782Leo1NuhZUbF3LVWMBnq7mRXcvoUEv2v4dsTvJl3WMo4c4kAx8TcoqNpXJemvt57/eSHtZn
L6VsM63h09lDqqZ/GOs6BCIYve2/G8lOVcUybCLXlJWzTKhdstMDeYbBTQ2EycTHqwtr4gZL2Xrd
c54XoKb63zAPRHa+n1nsqmDgONPPOeO5ijYLaIJkYFBAauBg89ihixCzDvHAmJnBiEvA9TUwThne
Sz2hkRXmaIiBtB9rZkBliTXW+Xoeq4C9o8lkLYPyv7cXV+ZJHWU28sVMzI4XKkTvTesqd+KOFPuO
ALSYj47S95R8uiyRVtjIxXo0V9Y4Lv14qK2tOvw7Dxvwe6zFWvs64UlyVCXt27QxIliuJYEgfd4t
9twKrRsxyo79YFVumHxWah3m6qdEbwXwjD0AjWyvYBeTVrmBJFQMQi3Ln2u7pyQ1lwoSR11koaYt
v7XdYK+dcOfH1JpznK1zLODOwWCmZtZDI95Q0XerolS4gcqkl3K9Mbw/Xn289nlwM4PqVzzxdQlz
vADOaQA0t5dzsEfz7bezgljNUmKEX6BifxzUNKRWah8njOOlNJ/YtacToLH1eppAXPPmACTDAVqs
XKkehwizobh2KJ2TOyKFjyJp/ywjw6QIeyf34eFkRFGmlzZLMtbOB2edpfUqdf0CSX3pN4TgbmYm
KcydIIzJbN2XTIlk67EVkDPQFqEdJ8v7YNJhPDGTq4rq+chy8FbOENZBBCzvQLKF5GdVPlAoN4YR
PhthrKRsoYgA1i6rSqshMDm7B2y2yz2My1EzQIFMxGUITOAyiOyUM3DGUPmJhYQQcmFJliYhsmT+
7NhqfrNgsF6tEBwa2glUHOda56R1daoQ2WY4nWF97AuduWiA2pCzBBtHgVflVAbBtYk/SVNEIJ6K
90/mfNwT6JCVwpDFnmJI1mYsFo0rJL0CmuuKoKhBruH1lsyiZrobDRahgQzn2eSKPdRAuEBrSpxp
7s0H25+nkVLIz3UyaAN2pCRCl3k8fVK7ARnW2kzlABfC8wLqQv6AAlrcbj9WzI2JoiMd557uAp4x
fnSGp67+wZJ1crKuQ921MEEqWfTveDvSLV3YZ3nO6XhOyzkIA02+Al3sJY1iJ1MWuy1vmOAF8QLa
KCKDIh/M96dsHtXCMSIxgcUeD1P+WPPLGldyYalJ4vSpz3hkbmSvL0kwppcyarO8TAk9ijmdal/t
w1NT6tUh3ZZaEHYcf7ODSPsN8SO0znH7isadIHOYyuKt+69ntm/fc8Q7GUFoWDfAaZ7hHvJxs9a/
8+ZzvDplEBDbkTWegc4IYoVuzePznzf9jWJeFaS1hDynGSJNMnqWfJRQVTJ/9Q6SYOWLXKB1eq/Q
FKHc+vcfBZ2FhUGvUKEytYX5O0HBbbgkBD6SCfa0h63SyBMEJvREak2maT+6z+/bTqy3Jw1j2dy6
98ZOgo35Mh9j0dPZiud5HXU01OO02MSUoJEd9Fk3nmvHni8yNQShJlmfePZj3a3hxbKzfxAVZOC0
8+5ejxMuK0qovxHds90kqexAM4M4k+mZRPoYRKgZLa8j8QiuUQsY7JzjR6CgAMuY2M8/05+WmkLt
1dZ1liCOL6OaHKgwq9aki7wi+/eX2KEAHnIXY9lY8s7gtYOkrjlcRDGzJVJTJrkNI/TH5m+JgL+Y
xCr+NcHEH2rtl3EpBJtBZWW7lPFaSF0PjREOKVocPcjQa9BN4qV7DvvqC9DakRLe7Y1QexZ15MdT
Cf2TI2FOhSddDCddQVTsWMMjbjS8YyV6QrGMdTLmM/oLYOq7/xqG0ErJNW6dISFoXsVOpXEU7YOf
ZWd/qioPWlT9giFyCz9sWYPdJexf0AKNv+8C/1tDxf7hKfNFfmKIA+HdXNsVJAEwYQ6DDkKhVOjm
GaFp9yGHfMjitoqFDpJbaJdiTBukqdU6Yo3E5Fti1lXUXiANFHqn4R7l7a3snJ8UaMmJ4Vvcyf/a
1pakv0LUiVeSiJprayXNDuIAWZsUtwxI64o5inpU/vw9rz1WYkOTvRX6V94cK3CL0SoqcwKjceXL
vC133nld7BuH1aMmcbTUxJm23P3SJzT8NzqgeRk9meVo4jTx9tMn3pBGdQKXCVOYgmPU4PpYugB7
MHAksD+BbzxTI2DvuuwpA8E9NMkzw4qHYynsfr0BNlRpdUTn24NduCq4B07rO8UtYdvUy+xe5Tlg
mAzVR/8WcxRFOLM1b3ulp9Jwb25DWr1JeNyqv6S3pITc8fWOOExBgH36aUhtNKuYl923mCiLo9am
QIwoe79jSuuZgUbcGcgLp/PPGAG7BBJeLYt9ul0MpwP6fEIt6xXgZ0KLydWI/05sME+ir0Wkozta
v6ycpYA/EwC23PID6g4KrBSUGMc3sqDEPfLpfvnEJvBAio5//GEguP0r3a8NLu8piVDrzYk6Vl5p
EohsmKFz+e2QoUmIG33uG0k7o53NMNaVhsfvtnYVrK2vBpIJuE1B9Y0AUeD1rscLUq5tf3LTRWLZ
7QZxuvPyUkNGBzpLsWHF5h6/fQVZO5v3CbgTdVM4wGSjmDd/oBF22QaUwxPdMDNUk5aBkT4Wea7X
yzDOXFX4XWBkJNRGgOi0DADlmlXUY9fjnOHLKcoi6zaWnBxni3T3A8YTLDSlkVJ3ZB2kz7US/sIS
dj7Ko+8ql8ELKpBFDMn57wT2E93Tsxob2cUNsX51qG6ZPscRAIRJ/XEn1QOnXg37qaUZATT3VJ2e
LCg7QitwXtcVoJMxk3zG2bkQekK+VToyDXKVVpi8hrC4jS3RY+2RypH0HlAEJ0ZKpM7htlFZxEau
3oIFIzSVHrYXg9dqfAgwySJe/7zTv2kBXBqDCS9F7lokBpK53dRWgfJL8K85NA3I/LFk6IZuIbxX
7PsXIdUkiFqzhD7iFinKM+6v+QmO4k/8aALzN1U2l3Ohw/2RXLDWL66W6RpeZ3ZxslevQxYtPZZa
3/ciXi4Ql+PDsMyMnnUxS/FQEQ1fizyuIwUcJlp64QYwa+QH/CZplNMQHdmZvS8ZHu7zRO4I81y8
4aqTxQm1STRIcJUfh+zuUJ6eyj2+rIoEEPqVc57W/J3GOuNn8hss2ubpeWzYDBmpSMlemGeveni9
y4v0mH4UCvont0tO4M6ZDib+bbPALxK3NezrAzQCtVJ98wZ8SPUIdwV3BB/EfrZk8sn7ztfwJILl
KlbR8OhnHTTUP7LCkpmr4CrHj7Hb7rqhM7FqiYOZ57uttQme9XXmrd5xBCnnYCloYDgQm/N6rRC/
eu0eWodP1RKQNsXfBfVc5EgTgnzHX0ySLVdY/BXQqEKa5Un2fs/TZhmsJkMSrk1ONOIH4YvY5+Jh
v6xJK8kSRNlv63F3IJDObPsvy4Iizlo+kchHBwIhChURkMSXXUV0NhxEmOzwyPp8MEGrGanxjaLU
ePlsLA0VvlvB/4EuJVHeaCwSijhU7esQY116kevRyIWKCwHtJpcKHSjmHIghM1YtQS35kjINOHSi
pD4HJcRyPOsdtALG9Daakp2HV37b5HDhfAjIDody8kghyg7aGunUbqC7wNYFmwwLN6Qct8IzQDY4
5i4UqOdUOJRxyIWcQIiby6HihzgL1D4LEgRXEyqCyMLAKXnuyZBSTH3w3dc6/ghSMemS5xC6eeyQ
I+FgTXPi8REHcfbxPHbFDUyZPMLvkgZoK+BxDbgZbPfBDCkvp5W1h/Bz31SHzvPSLjAWXdFZJ9Sf
eDS/nQC8eMkOTDLQHF2EXhdkBHI7gqVMYudhm6mnKMwx6Xr6GgwTQGy/28YhJrA6svrQlsdtbqf6
IERP1JxWKIMpSYujyKHKn6hCkmc+QQgjVWhsaEKbs/ZsNcJIANqp/C0+uaLO43eybHaI17EbK2MO
sHEDxn+Es3ejtIkAdrDmUKAcOlYeEOtzNqlvHLpyjxtAH1rwORM/DIm+LKXw9f/7Jii2CNdaUItS
0MaokTSsYez4cE1ADpiDrXmmLgu6T6Muttd7/FGhbwKW2TIpdHe6/dqV331BwyaHD2DF58WBr6ro
Bcl2FOcI4CNUgdqDlk+Rhp4pJ0KXhb2ddfkeqX1SC/F3g+XqO7u1QCbe8yuayUuEwrOOe1RMWsYV
Sq4/jWAhK3yhDY0FGTIf83n6V8NjG0ktIsmSRzhdS5NiLe+fmkxLKJVnQZTHxsL3UQAPNYZDHvbp
0Nj/7ucB9t+IrgS6ZmefvV4c7HdxcOJk0Fekcezh965f0xb6a0BlRIPVbSliz/JLEOROrdhismik
4uxqSkVpqUXn1eqj8tRxPViJWwSA/17JLd8v8bXkAqJPytToY7ZpYgqatriXfoRhPOKe2vBXZ1wW
hX6QSmvU173lLfXiPeV83UhWcYzy3mR2Q5cH394N502671bM2YLEw+yqdVnIoO5xslF4vgqfozaZ
Gq3WypMrzOo46UJS7b/ZW4r17dDAVpZTFYXo9/D1aFIjH2U9NbktyGFVTh5dmDXMpN08V1N6Fl9h
040qEK8FKsOVAgbfRD6rVo36vfCbUb0g+VPmpIMcQn2Ak35WNxryupDkencBEtTyKLfG6XHtPBFR
cevOoRVh3PANQHey0FP+qvkz/t1UXV6IwZcYUClTM61YHRlkm94xLwORdKVSIHPjqbWMXsc+yCco
rFefEpxeHMTrJGPNoKbS6WDQ2l1CzB+dMrZAdlFeoMZ4huI02/zGcR+Zod40wvuAHLPofabKAtMB
jEIfYs0Eoj00ScpKq4Y1UU1b5RoFVyMYh5OZ5KFk6fnjSZwaGIi0a/U7FrCgmaBbe32gg1WpCKUo
VwlZ0uD+JQcgSYkiSKM+RNZNjy1xZ5MpYU3JCgzVSkaEBBNQQb2hubKHx7/6prudZUcdtdU1MXHb
bBgCqyMAkeRm2rv7rLwmMtS0dX/VjYH9m4+hNEJabDXjwZq/kWNkfBTEFpKZoRBdormOgPscUHxo
itmFEFCtv3KD7vcnZNK8TdNc2e4P1fJwe6uLpqzpCII+bMoHowVVKvhrEYNM67Nq4gSwnZbT0fbN
l6BzNH7OLKypB/jC9Ra5U7Sj3JA24Hxc+rLMhzKy851nUqMHjvAccPDxUN4YEPlCfizVjkaczClF
chIjQ/CaN4hYDZi/JqKRN2TIEi+R7MqmO852VpjvKdZul8rVkqLQSDpcrvxiGR9sLoSxyuzGGaRR
R6Om5WkmEMjPMsQvN9J+VNbJJVgPi5p8exqkMSXXmAmBXtID6mGQuUuVc5KWu4av0Vnn9Vm37OKw
mF5n91EtcsZfA50JnMtztnvOLblXfyrOxjjbDd/+yDa73bsyfUM2hY9ueZoGfTmNaz3Zj39k/Zvj
/y6oeamMimr0goInwmZrAGOMQSPEHpV8ipUESlZi+5yFbOLa08JQ3Dwj033ywsl4AEEj5gzSdyl4
StnqIAeB/mxPdwn2R1LQEGlRJwtsGspzhaI0tMNU9bdGz9uoA6vf7u56RawX2V7u+kHnUvn01UY9
VnK0PwOvkESVTcde8bV3dLt5TJKPgmvyeapBiGHI5FCpmzkdgZDmRLKfVonuCVWls2GV1zph/nCF
HB5sGQgp03VCx69XEmjxpmUBXE8yHmahDvFCgisoaX0qiCrAzlpl1gtDBTMSf/3Z2jOIQvtKuVzJ
Ei8WE8IQdn5OwXCC9NPQLtIdIzK7/17W5USe3HSWWX7DptuubtVET8LIT5M/gAOpz0hCsFHzmB+8
lTG2kRAf0btC+f4sVkrvyLZM58Xta8TV/8reN7zasvixsUh870JM+TCivOuIf2DO6o1rUbgVfUyr
BZKG0C71zJ/2f9P7U1oIO1u6TdpyUN7D9G3uMFz+62d3cPhe+7RK+BDA+yYU+J3SxDjDKbyBvCnD
ETj8spDM0cC/RX7DNO9JhW7EjHkejKCRg4GpzvZk+ygSyX+ZgN5fshNjDoQw61RENfaBaaIZ+lGw
+yaPRYjCRqFDRXOo7wLflLiAYt15MJLELYSJU1d6os1Ty/UbzonP66ScuZXEwBn5hxs9m6zMF708
JnwPEvyHDCn4DJphRNfd1/Kb8maMAF/BOrDAFzkR+BY1yPLj62yuAIwfTj1tg5uHnp6iwB+36rZX
Ih2JNT+QDe147cxUeJnwH48V8RqHs0787zdDCMo0eposME0Gvej8XFpsfBEvtaHYU24UQf2rmwAO
hMDg39ojVU5wz29KgMenzfFiRJOx42QOBgUFUlSrkoHyPeR0mZkTxJpNmjbqi6CudfqEBh/78MmT
MVVLiApDijmRiUgAw2MFJm5O5bltn7QNQsJWFRm1rSOJg+4TRVZzy5dDFs3ABvda/yrJH/tD7RTt
pUAVPZ+kmO7zy4CwLtXylozXqkpbRLjpzHAT4ZUo71Q6X3maTOYAN+vVQcBMyjYZa8yzXphXbkZa
Eg00lZxFkyQhPTyYP5IxnFXReqjuhfu7UwvoUmGVu5fIe3P89OD8u+G0WHj31IkRhRIBpb/c6FD/
tHdTByKJ8+kk+VG6eNgcEZhrdg2/42M54QKJpZJiQb+shfQ+7Tsb3d6gSO+ErHsDNrGnXy0I0SXk
Yr3EGP1yKLHZ1T9OV10y+KDA13ldJkDKCo9iYjlzRXsIMJTMvqo6ZhjrkYJvyXTkFKOwlKi//0Vf
YH1CRJN5pjlkMml8R6EBUXZMmimbURvZWhisFOn+mILoCdm46X4LGyk130CmAlErjewjflc+lbny
fQWv5AeSv8xfATXbfEnhBJ0aLmtc4UuxKsZgeUAacJ5jEVSW7ploy1OBTD2m3o6nWPZ1zw2PMdCe
DNfyotx9XJxNQ44LdZ4HsGbwC7oVeFNDvOURTcNkbrw9oKqviPPxnja+/SY24RXQx97NQGFzUJbV
ZTQjGxj9CLF9omLKg7J0TnMd0lCyGVUjpHNA0pLIxl5cxtoaGwckUSYrfihMVGenpjUDQosQeP8T
GGF6uxLfcqlEsdLnTm4HspKpWolBIGgVQPapLlOqCGF71w3aBVkdJC7pDYzd5vtwO2opqRfWLg5y
hP1vBTjAuID3MQo3JUBNn35ExtgZGD4us1XHj9VIfDaksYWOC9KjEX4uydqH1SaEimVPCfm2L3gN
ZIcxfQX8h/9Bm7T7LD+SM5RFzoCCQjXrQTix5O58P3Ms1aJ82nB+66PQaW0i2nPtyLhGkUD/XMsJ
hLO9tmddwLG09UZywHhhJrfJIlfqV3JkIYasjW5pn6MH0Kvmb8u1RY4Bg6GBodwuYFF6XIURgqm1
kJIc6zCRrxgRAiD72exrQPpCWpq59fUcuiOvDc5RsWvZG41wPHXTI45dG7ixt4oEt8ZuFrKy58g/
YztDQNzu7mCHjzUI0SK+ZlVG/L1MNygUTMaYuGz18WpOO7ZY+KXmhEYXmwvY1bv+A52aoGlEyB4Q
6GPfMfRvZEMivqCHZRuwPRq+6LcyWbNmTPx2rebS7dZMM97tVHrX5zyf7ZrZ36vx21sj7bBRN0UR
0n02/zM1F0KT1mpr3nZ7D7YWEzYL/d/bDYOvxC9P38b1p4TZSxi/PQQxQRvrmJ3qMvs/WjBByYAG
Ks0rI8Euwq/8bP6D5SVieAc4o8xulcYA6WjGmbZRm5/E77ews9XT+ptakvhGf5olUrbEe6jFFMLe
r0FuUV3X62dBhUNGosp2/dBzvj6JmdJBEfJCo+ZeTakTYzukG6I2jECVoVbLt6KyfOYK1sEkNYjy
+DidIfn/djO+hkq43gxRDTRsasbKXH8qP+H26m/ZjbhKPRZzyi2H8e8F3Fz68Uumi+teka1Zozh0
+S0enpchK6EsbQqrKxuD4cSFczqJ1ydePyW3JE/3qU9VguHC4MsLMu4fGG3wM61Npbqa/cjLFk/c
pcrQ9AVUa6Pj5efxE9OZnF0Cd9YHqdej20FALv9dbypPFXWZGnb2uRNt/h3EPJ5NZxKgNU/KhttB
v/TbVJfi4g0z7JnANHhXGDHrRkhh+9jtgN75vhhKdUNUscUzK9ys5Gxj3IhRRReadbGZhXuzKJEm
7cL9uNewcUnYFRL65P7OlUoBPsmnM6ntkVcB4OnW05vcl5A4cxyJ8uCRwQ2UNr+eSxDlv8jfZ9FA
mfV/zASSCSwZ7vJlgrMJlrjcELwA910G/YcvRFMieZu7fO8d7K74wW/ljs237fbJU9oLfSlG/7NK
swBD/14cXqVqCU1tqicg6eHhS494/8E6n/lRlmaPs24okCY9EAUl309SnHfDM8V1XCowttHk/K6S
KtdkPFfSUCAcTMTwtL03Ns4J9PJigZ4PxymIf1C7igEWNY/swPehHdC3YhIjbiHu2dB6wPMhDRjj
4nT7tMUF2bojF5wsrHxy3OyglPdLhIiI7UxaMT6xB301y1SOP1Gvo2tJQROlQThZ36/ZWr7hob/W
nLMDQ2zHQ8vy0gKHB8NO5U1ZSFvw0lesZbkN97WkEQKPUqTWiNre3n44j8T9Ucv7FOWHhaIcx5pW
H4AgVldBt2CyfUki1bHa0hXMm5gVa0pp5pXRHmVk+lw4AaZ4lQzW6JruyGxuEdXi6/d6kTyFDx01
CntwhBsdMXVqBKUqxobWi+tMmQbrcAgOwZL4xceuxH6nm80JLSxQ3icdUxWPk7Hvho0eEKicz0Rm
FnD8OUBNnaHgI5ZwMgXLdPU+uwNOoa9YoDvyIbinIwkkEGR8OPBaZ1lPCrvgc9XW3xKgLVvtU7o/
Dsd8cwvcNVh8lkQ/evwbRQ7IkuWbvaOV0TklGlu1v7BrRS9HmyYOOCTO4YU2xranxRLedOUQr3/e
5tAi+VYjG+J5vOIle+5e9SxDxS/sKlox9bcgwzgJshwPeUVpyJt7xRmQfWdzzcaoa+9hS/jUPmT/
Xv+MPGWUN4EEGpdNnIRB43QPVKS5g2wAbhhw6tnuM044gcYmgg5/kXyBgprE+7XlNAfU/Y8MAK8z
vYU+SiBDrpC7EZD98Jy30JtgkvQTh6urLKqjvB6GYIiz4nqQWnjkz1KJCGIAisx6qtP0ygWJgy98
NmsmAWYO4pP+C/7H1UV2ivMyXZHtSQiVs8/5si1Kcff5m73ndX+vhrOKQwfakhcl9AfQ2w/gzHu9
A+Dcs7KxgDBcpkC/XmwPiyf4RHo31GmWOxqHCDGhdfrrR8NWaKOxDIi6RFYUb7sthQhjcIKTFhdL
3QBrVf/GdLUdi0yczRKlC/iWmq4VJlT6zbDJaME/M65lI06Z//BGlNkJ6++rIlLyinjEZKLcRYHY
xmCliGepdgtpyst/9rMwFTHjHoTgkX4ZgRK9gywdiz/gxCsiqmONnFsif5oHZKb9l4erH2/ALG7y
bJ2pL17BeYNAfAk3D8olHje7hKZJimZyg2Q62QkfapUK98mhiBaDA3ntCiAcnBj7fimWV7mKVyzY
9MDtUbrfIa0HbZpx8lxzkuERQ1fCZdElhuMgnxu0NqWU6UuMXzSy4DLeqV3quu6w54jgL+NuxjVN
0RGn+ITVsW0H6CMpfV4v1BP+VjfeVpjjPPShQROc7/jKBDVql5FtLtCIIT0EdF/BhmzV6ohcGWmC
0cCnRpBBGwPwP1KCmN1T+v3h2qeOKOAViWDjdU+X033ENhdI108UCxRBGkaFYk2TBTmRAO+6AcJs
Kjqaj4PSD2VBq9GmdhGDFmKwFg8rYNCaVB2tYNBDDBfIv1iXJN4hUbvN/euTH1MdsvumgGiwq+Hj
aHCcAZX9lNyTbLGeFqQYCRfQwedR0eyb55A9kq/s9VfIoH4FsgTXLiJb9/cVfFsb5OxnDAAaYvzr
+d0oyf03hk/AD1YpU8E7noi2J/nM6uvpOKnuL1evXO2+rQjjrXvW7i0ZTLH6WT/X97CN1g0MG0Md
O9YH+zDu95q0fMRYciRTnVK80RH8umDy9Pgzf8ePMptulolZe8UYbTROrP9q9wM0X3eGBt7y542Y
Tev9Tx1f19BSJ0o5CNV1uYBQ8HHPr4dUG3ehB7RmqVfsbc7DPmkIZ+94zNpPCriiCCK/2W9hFs6d
LcazKtizofHNfEVoWZNbfkS6WKZF98MJ8JAOMXMrFq7t23Vlg/i3Jyf6Lp1meIcE4OcCThoYMcFY
NYhUppceKEakWuci8EkeO9W7+QiKTvmx3ZVkSVcjBOvbAJcIX5soSgUs+IU6Y88nz+4o26+BcHLp
8rrzqyutqY9nAtoV3zI4J7JS4bhZkRszm40OY4/abOmmf4AXcuNln8PwZg23JrBUzurgQHUiZk+F
EyEBbnMIhAuGPCI1djXJVpS5j+b0QsTLMMIfYc10/cHi6jX+z5XK9VQqU/ub0m4w5RhGv9bSmrr6
e2xSNOnhPhW6iFPU7eUPxanb5nQ57NcmIS9EKviljXhygqQYzARRrXiYoZqsE8AWYPx8u++E3kjx
cktvajQRfidxG5KjuWfzoE7hy+aTU2WvDRXnr2NUdGL/I9gXnZJpykDq/LRB+heBeP1m6FR8t8Vw
JLMyznxDZPB5wvcbuplUyWFmO8eKajCun7HsKlBC/EsBQSnSzYa+uf+HZfSaB/wuUt11xL4VS0Rf
/oZJmFUwYx5hVTh/AzF8YDQtnoNCsxJMhoaO49hbQipILKbKnNavRC3GU6h0aAlCJkBzOAPN/h8S
DZZGfu+PV1OHrKKamPyk3Q1gXt2OTtsQF9ygS3YuH4WqV4KpZCdS6TVU21S00Ws8fgNgjLsXaQWB
XIdg7ZOr97nCxFAE4xCACnkUdl9digigGbfzj/sjyULzLgjivHqPUHFftO2OzfE1nF+PSClxFJWk
7vkwI8mJvjibO6Vy3YPsWg8oN/MRGi9fdJfHvHvwiEW7FfV4ucQLzw1/E0o3ZLdhoTKyizj/ojYt
cKO+UKMjx9IRF7SHVIkMohqo0OGQdmCU0GqZyNM1MUj/DyschaMRCi5LEG4A1QF9DpcG4wi13hQ7
7FvoKn8YlznpVvvmvt9oGZVfauyDH1ZSO+ITTag9ndoaKVXa0hfrW3fJNr9eOcI0OtzH4iowib25
vL0cn7Rf5S7FAmKonQhhjGI6ROp9s+qewM2GI1+I/AcFu71xH09NHbAwFu0Ck48MXAUSvQCFleCX
xRiw6Rqj8H02ncM8MGAEzSM6U2xVdVa2t2t23tzh1PRlp5/2J7cZVeppj6AdeN7pJEuOe5fhDTDA
vjXwKx3h+DzyPdeh/H0GaPQd1ArADBvauza01d6aMeWZJi7u4zHbl1oxYpop/qg8VfnUWwTg1zq9
yY72nREhIVgk5b36j/kpWasAqXrMkNxOyYdR1imgJc/fh/UrA+rohDaY31u41agOHTcLtkx0f9Qp
X95MWmDzskbMD6IAWV3oYWv5/BE1P86+RLwtQFDjeI6x5DB/ywAPA6lZ6mWzPP7buq3z+TbsdTcH
n5M8btwdIKPaXHSkYqg+ZMFeKLdy4GWBhXe3oMYdS8h+guYDdT6RbEAfJXG4X4BjfrJZ5NQFi5EQ
9hpV1OoAH7fmdtBeGm4Ec3sqyKPMdx0gJYaAaSoFfQdJ3avonyyYCJLeddrOovyS9nyN1c8zpt9M
XNNDoIOOqq6AImNBsaHUeC7CbFBZGHHUM+XaIAnyAaLNlaob6LeJAGFf4sxMyH3bUEYzXBxPa4TO
ZkyRLRXCqR/Hup5RsUIg4MOvqgK+NGg58Qwsiz50nmz1FjxrerPk6Mi6n1lmkvcoYXvo4D0H0Gg2
9VtSbSStVYODcRGLzjg3+ZHhox1QjNYitigGXo3+laxdJ3t7ZyNRM01bbbzv6/9bWe4+SWlOoVUk
E/Y00a5u84BvreNOyJHODJI1JilMjly49Geyzoe1wE2b3DHl+wbSCNigh754B5zaH0gLa0EQxQ9Q
wz3b+vWcV5oM8D3C2UHBa5DSJtfa1i9ILTYjA5msnM2ZPYBauFOswWPThaKV7JfwrcmnWwCxVG8y
l7rb3YXJdOIzKZkieS07V35wpssfPTQ1a0yaVwkzdOuEjFjOXrQ7yguMfiqKJfoP33uAPXcTRkxN
9wbT85kJYTmmb65axV2Bghr7+bpwhhRZMhye+Z2wQJ9fpUvF3Ua22swoGFPOqg5UqAk2gbmpYXnb
LLPEBvziYolyd80WPt57LX+ychOf9fYoyVmMS1pzTQYSBL1d2Nw1nbbsa9KJEhlfHLxYvMMTOpBR
AELlspTzDsSpLb8nLDN0tMbPcFSIxz2K0jKyDuiIUikFRNh+MrPTU3tTFbeSfP3hjEP4kA9nfht7
5R3KGcar/v/jnm5wfhz1/cR7B24aisxpWSDzjD1x+vT5+W9tUtUId4q7jY+1qy50xfxs1lF7hkHk
JgXbn47n8Gf52eQkXJlWCtoUHF9XPqxrsyYW/chQvb7ctDvrY0u3puFgC/QsC+sCN9E+YipDrwEq
BHqTE2ZAtLDrXn0KR69spglk30yrJ7h0Y8B8RevB2mfUEXT11ts3EZ2rTIAru6/RVEWW9V+2moID
CzBjaAkEO2z8Gry0IiOEGLr4toyhBoQcAPJsEsr6aXgd3SCfF/eNs67jhmBLYwuYQ/p1ImthfboZ
W4z/GhypbCDEtrRIzcBUsxsWp6cmK0I1pxf00zZbkC071GHryiPez2GHyg5xSVOPe7qo+imY9FZB
zpARCws1AaIJ3/kWv4B/A+x50k7d3kDTIsIvQaDHPomjToTib8gvQ5/ORLfRFfmycLIE8HVMSE0j
kI5m8WGrbbcwppPGkVmeCLJ/qnoOhXC5tYH0ykfpE4p+cGQ26Ms40KtrN6sK1lADAcD8JNl427zZ
6gw9pOJvPId8Qt0YhIUAG0GQ/2R6dKTK0eMBWiWms6tcBCgrKQMwGEWJP+YbEjTKsXjDft5L9qxs
48R226O4uIWyskVEoKEqxDofMDreVUgsIhsFWOs8Ugzrp99TKgfafN8TIImLhar3cZmZeGMWyyZx
1j3yZFN4I8vCtDkP4eeEZlo2thoSNGw0qmru6Icb0PVuJd21a9d/N2kL1yJQDQGrgHIfhtOCnEXA
i/sJId4mqQHJuss8oBgnL1jdPlBcTSq1Fs4b1mzdjjH5dcVL4Ewl7YG1cF1C3Lj8M+zVKCjro1Th
MjJecRuoKDLogvvtqlcJpns4hVe22v7eoxAge+i9dix2UoWSjtEcASvHSDVsPCsW7HgHWjPqlqEH
jNCpHtI6XlyvkOPyy1P1CbHoBQzLaiW9E8cK6kGFpFxvWs9Zk8ai9hyT8m4e973qRoO5lG19GK6M
ntOs4U+R+k0PBmKMFJ8OtnTVfkU8TqeDmHq8mmQPXLnpfSeDLP/qKh0QEE4lm6lOYtw5oPp8EVIr
LQj+zKOSORAR4S2baBDi2lTQUnCs6b2V34Jmu5s6qP39yAWHTffqb+DajJcF7S8ZSOAPZcFV4lzn
LLHnVsQbilKiIDIrIqK5urz3nDcNZ1PBN5hb906sRNoL4D/nbhPWe+dvB2SMKR557cZa431WyjrP
esxrb//p6rTjuzGonnRKqYHWnDwCOAST1rA1qVlAgebgxb8RTibMscvDo8P2gsRNoo7zhmD9Z7u0
S3PjA50zyNqMxXbS8jU4yWmAHAU6nt3tJAlzqH9uudGXj+9Y7VW3ks1a+BLTucNdCEd4VccJpZYG
PFNhyA1xwPu8K4wiYjh11Eq+6i4l1HG11YCGTj38TdZPz0L6l6UgINIg08W98QMRePGgmmPnFI3c
qSK44m2DL6oMzXURnEs1JAt6QpM3bMgRbdFOy7o2sBTx/blpdBgxEGxP4OdEFH6jRRw7y8cdGzes
eLL2Ttphw2B4xRsNDph9KLxWbiYriBL+Cnqxn7+5SAXpbNQDp4SO3vtV7ILmqa1BwdBRpH/lTG3f
y0B9wrtYnKFni1Q+k1jWxnVZXslEMQn4P6BU5x9bu3V6k0lH7NpdES+7cC69vMADZzDTeFFBr6Dv
X61DSD4g6oqNrs0pPxlEoeUCK/g5SzGaI3YCD+9p6NSUmnA7X1ldTMt607j+bEtrvXeNicqCHLjN
8c2JVFg1i+bhufoinv7tLErUdGyrUZQktUT/m7Pe0xO/NZear8M5ZFjjOBA45XVI//9TVZZ6eHOm
e58+Hx8lQ7nqVn6+6MEALFiX4Ht7NaPBtso1TnvfOcQS9JwigqEcY8oOtAfrv1Wq20DFJMG3JvXB
gZ76gq1RzIcZUQldldaiyP6DH4BnEhpKBFieg4c4UZK+CLKWkyx6T3Pepn5FO2Th7pRZVzf++hht
Fs5W5v+BogptwegEz7RF9ZpJqhaHsaeLaCgzxOu8OS018N9XMjv+2XImS92LwhvYvmQX7phjNHl1
+oNjXI0XRNrfohWc/X99MfG2+8+puZFIzLIi2deGj0MRC6YdUg/cfINlIeUgAijl+mbHgC4tDtUf
tjyd6y1SgnFJhS24C3GL25lruJ1GMNB5yYDMYKlA872bJL4E96wsHr8OmUpNWqBwlRLtLiJJ5XqV
0CiTgxN42K6F+h5/D7fv3QQViE8nF82g04dVI1YUHbeEnvacx/pZfFakz0LU3YMLFEfDbKcUlUop
UlhD5TAowoXHTZnJrBj+yOb40zxFqCFHHjJ11+bMarAPsChW76MD71ayWqX0uHXWRiuJMXExxJ++
EVXXblFDS9uvISwk0Y0sGxjq+64yUWIvV6JBeUU1v2rfo6/99zF3lAPtgHoERD0jql7LYZUQFVnx
Ua6porLGsmLWp7N42aJkvMjbtV1VsSTT0t8wMb+jHlxhp8Y+FWKOGNd8fdhh0xk3EWWgH1QKDH1L
/HZ5AXFVddfL+ByFVqqL66i3T8gmBSfKqUMSs+Lm3Bsv6CRgM7BICoCyTQ60jXNQCbdx5WadzWwf
0OWCzdfTNj5FIEaacayqJPQO+eLmNPegynsu4rH+A1PwiWhL+Wt+3iycewwppbQzwpAxe1mJnqcq
6atgyww0IBdfHpoXyjmA8xT0adF1ceQUiBjH0nYf85Hi5wq5BnJy6UoccJ9ah24vRgLY3x5A/2N6
T0uVvLnUNS7/JtJf85dcysFA6E3GsbpVPxEYLsoOU9uzQOgsyq8+W8Io1c4/zF0qapXAR6X/q3aY
wi31kU3xCqnAGnnWGNfn2mgIg6LVi+fHSJ+GeX+mV48mdwK87TZvsz6gPaoEVbbJReQDUZtVuu6T
ccBykqtxI4q0iiTjqM/VO/2SyfLNYD2MfZXak5lTKv/2XHhr01L0ZA9CtkCpb0hLuotgmDxFEM1L
4yorCQOOE3NCw7+JIEmQAHZbyKrlp4DFsQJ+TFGgTBpKZ1uRbdLSh1FQRdV2vmfuZTic1XRTsQVF
5JtpBc5xlyt647lkbFvd/WuNhfPe23vwj7DvwcTugmLt5chffeJopy/NTFoyNCF/E78r1kWOvamW
q3WEgfMVdjCBst/aDPZBx0uoH7bU5cL5Ki/LZtP0/BU2skyKBa1WZvbNSzmXIlebjOS2DumB1gje
uNm9oUl61wMHwsq10pE/Ey0/DlKqTuBJsc3WvU44kFkxQOnHP3CBS/DRqQQbwJJxMFXcoNmojdKY
SihrAIXCnsP+OuG6hM4qfI5Q73TVgBblU59BNb+/8dXCDaq/wH1dRtGzkJ0FTjPkkx7WzfI/enda
PxD4b6a6KZGrczkBt40u2rXZE1PyhxAZpZPIBhz4sYydwGvpUFm7UoeOtXPKOd4qLA8ynrU/9nD5
/O1YtsQEVx5wAbmbYWR9iYQi+wzsNCe2q2t9Df8HbiRqKLI12Hr4SN0H8cKaQ6EmGzhnRLE9sW/x
twLmtl7eDZC1wsVYdMS+LA0jNqWIkf1m9IEszThRmlGhXZrOoCK+aKXk/1LDdSbS6h5BbFaT+xni
uJZ4A90regFMFGvxpcbcDecaohKrwqX1f6NTb3V9yZ7EcS04kBbEdBOdtvDJRJMJajjbigmyryGn
DIjxEJ7C7fB+k/BxyMHq31FryqZMM8j/Z7N9dQwHdCGk0dU9X6/M71Qwcf8Gc3eLBcZu5Fci4gLU
VvvUQr5bdn9lmMewZPaY9BlI9Upzsa8jz0SGy/qkcooJFgp/SNiestdqqoeZf3HpAyo+VnhLPbH3
Zv5CDacW9Ko3HFJwQ5VEbEazykDb3mRCX/0onSWezH1myelgZfuW35cWjTVcNuocUOJChnOCD1gz
MwUMTnABLxwV4WYIpc1UUCvn9SNd3GxrLrwiQyf5G2nKD10afrSyVtpoEiCE+l1FEvG5P3JUUqyc
2VK8b7WxnCxPSehxTV4ojIC1J7AQpffDqvGJ6s6o1vQPddSADJv01gd2+D5ouBIz1b/GbPb5yafJ
rvEoDl/7kC/USzxxnyoNJNRsD7PxnBMgdq5DCRn0LU/UcXPkHM+Kfalzdk5EoDqTmUyDCTqDAuDz
f4fwi85iuT4IbsFD4avYxQS4aRR6cezkw9cp6u6tQQlO2pMU5QCzcZ1Lc7Z6sF2ooeWg4pSPC3DU
WSzEgidjKCciDr8vWZq92wi7AJGaQfJG9KOWeKmGrSqHZEywoWjyPjdtyJWB4ddNzayQqAucXswB
xqlJCWPq6hk0wBGjZ2iOVGTTd+UwURDgAyi+8QH4F4izzvBiiWZEusYu2XPTJ6SX+hzY7k74mjqe
0FZ8p4+q0HnRQCEpCg73QZ9nNeW0ehi+54gYZsT1Jgf0LOV8hZq32MsQUGRAysApC3lulvShUAFr
Yu0aZdMKh9V9iWz94MGOU/TkexOdrAon6ZVmfRn2OkIRXbmt7op0vEPqvBEZOPp+lk679YgJoqY2
7H7c9EsmjJKdJHPbRVm6diZyw13GwfCqsf34cN7uDj/4TTU0SFKxS9CIlMxCK3LTaFiepF2SlTgY
dD/ghRS7erc9dDuoeUv8tTEIxTSz8oJFFBFdbeuDIkByIg/gWWqqwMP83qhiCUvoduVy1J8FrGNr
kSMe9sMwVsBsp/rrPur05VnAMCSAqXke8bDXJmSwFy2DO6rl27zjrfqJLOl022oTyKHGz9zx9iz4
ramHYZu90bf+tPQLH0B6pWfsCAo4U6/bVoA4B6OcDEQV11evn/SvzRenDxLYwwSUrqyASWYapM+E
UCGGzjalOqQKroNKZRHMl9Ob0vLiHrR0XLz+dLvRodXPTM/r3OO4mJh9H2JGBZnm9/uBbwI9bY8f
g+jbTyf7EdVvdPEnCQoCjj6NIj3X6m5ZlZ4rdjkRNXJj3d4jXFR2lcarUJ8B+UtVhijriP3/l+T1
57oIQP3BLjKZt5aL4AMR0J1LneLXOlSrFlzsX4V9uASy1FjrV55JIIyfxjxvHX5LA+jo3NktT4np
mjr7N2XeJRJEawxJakFfq/1gMG3h6V6lb4a1PrvEK2QyLEP9ta8ADvLZdH26QAl6BxVwqTqSLyue
vAgCyiUGu+aBawhh7wsilwOJybcW9zN/20wVUrGfnnnnutVoMw1fIF91FFxgkrk6TkxvSY1XlLJm
U7uOqjDX/H8ZRLvg0ggPcKZOQl04bMO1rkvEuCKUNOLBKsLNSAbda4OPctvpJeysNa9V61LbJ5Is
c/+G4JufGiNLNQ9M2yQz6hRq20VTQiOwz3sI9tdjOyV/yTQl0JOXfRkFhBgVzITkgTEVHsffKPCI
8gvsOf0Jx9W51PVi5QnkYg6JcIZId3JKdMiPVSCHqRBJMQWa2HrVx77WbUKCO1AJjxXCyKlwlC2h
00U5DvAfspiHbkhJpfNiM4fZnPe08i0tGRKLgEOgop/1n0NcbPdpl/fN3rlIWru4Huiz5MtImC5/
4waGdnBoJgWhc2lcmS7U1ASo3/qGeK3vUraJDG//xR0rCSkmIEtiwxWVwhCI7g0akhqTM/LCTdh0
T40d3e09+vHYbojUVg6ang9cMy1ptzgXilrbqoYYiarzjib+aFtIbtPRgPjGSNqgkU27geIba3LB
jxqV2sfOp9LLkfZv7iTfeQTE1OOgKUpPGPcFwoKZRkARVmI8oFVf52kxu/UeaiaSch6u6XZ3RGQX
u6kamDAk+cbwOEt0po1MX4P5rgmVfbF1SUdQNZ6GWA8oZa/+vfYr0R0rixv+AC+6pd7Ptr2nYdMM
vR4bkL476I4bbslf0k01sdNH9p8UUohabEl8o9B+S0VVzy4DBzdYpNExx29E1eEHU366AXjOKxEm
vHBMkRPLP9VppOCr0Bb40WNRMpND36Pfg1F5UiF1QC+TnLSM5BXYCnzfBQI5RtQ9S4vLpnqGI9Sf
eOXkG6ooNgP/gpda/ATJmYFCMZh+AMW8SUzv2XGfEcJCT7MEidwmLOPMtdZzG03LJds+ZxMV5nZn
h86rZWWDnOhRttTLpI/+acFUY/IPlGU5LURJeAq0MwIoZ4Q5dVe4UWi0ViQrgSEdA3AnJkM9Hw4B
o+TVi3CC01I2LqxPWCcYVvjwRr2edPSoVt1LXU8JC4EpNKpxDvOVFJcCq3KZdKP16jWO4nb/42gQ
foiB4nqOkshu65zqat3QluEXDG9hrFXe8glCtZkEw2D8s6d/vNraYJiNsCKnA2jqLV7JvG7sLo4z
Gtlc8MdY+a4m2xYAJygxlQ+LLl7DNL1T5XsOSZi2cnpAALLEvpXinyzlZDyoqZ988t0zeJ7IIvNY
2CEhQNmcAOLitPUxBLBF0krRJvfU7B/O5E3WNzTX5t/NMNe7fXJY5nqFGuW4ff4+2fxTs9bJrSUv
wDaMouSeTwGRtJI2BRUskYHNpdv65i0idqxgqHKb1YeKWc2dzLtOWcYtmZEJ+g9pzC3xhmITaFPu
GxWYDV8UvORyJhQkX5ybh8qSgUbAqouuEy3jMSmeD9YAE/vTGfCSzC7Pvd8b+LY4NINNe8jrxUCu
xwgctgdzORR4vLGKxr4HYSxOJhMF2Iqmk7Kbv8x6mGP4WquPm94FqEtT2nIpnJ1Qw9+2dsMki2v9
1hHrvY+s5/jXiQOnJjhfiv3v4Z1zaaVTo/A4OmQNcIp3+1o0cxURqjaCwegieLzvf6bdAAXoryt6
mqpRjbiRVNafEUMtjc+fOL4Mzn5aUtDsonYBrTRkBgRSluXgyozYUUoJNI4iA5eRE8/A6ZY/7D+U
u7qfWgOpnB8DGPIhmieyMI4vj1ECcSfxf90l6/0oEDVF/FSYI8SVPnednD97AvgcnLow9PrsCYVc
PCdaWqgFxFeaNlXrumM9iVJsmwfvcw3Gy37nSkuXXYYzZEDd7tnUlvm60AucGFBqbOpwXLxwpoF7
6z7LfaZ2hY9Cxq4y7a5PUgNt49mO9Mduwz4ziRMnQk2rKyHYaWYUIJ8Ay7awxfktTNtE0W8/L6Cp
tuGFB+eG3OxZBCMpZ50j097ezKqqspm48zG/HBqt/6pnjpwrW5tcU1cLCio8JgsAHAWMK7O4oeVQ
ibQkuEg/z1UEod4+9Pmuq312qictz+Av8aUeJJGHHkU66eK3+E0Dwk3ELStBubZyRuprMmAV6PrF
76McWHc6vJZvqCCEikigZpHVbVzKSLjhWowXCKQpef3lWxwSqztPJz/xJkSiIsGx38ERrR5I/URy
8pB7n5SZXfBzz+k/a5xV8Mq5RLk6OsMvLYBtNSUXfyf6+J6deEYFBh7uAt9flppxccOkJo+OA3OP
rpACPVCdCkYKHwL6l5R3RmmJNaz5RlX+G/0J2CHqaVrVNbapQ9wplJa000moj+8zAL7AwYLuZUDe
xHlr4lxcnkdcd21MYu5u8g8qvpnuTaMmjwA8X92BcixiLMni20MazB9a1IqVGfWFlyAjG7ZX4rkR
9EZy6+cVp6NMn3MrMJ8TWCMQl4jFTSSKuoboGYi6VB1aF7m5Pl7/K+Ho4Rknv/AXeSmxSItJtWVq
hyiRjFGte/0r9pXFz0FzdHQ4Acj2gzrTmn9NgqJI7v4jzzud3JvTUu/TuvpcswsrrygA+hzm8hn3
v8AhIhs37ZU4dY5DBoN11n8okFo+YEwcXlXN+RpKaIVjfMuCljgyWRNtqW01bllGJjbWeIITJ5Lr
gn1kC5+dm5PSo+Lh+QMoO4a2zxrArD3/UCl/7+EiSRLtCX23Mh+U5b/Zzc/1xdhdyBNskhc6wtXW
mAUSNXQtDbQL9gVnPVM69V3OmRzVrwOF+fow+H7EDvD3Leh9UtW5L+cMe/yxwEF65Riof1Dy0MX0
9GVYX6ZcMOxnEyeNCTjalUzIo5gwUZbLkhDIjWP/jS4Kl9qLB24VLivOlwrk9WzRJirTTXw0mCEv
bZ9VNnXP1H5ZyHzvPNBebZCbBNYDzbZF3YBHMLedAoKJsj0ssIa3/06jLe/8ekSxjXNzPGV08Nrl
JfLOJMKV2yHCmSmuAlnBIUKfg7L1qnPa6dnqSJmjNTRglcMWknNakkiRn+24gr7OQ9+uPd/z5ESx
9kICDT/x1POLePLlKOXC87ue0BIEPAwJDJFa9wal+4jcXonFbwKW0InJ+ZsSxuwu6wzp4ezfa7bM
2XuOhvH6ByLpNNq5DoZLw4P3Ab2oX5vAP++3AzryD57qJ5lKqZBQfGE+89F3MG9fib35i56kCbgE
9NrX6paa5IeiLO8AAajzeFg/Ifc5Ce+tvLwCYMYKHPyybdT8CHkaPo55E9F66wursiYXcXJIb00r
tSF3XqUzE0c1YjcTOpdMiDuqLJKBsEanHqL0uRk0mDe+er5Kd3XND6+JxwVvW6kLr6Xmdrh1tUNJ
9hWw4wZGmvgWLuOk9CK9NadMWKsFjhm+LPXlP/dtVev9EcOKgLePu4dEYyTt5FBEAZrZT1+IeACO
MkdzF+2/YNPcHQU/Q39NCww59+D+RwKGvf6RcYJRED02Ahmm8W1BdyUb33tkHG6ClvMDpYzw0vq7
IefUXoxzuwisL2AXWns06QwAsAOjQ5uOIwSs9gibhdjY4OmUexz46LUku+7nsDAH6178RPgmn4Ql
Mr+HrXukHJUjO07CYt6/5chcp5b8Fw6GvJ3Pyq4NjfABcTWMosyZUIiHVxJ4SN/7WvUHSdyDZAN3
Vy49UqaBu+JbnD8rPRu1bZLvqWgnP1fa9F1z4jC+rRUUnvmL+hr0ghxnVyQ90Gb1fbCixaUoWrkJ
brj4gySpBH0/Fnk7gjLGJZUfUwJvnON3BjqQfPCjdrgaNim8XVye9ZeEJRVgRINceAY/orQATolg
1Fv871jc/3X2lsFinjjgiBc1oLY+PyAdFS0bFNx4sMiWhjV/KVcXCAlXQXgh9WYwI32buLaFyQdL
D7kqzxEL85QiTxmnZI39b37hi6JDZ3hUJuTVg0PDZHXdYvvHzkuTzQMLwAMX7x3jn623PqKNBifL
RCFbYusw8Efo6AVqyXBNt0Rp6y/sDCTgB9ZopV8BnMLfYJ7RxoRqamV986RN8WwEql3+9jyc0V5D
bPTrRMImsAnNs6qct4vT7ZbBYI9fYwiTMu9jmgviDUZ6M7s1XysrYTKl66FC81GuZXGcQP3Tdjgj
XWiZQ5LGV6MDjwLgUwlqSks3ETTUScJHZ0AR/lKjVCxtBvLLF/6+leTRrnx3Hs73+yEQO2puDRnh
3oc60UJkfrjX7Lp0PwECePvElOylD2m/Gssp89lb2gqCnvY+05KTwVyx7PKcDEtgG7GRPFugXhuj
4F1LXIv8qSact9svcRuSqYWGeablb8xg4I7ZxnjUzVu9bvRD5fWdmC3xdSdKC55B2U9eaz5f2qSn
Jy/e6N9oAUEADL9f14ydQTeXXF10M01Gv6EyGvT60lPzNt2kmSI9LN4tybUfBRKyjtiQEvoJ92ca
9ZRd3LwqI+HOiIZsHn0sWrEMHD9w6qEGESYCUBXYjDkuat5mzuSg18q4k59heGhMu5QW+NYbpsUa
LGNcf7cnif5Jsgh8hhra1ZaLfjyn1ezxTV2ji7STMhhdKu1hkfiN9UFw/BPCVyp1m5GocanOEqpV
2C+3GxyN4ZmcvzWn7vC8LiTIKa5I8nHeA1bAsaTj/7SpJ8uqZ1fikHGrs99/WtHnI0BnXoko8YQC
iSB6l0M85eNDgLDzjnIgggIiHiyTh/8mPRhiD3ar+BnWLk8hVKRyXg3Jiym9noea5T7nnaLTFWSr
OTNRehrLPs4wsDfy5aGl1R9VN/FDiYRcj0sDOAUNdB0RKKyskBh0Hd9ekw42Vvo861jG2HAn2Tbn
jzUwiBCethfHNg988sw7GO4XcjP0M097HwrzYPK4wrC10UroDWIl7c57umuMxryZ80i2ME742H89
qGEylzPQjMvnovMBUqUfF/cOcCYOhDpETKS9n8wL00jxkwEyS9kOALHEVhD7+4RBVgh6UfUarMiF
h92vqcBLrY8g7LUkhzqzYQ3AHJuJCkgoviE58pZ4LSoCZrC9Tl03Fr9wHBbU3wWvwAKKWSEwHTJ4
xCP8TNRP+iBpd1piNAP6hz1lKE1Cl46tFh9FLFQHxNgk86ssifLeav9JAddmrpWh636s/aB0fjmZ
rWY9fRCIFjlGlYEalSdRPYEbHvhBrscuBhhSMC1dqZ9lpi6ULAeACQoZHyC8beLk0PCCYCh77VJU
ETzApFAWEWkVfSVc/j6717pctjHE7RAdNrona+WaVG8D9WQA1EMYtBh6dsFAPzb1ggMTiK14q6h8
vsqFd9ggI5C2UGCYUo8zx/t9a28SnNzZVCpSJB3MIckJ/f5coUGJxxz3qtVfJekwfXiZ+G+ki6hb
ln3TfjnmdbZPba5PcyFdsvSwBmH22nk4IKb3edVcwnj1hchR1Cm0yKPhegp1nyxFbSxJCmHc+8i8
b9AZdYK+OJn2TvvWzm5OkBek8DdWVaGPfqLqIk+H5dRTGQ4dXjlID2hbkzqi7KGBfpqqcoxSp2i/
U6Y70saSLWzB398Jq5Ldv+iZ4mNe8goOlNbKQnMZ0S3/m+bCsxxN1WjKXTZnq4NSetEQqRMLjd2H
xlu8qBipv/qW64DRiVytFQtQOXvbU+p9jZBUOkeOelfgauS+52BpeK4XKf9neLa62asfPB9J/krN
fv78Jh/yb7B+rjAbprL3nWj3+kuhl4DZ/2tV6Y8pS0zuoJVW8NUrPlP5KyrXngel9IiwANHjCBcX
j8xeFbpkJgC3Fij3wihJIJIfZKHGS98QYFVE5XHdFDMst/1/KEqmWepVWeKmJ4UG7v7vCWJ276zu
WLpTRlAwuJJk/oLUPuaA0zVA5Z6WX4iNC3XWfYnJzu8eEsqkGCEfwqy3A6CuZGR2mF+t9oORPiel
pzyd9xbWkqHKMlTuJhLgAh1ecCFiDtrCqrq93xn6vTa5FglZTr6ka++R/3fnlE8LOCKOEojGDBwN
XxJFDdWnWAQpq1HPUNQAL6UpL7RW6XQOjbCYg0fv9YMbghBrZaLJBZHxnC76EbpxyfItfnTy6u+2
f/kWhlafnB5i4c07KLSEq/jajmrMzLinXJ9dzH2ZRgp8iaMHs9/XUWd8+0OaiYrM50hz3bCtxXvV
VIlr5FpnPuws52x0rw6e+NahHYzojAk5x6+vs9dCXmTbWWUzqcPCOgGxgXBcDkHAFsepadfNrjiu
xLs9Wij7V+FnXkHrTzaMwpIvWyUbp/E4yD20NaXu+5n8LGhWSwoSoi077bvK/NtfCJhW4u+4KLU/
PgXNTKccwEY9yji9UMc4F8l0y7/eWX5DHScO+K8zn4VBRjCluJ0Ul50B1sZBox7eLUdF7EmF6JDY
K++MUM6XydChCHZDnbDVRXU3LEUQTNnMXvVqk7PB+Rn7ZPXFIQKiP7Aj4PGCY5rvy9lQkmGRVYG7
MG4TqlmzrELVMkOGqezSnbek2WuqicAwqM7dZL01wDDxtW5HgwfKLHI93gRPA3GrGyDHoFKOTzQs
/NgVhcpv5qwHzWXqnyfnTrM8V99zjSDSftRNUdGvwkSYiN2Wn2gnhs73VHVztDcMBagtDD6cuQUh
wLQvCMRiZHR1r/zQH+uH7x27pdxbhrDNbH6/lL/blx488A/pU1MskpCffJGO2Vo+NHHXo2byGO5w
KDZbck4d5cZ9GsblasGre3W++CwRTT0l4NvJNdruC7bYAvigdGvfn8k+KLcPvTgVtLEfFh175vbr
xvvN9iK4TqJ5PaEDKS2KUmEtifKKrSkzpAPt4B2IPZMdDA1kr5YXmHse6lsXfD6B/KJqWrXDFTSk
qb0qlpzSE+aD/MysMFrrrAzlet+u/zNHePTY0EDTQ4FjBjqSQvrqM4AIqbqv8pcSlMtzO6CfwBLq
Ql1nKShnVBmtE+aDRR9msDA7bX5Hx6K7t7qpRHR2aDjo9vMrqy3fpYGVFb2Qh14APLmqoDqdAFo+
scNPJvRIfP2cK5NiDZ+7wk1asEuP1bNzxwEG581Xsk89GIU51V9fXTVLLF+EJtyXmbXDxvkYZjlZ
w++uKG08lLCRz+SXQjIu2N7amF8DYNz9ZAHE2FSsbYjt0mnbs19G4XVUlz8TlWZvrerGz43uJeSj
Sowxqb6/y88c2iW4sugvx1MpWlbb21KlZKex3P+wWgmBQ0HYFJbIuubG1ho+/M4C3beVPQhoD4Ac
2/mewGGAASGjhuUlKR/SMJy5dV80Iq0tV8X8ehPl8UG5ZplzmSJoNMb7hS5JAk3xAFAtQqSCztEw
0nTYn8RiMbEfMvH9dSt/6nS/MYwXkKrO6u/fbpGB4B0simr17EhpQbjhbhj5nvD7YkPDKIrgA298
ZLwXL2+ScQUkShs9yEt+Esp08CvH1XRuoXUcNAHTBS0aMIAfxnw/V7etZj1CHbw8VsGKm4vOnqwe
RP3gamZIQsp2zlkA7komJXFgSUrZoNFUhFrpCCnM+u41N1Ii4lx1AQHfRcsuDHV94x+zhnBY+Ws2
DNL4fm3D8JHvR3PetLpbaxG4nM0EleZZumgx1I8jv37BuOUy90KP4Cd/hzUM3I8Vihf5ESKugCQP
MY3PAnj5tbtjz1kz4wXCH6PjcsNyWZjlYqLhlXTYNo59k9eAHpG/Fmt6UGp7FQqknVW9n5UEEiDi
B0mcUXykhTdLMUMw6RP98nYKVzqwbpTcZsc+yxRly9ocspw/hGvIc5r3hlcyibMJEM1qQbMfLLJy
htUj0GBbRPahqfTBLvjMxPwAcEJzydJDFEqfMDfKVyrtq/98hnGtVvWMqReik3FlfVX9lMXNKEx+
DysXeULZOGAZsZup6ltMhuL0LcmlqunvxkJzflXxfZtmpzdWYrUppMK8RRYd59PY6StJEkzhZMfw
Ck+UQERL710zQu6eRJaftdBYSf6wlyIWiNp0/yyXIpTPs1vh/K2DToLQxJiE2TG5OH18IhrhJhtg
YGd6cVkeqaYjqpDd4ykbv4BskC0PKSPT9YKAviMiAFl8VR4OAGmLY7hglYIvI6Ktv/5Ji7N2Mc+W
u03096Tjy6cIBtR7RGsutT+70r4KLnHGQQvaiX4Z3E0UU4tAx55avDl4UFBcb7m0OZGzdGf7CZRD
8gWTJCyXA9ZvzxBXZ52AegutUlDdxhUdfVNZClLyx1hOnzdHMDy7okzOh6nuabooLDrksBFGinwN
H96/GfT+/IwlnUjm54FW3CmOIOXwaTf65cYjWLV08TSJHlxcWkGjH7USm5r7Nw0eGihtYHJpsg2N
J31+QvVHmLDU4lTL6a0/ItjmQgrxZymDA5oaJSBOzSauT/GTMNvcJrcMRYc22fABj1cavpEpCedV
KRqVkGV6cn4mMeZCxxk2l2MBknK3LRA4kGU0Itp3R9Sj38OocF2j/prf1ettR/VfeDn/PiHCNKTX
j6lZAcjRMm7MdyI/Pi4wNBl+h7TrTxleS5Fu0ginpRWh5wz3oDq/KHJps/VqpTig0YRxbYUE/r9n
RCUxNlfR55VzVr4ZrkIYChwDDgjwNIuObRbyYHbMwt9XPQY4Qb5LAOIw4vbWteTU8I5TXO1hjsaV
acjG6va2192dVoNBckzTkpYiUvM+Rzuf6YzPhehMypSMcMno5wLFuJrDuZeyg7XBECl2jWL91wEj
+vfFvlgHgdJZZxvHu0ENbXIePtOmX9ZZR8VIyM8EuaZmGCKCjb51hv0QKkG1jACm+aKCOH8/RTch
3ZMU1YPZTl6nhFgvg6e5gY8KMv/ZXafVGIuaC02l24/hzMDi6HzUCJSErJ9LpNTOfbX9CsblDNxG
23/2U8wtlccZUl+SBnY+9Vzyj5pAroU1oxEyOfkYW13wcHf4fs14ElA28twx9wG/HB8+CeXnCME8
w4JHVEKofCOxYC7uD5eY+bEnIJRVK1bwkT89mAcKdMx1x+8wmWkz+R2Ok98e7jAU6DlNfjQ4qxLt
0z2oWdsdkTdxg/5o1JHGCTIEjK9tunQ/T9C1AsTTO5/3dlxfGWKZqSt56Hvngggi7E7LlEasPiES
0ksR2TYYeb0jxZA3ZVgJQPd/vB3CkzEcWuxd9Dxpgl4dPCOHjbqV1rZfUb8Xqof/XybF3cnWLUwd
d64dH8ZuXO0FBPZXlAhX/YPPmgbBWDtNBSA66xZZJvgQDRBlpK2DmaEABbTefUzl7ybSrSr+RqO3
qb1hSAaQhQm+yhZrCa5koihodNRim4jgi1hOJOdPpKFhyOM/yPY8pgYcXTSykjGrGkTcnlt22xgJ
E4RItGZnC6ekGWJ463aDpY/9mB+JqFpxLQp+dq5Bgw1+XsgJUS2ienW8zFR55fia/a8bCRpIhEdC
fkizyCW/Rmez7R0TiPxm1F1YlE6K9ytIJV+hd+ONmN7nmmjDuruC8e6/3bl2X2FP4K2fn6GtWp6r
rBsDKRLYXjgB1z9pfdsYCbJpNEQQN7H9XnTtEMJ6KaJLvWZf5htKfRx/UggijuyvrF9iaYpeTvcZ
CApLQ3QMQ+xiZybA/NWhpZRh9HbxpfeCKNuv1poJfVU41fMF74qWIMXr2iQ2pTKFRoHVY5kyHw7m
DBGGYtdXhB2LWWPFsvhIuiT7p1QIKkw7cHKeTC+fYuhU5k0LGlSk7XTmmka302CtpdZqdKz9ibP3
LXc8D/RdyVnJo78sIWdqTgLbG9RFDQhJkzLIW0elib29pQhjjMPnxUsUsatYz5+EjDT9xCVIAaaq
cgXPLVl8VVlaJFC4tjr/lVrn6fqOKGzHDjsiDKjVADkfvYD8PGMYAlaZhxId4K6+INS/iN1b8LVH
M9NSgYBG0UZEs4xKXRIoXH1RL2J22JPZOHolJpHXfoJVIKhnJykaA0T6zlGk9mUGLBXN3Fcx6RWk
hb+zbI320TLeKfiImRqXeM3MKZOdDeLNoA3W4kOfDPKDSRpgECcUCOVmdq1RDwy8EZcA9KgETbNh
HMNfEDsaXylFuUa7/KHLqxTF25/ZcqG1g/6ZVtA+bELmHCgmcAvCpXg7lebtOSJ8ZKW4E4JyqGls
yTjjCf8D90iRSfv9licKEt9H/8YUky5b6fcC93P5k5Hso/HHH77Zuel9fYekhQu6HaF01eqDp2vg
Zqvg9eSh5W2eZiVatgizvHqkJQs55VkuAJ9LgMESdPVCHPjidCuGnbmdI6d320S0IvVlkVtNkJ36
VLerWzZQxzvKovLgZEKss89UhCcWvVogF9ZbmdsOe8tI/r7KOlEFj56sqXKlrkIcOut2hgfOgcLi
lvbXZYXzSwMJj8tckQYfwLuRxWlvECZhhrXeJQwh01o9nF48J94rDeMYk1rhHdgVTAYNjybp1AuD
CQBdRwEkEaJ0ykxYDlGW0k71NZMuyaAvlC0VtI8OT09Vr2WhgJxJ142B6t/BGQ86p2zysIbNHgfA
avDVAr2ziAF+f+87M8lcWWpSScxDqN/KOTSEMn/mi+/hqgZTketNkfAzMyoiO0SzpIlB/FzY4P8l
OHYPomYszp2z9HWOlBVRAVaAx9VMvla3ixZyjFvN80OZ6zIADF4fpiLCrl4i70kQ6e3JZ0u/y+e3
skQ1LXGoAbf0nvKoTWhvYLhaeZ0EizDvdf6oVL5ZSngc5LPE3wxywNAVWiL4N6XnhFjM/aZ1PYEb
UsowgAhjw0sldXvALG0qFgwryo5+/0YsBzN0TDgOQ5SdAsc0sdpvMMCCMxF40eWhU4+DFRynzinI
+bApszb8kcLb6fLrVKPj4LlrEg94Q+jxpd/I/p9fQbHnoRh0VcbjPosou862ztTuvnb/L+CaJNUg
OWcerbxA1Xp+PmDeA1qVm9aKqziaRYZyYA2r1ToJ4qVlFx1TwOLcXYZ2/rArFoQtpqNmMvb5canh
g/EhWmqJ7G8JC8nzTC/CMxDngV51sQKz1ajQT0MtsgSF2EYm9ZwOv4yRpohfDO6MounSqA97hDpu
992sq5GhTDQ/x3gKxxbtRqUvarRRBoO59/iD9g4L8zzM1zsQkR/wpuKloMRJ1wyup2S9W9vi+skr
NzMz3ToVPIfnd/O5+weUcOPkVAd9sBiN0hjYY5mELVsQIY7BGe6p3be9Sf1BUmeC64g8IQ4U3wzM
icuG8lmF+5DH/5cyUhioqHve3hYp+wE6gu8NYbhbZVVCHzP7NICEUpVsjeFBpaPzUgx4CAYuO624
ZxIVtUUje7ObsFv2hmSDrc1q3ZjcVrukY2qAoRwrTbPBXMZyeT6hhjCGvKNV3jjx7qoZMkzUMt5A
VXrcx3GE7lQKKLeZu9i6I8Mfi/QpFH3i1Al5a8QovOwx+TzXnjwHd6Mk4nmh41MTWL5aT7/r2FKO
m9N3V3+G3qNZLfGnOwV1OG2/TyXnELBg8fluoGPcrF9zAhUfNzWm72Cnbw8Kow8qEkd5tpnjNxH7
PWRivIVdt++Zj36MMMuhhFEeneysqHAz9OaDeraWDHxCQ4iRM4iMXu+RhTbGU0y6w9mD6DZFF2kv
4LvC8EYltgINfAWjXrJD+H7GwBp6PAqRYVmRlcSRupdaLNZAOuAX9Sbo7WGOLXDcWnInw4irHCRU
US0cREdwd/ywA2obXD3X8fgf0WwPLZ1NxJ6d1V4BMNe9Ex3/SPY+tLjS6lgyiE3NhS1l/V8Rt6IE
sdD9tyugaayVchsbt5k87xS8Wq81O9eE1uP1vSlswhPdia3/1VQogSftFX3aOitrPLKTe67jjaJt
j4uDrSV1s6dKn3ZyMbPb31kckzJaNEVAQxgWUbeL7ZcLZ4JWUU7MUsDtb1wO1HJE1n17YbsKu/Nw
OT4vIpm7cj3WEseW7XacLopa7rgtNgzPF8oEleMBGkT0V4OxpopEPlhleSp2dcUaY3HjC8TyoaaC
/zZPPNCuc5qUMrQGBU4nw0kzQ/I9z+pt9qZ5dGFXnhJ/SVTt8cIUE9DeBQB7g4xoK5w9VWs1TqRW
Ft91gfktEi5ssH4yxpkWC31FsyIyRxmZYD/Me2vS0PYy4nEz8SIXwuLkMIhJKF7AHqk9U60aPQy9
Qg5kuJQAzxP3X6qXbIkKXEm89eXBbtH3ovKjs17H6IEqPghUc7R4mW9l7xC5T1pAhBwyGR+TsVCY
QN9fWaMIvvTLzp/EVpTJw4q1JRa+P+IqEAqBr+V8MFKIUGVFWofbdOkMPCV2Jzzpqiqymo30Ute0
jtnlxyllVa4Z5jXgABWfdw8aCWxsNj+vZVJbfv6JndGo2wAcbr17uMMbnI4WVDP4+MdOd+4NCE8o
iuL3EztVj69lCMbHin4hEXISm2h/20jKTrCH8duQzE7YcO4NYEiiTWDeWpU0LZHcQRT+DaOzMzTA
CSeXX3A80/q9gpXD4YK0UMsxxkBPQfBMdFzffn7VV4RESbGDVUkfk6bgG6c5SG7iPE4tSQtT0O3K
ph630obS0YJ/4GsCtONaO+HIhIsiWFS4cHz95c1tmGrpTTw6dOCxV4ohsx90ozGlfM4ZDjsupYBg
XdAdQ5KDRNp//bdHgZYwEhTkYWnhogDpWwfrQnP9HpmvLAC/+QItglkqAyZVuDwU2n3zwclK4my+
+KAhIvaEOac7PM44pUX2vmQ/K7kP1PIhgO1+yjEajXSimcqJqp2+JS4z0nJvpEtMbm05JWllYosp
ZSe0hop6sOX1u6e6XvQgKMw+9Toz7hCrP5BXl50ESxuJuLJxrZiKJrvIL8uR9iW1NJKWiwoTFuWS
4tXZuAn61IgtNoqi+BvJksfy/soVLG8aGPXbrd23ZptrEa5CCtflM3QeYEWXRGvsqEWb3pZYTkVE
DcXzCNxDHF4HGqbFu9UDQD/QzmKmW/GXwmTY5THz6jVIqNJK41V3fLXAJIh2CYDfzaWTBAdExYFf
PjHXs2GfH82MVBQmHx7MvWAMP9PLINXBSJyaSesN/ihulpWqjonqN03s+25ut/r2eT9t7FkXqBg6
L1qYP7tsEuUbNc6XcJ5udg+XlLmNCyZTZjfRu9TiStjxuenz5aJWHuYliMXfTSHhyjntaOwmD+JA
3Kb3OgqheBjL8DEbX1JPtM1U9n/hJSNUDO2h0FKAICE6Wrezbq6CzkGiyOyDXVCR9yTjIOFAlLbu
aHz9G911wihQyduIUZ5caOoKokOMvgqSkAAUFaOOGD65XZGNjHG8VlfE98I3ILZs/XT+pZRGyosx
mxANChGzpGmtBItCBbfXSt3mYMn8T++3NUx16BkHBBitzZoGHMhpUZHOtFmiud2nNQsO7O3yuNLX
h+ZdRWEZgNzvyhbxyyXHPnaCybzCiqFIlEPC33Bj6+HOuonMDHP1Dtx+N0hGCqIK7QfFNrA1qXan
HOuMAzHxbYvlVqPwr9V/IKuEpUUpw3jkSzxYg2WqhCIKMF9MAhcJDnFre6RS3K7u9W3KFm3eno7u
DFGmcIMAwS94siFwew+4HpsayGFlTJPJmwhFTHhFeBaZEEQ2ulKB+UO6mIXz1mHwXIFoV4qWb1M/
EIkwwwDpIFuQIAJjzLvYikZhRqPuAj1SEErVwpsz8USyJoQFiYX54QuxC4a6zhxH/LqWmcaWXJC6
n2hlNCQ+QdzfV7QgVZ4kh2qdnDpNHHIDPkFcA1nPvwIH3k+T9a1mgCIejtsqjEUEuhnPApih7HFe
qU6EZucGi3wjLH+CvxgsBeBKSM8NZbri07HDysYBpljjnGN5Klm6X/wWa+UPOuV3vmwj+ExWnEa6
THlWutU2qUEB+9vSd/Danf/Ibm6AKtidSJKNV/B19IcbohnZXEwmMf70470Ar/Ma3ZHOyrPdLdZO
26A5OSo1Is5ndRsB56EDSbJnP4biJrq5ziosFvhsb8Ut9EdlBoeLmsFHcVWq+7Th6F4ZoQwS/iNh
ECe0K4j+lSwzWmrFZYI5aeyO/svMXp6DJdSWUmdlNEAXaHhkGUgY7DkceiDmt7X02Wb8aRqStLda
hmv7gSZws5PCa10FDeP/aiY5Jic6apspzQhiHeH9hMVFCXJJh541Xj4Zkf0QW2jEJSqzi/pGRkqC
VbNwMRuEZtEczq+d8vQTkvtYhJfjNJAaeYc29n8sYX2QCLzHxHmzaV9DElQ1bUJa9gAoh/Fe5Szy
yyBDyw3Foa+wNPqvr5Hpuz3+0egA0e6t630/8oCPVJql0tiDlvDAqPb5b7mbhyzo3l5w67fb75Hw
PpquQFjKdq23tHrGiC0an35JIAHJZNxy/CfF2/lLXz73YpzBXqxPuD6oQMdnq3TrH+07gW0tKovJ
fWEeVcqn/v9+Y8b6HQ9aGRgBm+cMfAp6Kfl28eMzRhb8iaUkRm7uITyBs2Oe7J4sW7f4A1FETifq
JnLhOn+CUVzY0skQ1F2oEARbBfQbCl3NxxNlWKNeeWHaOxUlq2sV5xWmxFTYbjjRbQa0H8dplwbt
1RXsgCDW0Z3YMpj73rEv/pYMpRMwuYD/434mi4y08ZqQmk2jx/i1rUcbvMccsyBKMQo302VQ8470
VaoES4cdRUVyk5Y5dufYVwRfuhKljMpFuvOnr8yFAm5GGaycIvvB61TDbyuT0XLBiVIEA3uXHQ6J
TFb9QdsoTpUF12ecp1N5wXOe86DJ8J8bEU1I/CrEkgMZQNXlMS7jp2NuUTfQv84JslYbcTdbrEj7
Z3SS+RPMhjocVvSVt+Um0CXtNFMwv47BD+vGx2Z2J59lqntmjBw6SNSyWsWSJ4dZ1rHK6YX4VTlU
G0MNfGNzUQmMd9WyunioGVFa8zq8Ob53a87Psdy/2UIxub1VriG8ceu7m2imZPjLWe2fn7mJ476F
CJ5WDvCocTW45Cxo3WInmGnnWmsAQxpuc+FvvSCBjfmNUEFMjTzY6BJI4MIECfrIXNbhH3VTI0dC
KI7fi1D2q7bHdMZBAWdr1gsN51VIs3/LMLZBNw7vDgbsmTQ5nTJYVGjBkXjBeWuaAx8qjqmGaEET
NM3g1k/tnGF4AsKMQYvyYmMyuzVUSD/K3D8BXwYQIwyZNjqpCa89/ZLwmJQp2AWljBKuJBCTcXhW
cJhgroyhk9HXPPi6Xp5M30ocTeyMO6ANqC7qA80Ii+Cj475hrDY2s0beq2BSjmgqSP7XI8q14n9r
HHiLdh0cWM4aydCDptqQPRav+kiv4b9voydQLhCrWWA/OhSn4EgqX1xxhQ9+VfJoYf24ldxu+Qkw
ZAWjwPf7y3s6K46KBOgvKjpeCmLYpxp4JpXfWQo4TDaLEB1koGZlEFd8gt7KgE8L9ZHNgKfI0b/4
y3/cXhkk1STdu1KO2wOHjTilauUVQ/kYh0wtHryvEoHxXaidS9RE3uPv1TY7Ltd5NmDGvv7xvMLu
lGJBC68sIcVE3upQEfXQ0AMWhNLBW1kZXzm4LBMU9lSeB/Uzsy9ojGgjCKc7Lkf3ABdPuB4sO2gq
H63Hg84u3sa7nwXCllXj79mrBtG7y/W7aK4q7fblFDFh0i41SLU4XFMH7N48CxFqnWnjaKPoC8BI
Rx3Teal9Azixu3Xr4BWNVeSOEC3uxxjIfEpG35LP1kmOKUBIjhe46XPSWUR17Qsrd2DlDgNs/pg0
BHDQxqigOHugH9GBwwEhx5a3rSPd8oClCoiqFavec9gXC1GJHgSpbTO5vpLiKhTNkDY+gGxPRzEs
YJcW44aPzNLABGnSBpu3KQADANX81kBvg4WoNYcu0Lio/APmDZ+XWxK7pDVhEdIQZxvn0zS6axat
3A7cPY+UX3GzB1sYlbGsREzzNCGG1AlxaAkH9mTlwzBL7leyDygPCdqBxtlsGOpEkg5wW03QozaM
mL+dZXwVOxtDNhyAf0TcD+/TwN3znGxogfT4jP3S3ki/uKyF0KMpwDOx0MAXdD0XthQ+RMQKgfRt
W7n9IC3Mk1ZvOnX9nzF/dTHs6U73nWm5gaw+Da40ejiMvD3Um0p610OPyN2A3AZsZoSuNcCL4dqj
OXBCo9iHMMUlpMm4T4eaFWK7aFU6CIai5Ds/PFH6FwMq34L+wETsPHzNQ6xhMuDpVv+BGayIV4Ir
RsT0B9wnBz/KKUeVGuxb9N4AEBdySXWhIe0NElRjNXcWDt6zJVaYilf3f7Bk3L4DaTZvBlwkgVAI
UMRf9cA+lQ0LpeHLfPJWjp9iJe+5RYzwuGyKHwdXxPnV8qHWc5xeE2yVwvOtm4NY2JqASzvyg8Iy
UQjxcKkc6JHvHTALJTGjJoSPlXlFtstBHzpq0DXw3FowgamQbCmA0NAwAT4l95WZbg+VBGx6wUPn
u3ekFIhtTXhO+2dJEwmtxz22oKqgm8t/95LvTYMfR+P9am/jMaLLTZAVq858M7KlwOwFaVTfu6e8
X+36ddaNPGCnkIcG4+EBbtmura8S0MFIOnh18UxBZ2upuG2iyZpFfirztRU2J5Iu+rH1HJXoQS20
4xaZ6wIwnLevDNsA7uLMM6xiS3uEyV24rsPvsXcYIl6Bz8z6b11Kif2D1AD9Qqzv5b0iXMGSvRok
KOu9Cm10c466BqYwyLsj7gywZdkyedZAooOpI9FuX98HcDsVjZw8onGP1ns4txuLCfNwtaBaa62K
+0QlOh8VQ3Dyann03YqJwxj+i5yygfNeYbP1eKSoRoHy8OqTTwU3ZuMYDWnLuEsrZ078iuBDBrZC
944YdABbHRJ9uRDdOZLPL2KS0NsIgzprFI9Kzuk7FWWRQ5am7E9LIeIiTj6HsGV1+U2ms/bIEOo2
hQ40d3sZc1UWHF/m6gvSaQ7wULi4d/SXhhdgbT5O2009XVSSdiWSbev61lbOyLfwHo3aTfaYH+UY
3N2Eer/8OoH6KT9CYuQmigedy7BSTujD9pozlzvAPLjuBSnI07bcaMhJfkETfkyG2Erxby/avc5T
ukJQricJwOHDGXydZenjkoh4OY6W+KlhbabAt1J2jmTKtW0rynDZY6s55V0EFVQk94NX/EM0TmDw
vlCf+ZH7Iegt0i/+H4NKbotDi4SfF/RjiXf8W04tesiD2KfY+/x64R+xiD8uT+uB+vAZZAGLsLtm
p+OwcriqC+nHe2Bg3e5DJgAdRGBApLxZk13mbrnfvTprBmGKNKDPppYKMOtv3sqs1akdoehKOJ3p
8It/8wNFB5Y9hzdcYGsoldhgXvZWWqwzDb9rduWP04fZgOKWfW2KhwXXsutOVUk4ailiUSoT5kQM
8b+y0GEDRPG8oEZMwLnwXGyKtCyp90KxrbkTJbtxuyROTDanMzjHxB3DGLToIiIeWQypal4EDTEs
dLRzztp2awica06inHnJlMnSThJnUyBVwPaQHkV9ufpbFXwUqUr3oH/X7vZOeVCCsFXTRA7SM8+4
T9Jet+kvlyM0CUXZMpqGxqXq1b0MvH7LMvwrkgoqNvm4HYJ04i9TiQGG5ZT/ib+DqceLYWLYXL73
JqL9maAiwwyHBrtKG5y5LXHLBqBcclFl/+uhAmXVGpV2tybCOUP7po4IsVIcHJbrri5UMC7BzvCI
bh0Kx7qD/CdaebM7U6xAAfTwh7vvx1XGJc+WVrDlhah2TWvEkdgwbXZUazdLsLB2oIsTp5++aXND
BpE4KBrL1W9HNnesx7UDZ1afpprhnsdmWdxxUVbf7uqYzZVhgSUm1vMWGzVdL6e6ep/Quo3HFwRG
+ovwA7siuCqyoVFPLHKUiKDdy8vMexFzP4uiG3uaK3OMJQw8U0Uv8RqcK3lbR6exitLXtxGbIwjS
RubqgyNDpWXCRG1OxvzaKWEjYLiykuEIJdCtqfRlNK1dXX90dmwr/IV9RzFF+8BhWSWbk3Jj8uHy
BR3bpvy281eM0OgioZpPKLx+CR/Hv2kuaqQRLOw+Cl5ptYc2Ut7Q/Of3kkIlewOQHylHcreq1e3n
4o0L+jeeGTigouILztWxb/8CTPAbpl1ri/TvXylzOTY6zhhXDm6WtkwjF9Oj9hIngJr2qwnn/ZzG
hPkjRDQCVhep1ZdtBg/MCrWrnbTgcIyWZ+/qmaofgNSerZYvvbIF3snQF/Dag2PrBQ0atnl1FZH5
wR/98zP+Z/6Q8LAE31qk9Ei+nb5sifZ5boT7HqCpyi/cWU727CUAH0mol+KTonTsGWfBGhKYRPH6
g8ylrr0gzTCui/mG3xxT6OJDgKpfhPfrv1p9Uj35dbDEt7XitFsx6i6GoJ7lM2z4C9I1mS47cFON
0j9vt0cTKUGozR9coxdq9XyPFGIYbhQIi45tCzoolAl0HwqcmEUa5z7FBtPOW4nTpsONWhgTdvu3
dMZD1WQ87/jjJOeBXZ79835mQ6zQY/UMcpA10PEcdpbdVlh1WehbLHWderpfhC1iU1sQmwX4emeC
F4s2ma4//7me0QGLOOxhUb+/cnhoqXGldGiE0WiGZ96N8X2+AkSVbn0UULrXyyqSMpiJCti7645Q
cB6qV7kNtGrZJa03jmd6ItNjgel6Bv3S+0SOiHczjGIQoEWm5ENiZNRv/zosTdW+t9CBg7cd5jHh
Fw6X6gcviZsEtOlxJNh9CuZlaW+8Apfc9WYqlH+Nf3wcmosR3KYbSr78tNSaH6CQfr1hBXpRystG
TXktsjETJAqbYPlwNHKwAGq+xfum3mxp8WSoN7GSEzR21WzQqpmq9qtxfbSD55AhVkxiNzrfZoIu
5dLD/Xt9N10/sXwEnZk28v1cOGRcTgBG3g4dFeP1YX5SGzI7WPFdgZwznpzAanIMoMlImSkKVU7e
F0UxES2LOzF4Cx4yHcinoF2oLb9SorZupISu0itNt7ZQBb9e/4yFg1ON/eqVB6pLTD6Dqq5FsXFM
Pu7MXZLEMAgp8lfo4oQ2D3Fls5PT0lvgkJJJ1iP4nINFISIxqJtpjQZNoW7rZCRCEGEPscmR7PoT
Q2Isx5pmmKybf/WcTDjQqUEMHiw7IudLv75holAVa4xObeGkXm/0oWZgRqgaoIi1ysGKmtI4GF6R
b1NdQDGW7G41RXpakbJJCJKEE0nLIL99vsNtd17yXn0BZ31sWcWmCbpX9z+He0SboMc0DvdsRKw4
b7iFC0SX9m5Yf6Z+1Dr3tKc0UArNmXJ9Q86POWIcuwzK63QunglwROfvsWZQ4sku8GOpLWGfKuaG
VP/qXaT5U0WDtk3SXiqlgsPrJQgAs5xQVx9G7sye/r9S67getoIQncGyLny6Lxk3+Sv45T7niTQB
8HPeEz5E/Y6Mp/dlPO+cE5bdbVZEk+yFWW5k+q+fKSqHOCAVunz9C145+lQ7ql0z73Bytuxuq1VN
aE6ZzkqNfij+diywcVhbOPWku6u3pq/S10TG/DNOcBjHLX2Aw0t4fodtZtEa6c4TQvfWXABCcv81
XLHAbjfUTNTDKdzK0WxyvGlwHMzG54g8SxdmtMgbT785KOFyaepB2VhDJPxFirGods/icAAdjEcs
ym5rCKKrYwWM2V1KR0x1n9BRnpuknXwUBoW+ezrD+2eUnUX2QEqe+lSbQp4SVuo5vMCpeAoBJ+KD
dUnHqX2hyRucs7xNVMV+NXWB/dxZvAHP31gcTMRXB7ZKKmaJU0gv5G4r6JpxDbdKGKUaH9N6JiNu
s2hJLnIIjc1ExxeioR01Kjxq1uoNrfLPjpCt6/uEopj9j6FPt2kxSFQWj09yHfjp+82U8Z6WK79d
E7Zt0Iks9+eXFKqrIU2ZqMwsTbSZWx2C06QFFj5+S655VgM4VX7VmtDwRuLW6jdmGMNZguGK+Pg6
gL7aOU3cZMOidFbfMvEfVrV5Pynfi4tx4bvCNtPcWcvkpN/MKwHgqcj2ltDpOvI9ChjeEhgo4ALo
TETU09zuSdWuOJejUjIg4Jt/zgKcSpkiOo7XkOUdF6jDMRJHA+GNoEqz1Cfbgq/ev5uaGpJv7wTS
BKVv12vsUcfPBQvt09biVi8AfBtPadjzgxgwTJbVv4fP+RXW2HLLDsU/xxW5XTcuR72q5wou/xhn
9EjEakcZu1PDxsjG86xRV9b+FQyh6N6DX3JpNq/x1ep6JTU5xbrjHyCSnTIZYl+gZg2tXa/S2jt2
uMtaxjx4Cm/f6LQhqmwdS5WVIvxp07jwJNO0OAn8mGY0sdAitT5LkiVPyWJxA+9R8j3/AsqAzZGr
H4QChi1sE1SVHCX65vunsX4HoK+0vVOwyoKP7BiZZfoSemrXPzjA5ccVogemPwsqDnZJLXCZqz0J
7iF5/Hgk7J3YimQBAH/RVyD+x49NYWOmLqSUpnq0+JieM+oP4PoH9UWL5MuqE2YSfbhvY49CBOdD
rzabHAOyAhTZtfqV6AFAVRuBqaf/2keutARlGwoEp/Ck0jXWdovidxF8bwsS6s3Yi2i66Y/fkW8u
Sy6H7m9gIBSsy2eskY89MGgTnlFXM3TgNCdSJ9l00m2HKcish9vgqEmPvZCtsnrBdKDld9NIBFL/
gepXbldz4j8la6Z36Eip2CYPPo3lH0y2YY91OYBYnRT2YPDcYhXvHlwNFjpQaIRIGZ5n7GtnvMZQ
FWKD233kvTQw5VlEgkCB7pZpMI4yPgkZy3Zu5s/y+ldNLnrwIShe/kPDJbQRl6AQ3Yl8okad9Oz5
Ju1whfX+99nZJ6Id8Lb11O3dK2nbIP43EBVuZ8uuPuVEKzUu4Lvljk/K4GGp/iIpoArn1cnNm0ol
XKFtEdyIDMyFLUabCoqkwCEA5u3aycuNi1pntGHhczZSJGyRAAclvLe/jHObwqpiQFNj1odPvDuu
IHCOAb5ul/hEolu7hfIiGzqrYUEXYhjPjxgEyowScpuNE1GAjWFQqXbiAJOu3XzW4Rb80QbIHRSj
lXs/ndfQ7n6+fNINsIOM9NHtvC1QH/9svzM/JH7Vm0Vowi/63QoGT9eKqfyYS096zZrON4+pU/YQ
gEPypji35wyqhaq+hcWvW192ZK4/ikGwuaaxVhbH2eH8ygRO/SKloyjmzDsa/7/S3X6zzd4vRPgy
H1ppFd0eY9iACUcAOVQh6P8IM7SOh30Ph26rkChzKfihJHpwGK0G7pWIBYOFCG3l0l0ZKpCZmbgT
2jbuV+p7aLsGGyK7eIH12FCJl7qy4hQw9gkzB1WXjg7yRAu6mZnACo7++SdkWpk8Cq0G7FpQQHx4
IKPg/RKsZgLDUFmIp82js9/fOFuXS4MgJ6d0rC6ChW2XCLVRA3KzxFKgj3GDTI8a2HOfwR38YLIq
KnkQb5s3JixolyMWKru+79WBL+ZkkXnh9WpZRfnWoCBscsWC4cqV6A/bkxwFeRPz/iwOTQxyTHWs
17EqLq36gb7j6dVA3kiFgVf0FdOL8iyQ6JSMrYPCBU31WE9gFfsRF2sdLe3NB6Syzl76MMxXoUfT
CvKeVuQyE08fG6D0IF0vR0gQjT+JEoNlDOO8pmzwQr6C1N2NYzln+vPFOOo4xlYRB/mDpOr9KcqP
ztxkx/0220vp2YqiKjep1A7m3VDYM5zvLoBh7KfvIDUdljcTmzMvjZImug2lphjNV0JWZGAZHh9E
x2MbtK3UdcWxO/fNtJLlnNMXW27oIZTlXnwJ/5Ar4XxXl57A07J8qB4620VVGA5rkksKIEjMBCr3
vZj8G7zlGOFiukNjz47smjkeNhZcXkIc41dqUjMdHIQIvNI1BhJrxJCDzeolUawFOWkXfSoO5xLJ
H626feiChC6T87JIlaX1Vfc6RkJ/eg8fVAM2MuHRqLdvnlYx+fbHIzfJwHv45ZtNX/P5UClsg5fA
+aib+AHH2VEa0RHWmQtyMciax/P7w7g5Da85GH71f8EfnzmqLj7jWI9+l0TBQZFPmiKoR3OvLFHz
o02z+iKCl7b/XxFeKn1g4Jif12Q+h+6qkPFCHyR59eTZrd5yLAxYhP/TlZMprKYg+1QMSdckEdVH
twC3otfha88k9QXfJTZbEEqijl6Ci7MPX0Mom7SHngn0/nesCe8hqHC9tr1NATEvEaYP9iVuTaC2
1hSpqte67C9m+xnKsQJgaB1sgwWgY+xb/YYtZUIGPulo69hiutwelPIqr4b0xgISI6vnvWnFrt98
XS/ljmmHdfSqlwzwPfWlnGRUO90GkTEz1wubxbGdesLfS6DFvG6mvqnjeLJId5OXSBQyzk/k1z96
4ADsAphj4wIpUbP4OikGEXGzqY26n49i11wF/3hEHqfT9NZAathltL+nbkfRpCNz+3eIt74LoQvq
k1WnKTBs+1Rh+VYO4AqE0T2Wt170w8ioimkBBh+N+nk8MakaPT3uwqJ34DbgRPY8ABGRKRELI5a+
qA47+HmcTeS4m0uEXUgDZq/OUyv5IhQwN1/1kWuTa3hoF2cpOgbQJU3+UbuUO40aL1mxXYPSeYic
0vAUf4crCHNaef8HmXhmL0sYSzDoA+Cn1a9h4M3vFR1SNHgZNy1yI9uVuMA4BZv3BDxXxqvedrBq
9pbyBEK4rnsMcYlj3BQnoWYlfZfS83SaXQ1aFaoCSitJHpTzUHBgaKAndjVQwWQDLgpdQHS4RH8W
GsdrowM1LeHQA2GME4ml4XwlZmntXQif9pQ1qa8Ksrre1/TiOTKjv2+cQuWro7jtqb3sS3C9/cN2
5YaSEcUJ9EAn5NLxbLIGW1OXt1GxkYKc2ehvuSOSAoACSizlcJ0O09ddqTXJTNe/zxEPbSlJZWF8
umQaMcS7lw7wEVaZOgT4VRcPjylgSBruXRm8MSNLlZ0mcW+1YVHMHYf4ZZus5JS8JCOlV0EiUuxk
I81NFp0/DqEhWHH7qf8CWV3tV4SJ0qYI+lhHlADBWzH6NCxp3WZudCFtlwdMWLhubDX7zH8CLrM1
6By69b65C5kO2PfRKSAl3LW9peDbue1wNWshHlqYm8xhb3o22gAQTEFXU2ct1fyde4mgRUgQMdPH
ys74A6mfDqMuPMOMYeMpH6V34T+Nt2xsbMTt9cTajQ7b6G+nTy50FM/NCrRsYd14DXeJ2bBF8o7c
hokGxjbwYe07YU91pugrzap4QlTC/BSygxYhLADm8xeVoKjhRP5YlSGqVdOhKtVDF3ItadA/LHsS
ai5lD9dELEhTATN09O/6/OfgClo2AQAAs7oa1KWD7qi7dG8frZVOxWdgHbCJKDEfQuOKGxgej38j
gftwGJrFFCZr7g8lrFE5Kc/CJohaAsU2UpBRuVT07JV4+n1kxYZqEAI7klP8RygikoAABARSn7p7
yaLTz2gAROPpeWOmaX4qzIlB5tKavHSDqtdKOj1KIiyyKeG+Pyxal0yHk2ev4afwiuxWT51mDg2u
ZtBycZkE2erIZ+VqweeBzbEPJbgWyz6+JZCoD2nrAveGDNtoSQ4FWEP52UT4CqVF5Mp4y9bH6VLZ
jbkmUvHez2KaRd9m/r/iTJFA0mK8tRW/A6/wXVnyj7b2czvB1j+1T7cA+8c7HFSwJPijOutHZWCE
gtCwMBWIXtdLtmxlQpQOp9QYSpVQXoZw1X7yWiqxbHczR7XmDJymQtUPiTKZmev7uE9vQ8/lvwfw
s2MsjzxqF1iy+AvPDmIt1z78IruDHg23YPK79Kar7SNHDHysI4MuP16XbsL9N26mSIGOifkmM3c5
PWBCRKAPhTU+BtvX3AHPCaZUMh8vaoYmpEL9S7YPRrp2GUdLMiGAQi930FCxUjnDwRlkj3akA6f4
sddeAeotGLvKnSX2T7PsHNtKXhO5yeIV10+0C+qnRghc9NkaFD12dKHzT+61TNWzE2gc7SUzYs0+
H6svgM0TdozHhWDy1KLHFmGQzg40f77guUADR7G/HTLk4m3wSRHiB7cINGlclkfQjUJubzo9uhMV
jklC6p1qoagEsUS2AR/hTMtncuE0Z+pbD7sdobz9AYhAUJ6N75hV23sDin8lvmMR81ddL2k1EIir
cJCMbzHAqc9yMobsj175eSUunnykihMxEgq5GbihzW/5d93gEM0Cykc7D7z1MhQDREIHahqI/pJd
/MPHX6ADtda4S3kkDe7uujYewhQVd6MJ/oRkN2f5y+sWAg4cmjUTwZdFc0JzSDtIJXll17nDMVUE
3GXhykn+S/DOxIIZFyVGQP/Ip4nxZ4Z8dM7i394806Bcbz+/Gta2fPpQ7Dr90YciPimyFQAV7Mud
3geKck88L3ZpJE+Rk3MySUq7c2VbS6EhF8bmXfyLmhMBlepNJhEs96jqpEm2a3WJgFC7JSric8Tw
Cil+5A+YN9OtK0FH2IpTSgrhqa8fVmZsiPpXotoF4PyUQWgU9D0YUVBflsvbIdXvlN6fe/J3W+kW
D0s287fTxlnbfIRqssCpjHdHfUFfm5gdOIiJTik4eBm61pDnxd4+mLaSV4P/h2ggYFdRyRgnTket
JDifQeiKw8nOeWffznwrKDZ9ryKMKXVFWYiyE3smLB8f4ClUiT673V9ynEhp3OQ0zaVf6f2Cqo7I
WGWSGFJe6SNUf9CAo7Qav0EOn6yOu/9rI2dZwh/5on8KKmwT6A9YLD/ud8F7NNxBKFOIbNDjX//A
3SMiGHKGAPZ6VuuX+y9wPcrcjX2zJY0nAz452siPHJ9pX+FAkS5pwDy5O2y8Mb7i02bYc9oBuoXr
CBszzu+nxQNt3iK51bkigXbuJ4MVocIUVkZJOBIqoku1Le1D2Pd/TG7VTHEgZDxgr3CmR/uU8oXK
q294oMSw/mV8XUismfCMD7dAoYFDZCYIWdJuYQ9wLUq454Tz8ZuztlFBUjEyaa+ZC+yIJQBribSZ
9RA6vuIwyYssmQDZW58r+zhW3nwEja5CvAaOwdz4tFxOZIAzkFfaBhlNbMOgpBYDFUCbgZp2S+kP
5UqZ09n5KqV1L8pT4+ZyUFwX1Fs17GCoPtw4ohqLPcm4Kj4TezqzwXu1ZY5j2xcEIXwmtlz1VUSM
bh3Ow5speNJ3DWzPPslj1pmBw1AlkqxE/O2KAgBtbcOlMdUWvxjRwcv2MCrU0MYzH+ofdnBgieVs
Z9aGkzAWurkuuXQ7YbAiqIbIStyOaXye3MtdQjW/eu/mq284VKvbQre7DMBr9C+WEgHi9X7FmzB1
kZnix9VGI1TpXmtuQz/SKPZlIVUZwrwlEsUVIDPcngD1UZr2lpOLMW/U+WeZw7pVktQi+WfSERQ4
8C0J9jXQXb/756IGF1I+EWeT0l0ewKEGPtNR43aUWL0vThS0mqvlffZla++ZXWFv8i2a6AFI/5TT
L+d9r2Kozrv6pCk3Q9cdrTLP9BMlDwClcyS/eBa7N907dvbJFhApzysPoq5pW05NO1sH2ACxKl2r
wmQ7rFO88t3HGj6dupKz8PVE1UFh8cLbFQWiNXC35vu+E0TtxCgNdqNW4HRtA2ilNAiQNI4EHCXH
M7LW/FpcaxCNTX7vv3kSGiFre8Z3Ww4vlxG3xGxZXb/aUZJUJj3F0BTyGWPrmJalQ7Ykats2L8ZN
h6pVItOCrgcKcZxJhXiDjDpLtD4NZlyFdk6mrrF9wAMgKxHtytCroZtJpaC4BZ6ysg31BbiqyEqH
myz71BDfuaGP1G6ntuhhSTaqlsGRfhw/bIymKjqdlBILDpSIBNilruawfWVe/CouRNBeYEj8UDke
AZ3ugwLDp3AVbnoupRu6/1REZY3kHpSbuzcCvJiJ7YVJa4bXf8DBCG6xvjJqo+l+mUZ9TOx8vwna
PDoFgKeReh5fVrG/rYEK34J6JFf3i5pz7k6K/q4CW0mjIqIOssikQvClHjECv0C8ZtBl2B6Yv/oT
CJvYEFqicX/5K/wzMsJF1XxbaCzJbNWbe6Rn7HFegXAsClJYnnq4vMKfXs+0pwrnzNZYzZdth5I0
EHAviWYCV4RrPNz4uvgnOZNGobuzjx+LIDzAm1ohPbsrDmzfoMaCtyj5cgPYkuc6F9FbiW+uiI2w
l6cS5YGGeZjmabeqaRMBlI25wKhO7IcrblbNR+3l8N+DiBaQ6Iz+XnVpz5tHsUFV5Vy2d41CI+hg
ZHATPjoRUV4Bzt7ljR7yejNjyxG13jPw/njb+IwXWFuwr/Uko60SfK/rXA3qpEzUnpAsLI9vF1F0
0MRHg7fcT1GayIG9mBHAiNtECtq0G5tvaXy+n+QqkIyaoT89cl02/qJpMdyb4wSWT13jQeZOTTwS
kuwQuMRkvUnvyUw03FdKa7u3tVuHVikJ2MQ/V7AviGLVHIP6Ayp2jjPaZiTsu05B/D/tPyHdG3Vc
ZwlN1JUzdjE9SASsGjXTuwWmOl9gwtWqoZ4863F8iI5ghRz5OJPumBXxGQ8lkTo5N/AEsJf0EGdX
7F4HrgjUORf4zIvuH0vILp0wNRE9exWaj/S68C9CQol6MOZkhEGgC6kzAAQOFrZRhCWkuwKgVFEQ
HQ/qYDIBG8uZY63GNq5FQZHoJxacksveXl4X/cnk+3Svu5q/kCjWRw5ISJ/XH3kpKUs8BaqrXQuK
AaAA06kRhexjqy0EJQTuSQaKShMwgz1MYobEbjbqIs+/+qnUMvWAL5KeH1kbobEyoBPTdDpDvVbM
pULS4bEf+L0yYDTSPqm3gOg6QD8dCwsiuyl8b2pxN9J5GHNPediWBQVdMGZmNbozpaNzs4tN6qkL
D9Kt8x8gPihCtu/RjtNPtZ/2qVREWhK0WggVNyfwnjj5gaS/HUqHUBTfd2SLNcdv4OTcXEHWoH/p
+Ch1il74YSB0N3CL05SOF8M9NguABsJs7MlKT53FO63B0hiHK16y2NPtmyjXW3v8Pk4IdN14ZzjJ
EyHJNHnAKjkJtiU9ba+LM2cYzp3WpTcTOf6UNrenPPl3r/gXLxYr26Hoq8SAuhX+P31SKfFYStRW
0oMn2aCueehycRRtE1sJO75AYXi/cYDv+G5HytRDl0vDenymtLYHApwbj9sEJT1GXPQZ8Ry6LtCV
VePx6HFIsYYBVHpG2gwAfLfi5gXELn/TQEUtJDHQywU60bu7vAyvqwvVT4bvYfJYYXNmKi2Gn++t
fCtcHqcZZ19WjI/vYs7f2RZSrsfS3tFpBIDRVUZ4AZhFxlR8RqgREFgtcJXyMRoIPubY1XgugcSj
YoGVOJcaGvx4q8GQP2173qvO5yo6eYq3AhmKxivfvBZPf1YVtOGyXAOwKPUXvM3yqcsffbpxB06Q
MOPuPaKDXBDgcEbgpjm4g5uL7rhL2VlYucDsS8iLZjW5DFUBzME5y80vAHFYlNR4t6ODoFhyB+Nk
4Ck0SpqOhI1NbFiPVOMk5lpyibA9aP00IfQlPzcPKIiSpej392f0mMFfErBGxtWPnj00HFGuZ8sF
829/KL/XyW1HlSwMUmsC9Ew8z2JKyyz/OVJdhGI/cr2Oi1FNumoQg/LvqQGZLvSwj13cq0ATzftu
IISwpPwagKDILeTxQLJjAHjOgk/c6SNefbP8zcs7q2ILaUBRjSp9HkDf6Cq7+dbHPrPIjoZ73LAG
86N7qPiYMMloVclVUKC5a5yn3J3BRoAvbgqL6q72TdAf6wbKShPsjhnJ4ZOV3+vtQsyXIX4RLW+A
daCOd710tZsIl/Z0TfnMJz9tFtIHH9lgm/KVGYVgguUVMgn32rlD9dOq4a4yLzTZCic1rIruRQmE
0iPShlTnCtC4HEepmOWyQiu7PLX+v8n9bjR6LamVB0kRhmgZRa+7igmw/VW7lFNGsntrhEsg8GlT
Ckk5lm+IBzAuY7QaXIDmfP0Mu0ESq/B9tPtCj92Sjc2FBA3ho4UUvRpcIiVIy66+AkK05K09ET40
MPckmtmCeIO+jdOS97OdxhDm4GbdN0Axjpff9NHNZwOLi5fiHCvhNQroOkBj7wgIiLXxZmAnB28v
Pyz392xUpjvl919/Arb7i83795Zj0lX5yzI/cwIb1u76iYKrMjIpRNAHuIyMsRECLpgMTFwJJwBR
l80PNvdwL09saOzkJHY7D7pNpmEPBSyGNwJpjDNsxv5dSKFC+iTJNaGDsoenJ9E5jX2hFzHuIWyb
P88xySfOBQXZufAKdSoO7PyHWDAHVcmKZbB6Jh/1D3RyuZoSjvBECvXvxNiQHGYwSU3bCu3SrzBU
DXs7sKYicue/71Oo/DiFhNGCEiOo8BOsG6ZsfatpcailpdrTTPlnwE6oZaUaIcAjTZWzHzYadhoO
xqiLcqQOSGGSwQg5Nd9Q0Zyd3sin89mf3JoXTtXtMqqQEFUKJtMI6Ynx/uHPhArGQ/0wB2KuSbkt
HBGycVXUtr7/+2dA++l8ZpWEwvKzoc13KlwKTAXY1dgFnQRCGq43XsrsgdkqRnViIHVYum3UqAbV
o70al5Omw1ZayUdUfd8eIo+W5lsKYuvj+g+AYKrqjGBV/RR7nEp2x/ixDxUg7AGgScj9CLOsCEGk
QkBvGnH0LK4ZWZspFM3P4iGv/glEqmWaCI0o+zmyXudzSSH9kM2vmlqbAJU4gcah4dQGeRNhOle1
lefBv9lteH6KcXIyU34+w+1PWM3EFIijdMROk7gUAwRDQ/6n70vrfIy4SWzk4EybVLF4RSVPGOcG
Qz7aI4+uacBFim6X40BwMEAXYsrOEFEuG7On6jCIhcg7BypfUSTiEGIZmdFTC9LLc2H+G3umUT1H
sQEYNMtxzUWVxs4Wt/ZaScAmxkfFFKAwEnWgSTD3g3iqjENVFe/31irkmirQFaHQ0jrwDFmyOPIB
PT7aMx769Tl5IYQ5/kIY4doTAc8OTCnrgI6FKj804h+mkBTLrBS6JcnylU5lE3ekWhmPGcqndTZd
zWC4vUdqfdcfGb4b4tRe/AP2XK9fe4INWGn/xOj3iyFkH/If+nLv5OnWNcVoom/h9GyXyeDLAnwX
++kTQ7p4z8crr4TPVgWWvMAufxbAk9lnHfHhmfwO9IkY5camCXhusQ3KZwPWKvLi0XDiC+5/7sr3
IW/ZdUMWl+rYL4jH5h+mCDoNV2+PHT+Iyv+hgPJxxUi+aYLYBo43ZRStjUAfHdCEDE05jAyvdUA8
uW84LAuE707FsM4o7+kyTqsqHCgXvNKq2sCHKIVv6HsH+eUwuZT8MvLU+3aehFDnonOE0NeIm0Lt
k9LVhExLASCWHLjcEOOwJMxcp06SlicsX8hLjGqMY0hN0l8pX9vyuV528uizptMxkQd8Sv+aMjfs
23SNnWECNQQtSiOfl3b2lvU3qKylm9R8kchvOOh/Ce4w9egfbCG5OFh7tsgA1NuAZYPykxINb5f+
bWcizAkRSMMETmDAuWINl/QaJx0XcRiKBVhlcWRvsj2P491z6wuc56SvZN1TNMB1z6OMUYgyndx0
3znHutmUeFx7j9o47vhfw3GrCOJBFQ8omY48mR1Nnf+uolVh4QsOXS3jgAwS0YND+Uo3256Jafxj
0zlSaUrpSi55tafczXZK+fNKQPV7mlCLrW9+hDmXf8SaQUoIHTrCXUxQYQR5qPdvQ7OG6ijA1Cv1
5S/k9Cahb2bja87H6HBK7u0LVtNiO3tQN/T6EeIK+vfRDNdi8M3nKMPsfqNitN0mH+4boykJ2aJF
GD8BNUIgR7Yqu3ywbVzQXxP7qbzdNC4gvV3W0DrDLOFfa+dZwvUSMgjvTdMLr4RKElzxuRgUnsSZ
WTugOePhcUIsQLTWcNPReq2P6tMS0EcPwYPIc75+S130pzw0e2llCJfdLM5ZQNZB9bCADnFneooo
amQsNIMo+wGhPse0cYot2ohzubDtx5ukRBV6t9lZrNDv41A16tn75LnovFOuWSg3YZCEo8xq3Ywc
AufdGOXKPAYGKP6+XsTBKz6H3ABBgxoG9XGxjBgFAqClDluRDMeuqLeeYvYWdDP/IRLK/NpSLTXu
SfQZ4h27L0bZSeECOzryc2Za6AiVa0OPWCfA7kj5vGMa/HxImopxnwh1wTXcFKhoQYAmTuh4W3vm
F3S7+vXGElMaF4pfv6ov0jvQ9Fn+flQQ2gWO7CPaikSs82/kMViXx7HlnLZr3ee1PN7quTPl93dO
cejj2KigOPCiyqjYARy2VSJBJPFV5KhuGJvYSQxTzSAnbGATEzDMUIysSyFFJVr0/TLR8jH3gtbj
mdP4rsq/2WSfetkYCf9qtdPEM0P07OS9H4m4hDeV/SnSUHn7mlOei8kFAtnHByExtzHKNgTJf+SQ
sWOXABik51lQJXeSGx89oqVwaNCvEJMt4Q5rEmp1mDyweZWo4i3m5W3fMr7ay7FLgfXLvB6ekXUc
1BeAgCUxwGEmadLAO24KT7QwdiZkzLoswvJ40Er8PFKWvb0Jg1K7z3xPViVu/LmZyNzfq5gXsI6Q
dMhwpZr89iYtMNYBIxj5oWmjscKKjG+LdTY9XMznq5tk299T9irojPv+qx7VsURgK7gsCyGunJ4j
dnybwCrwRId082pddqeu4uyWPxlvrzcnILwTgk017JaAAXw1AZmUXiMpmEeZU6lNmZuxgceSmFTm
w+8aogVXtGnxKiVeyoKcvtF1s1IgyisQTMpCI/mWzVaL4ib9nxx8bDqc5TFUDYB3dYa4TES/qr1/
2CpG1lR6S9ogc3PS5nXDkvAEDNz6KZP3dbetsRRzyn+rezGAEyP+VkRHyOEXte0OmXU4fgd9DP36
9T/II0xtRM1J+c0x7TG+6YpVxl9Tm7RryaX5QcpqO4aFGVRaATK2DXArx+hRnQhT5GV3KhIeAAHG
kT1WQrF79fkLS1jGF1tLB5s/eUI44ibK/d9kPP2225SbsNihLTNoBLoRU0BonM40EMHqj80wSJlh
ZtiZiCNNoSBV/GGMfenEYKljm6ULYHZo2LbNO3xMxSpEk0/Ro3d4jGZnDMu0exz5O3aNKjlwkaWt
Gde22PXic0MCtRJHjr8UWX1tnOTCo9H+k0G0wCZw4kzFL3XQ85cYx6CtkGMq//CSsEZj7LuoxNNr
8CoUiw56ZwRs1UmPZhIcOP49fmg3JoVu0u85veas0KOcAzJm4bOOtYzOn0m2VgO/c5k6FjvUE6kU
qCFQWLa/LufvnBlDzEdF6eYysrlY54C44iKAIl4lo5ii03I5q/8iA3KONESYESv/Lf2b+W0lGpbT
fcwxGSXSpqJF+Lk16JIDVQlnkbGHyRq44LWAAO8Z6rzNqIOqXaBUZgklxHn8ClQpxpkGRlmGWrJG
uC3U5WJfv+E8tsQDUD2S5S6bYB1lJiNhj1PuOGAqEXJbvB6XzH+R1gBWctHCwl88DroQSsiNMpc0
j2r1rdSukaK6Tbn4LI/w0yIUdy7c+Q+QUCJLkSmV8ebVCAJOe1uEH1jW5iw7oziKPckCstKQxZXC
JUlpOxEjIkwsXjXwx3Rjr1NxGuedek87UyJUggI9OHK/gFnqEQ78YsQlD1xZfH3g39aq3qdS1C5Z
kuEVHigU1D35yNazoNDTxx24Z4xARUgHUlY/7xEMg2FmBVr+199bVQohQ/PMK2cO+yHTcPTmqTGP
NDcJ4vjWutOpVKZztxkf2KdT4FUOJowbaJOdXhKmiY2L1YZtz9KCOmm4KiI7q199KiZpLBAsFUoD
lrE1SdFSNcJlLhTAsdN5Iote/MQU7q+8CGze7JoaXzTu/dcfGvVhJaR9BsEvAq7rgJAOrYMr4paz
ij3rGsVKv9Hbf/ks8v0D4wX1Vi/ombEfD4ADELyGwojiuZ3thtiLGj7oJ6WiuUIMIWnhsEORocas
XsA4pyBybDNeclRdaM2uHt7yTVgOuWX2w2vwikUGGQT9sIXr8ZL3Q+VJD927q49lhzjaCpEfQDWp
GxRAMNGK8YM4ZeimaYesmV4N1GWW18+gOb3qqEJDOG68VIRF/cTApLK1jNXwkfBvJ0XIoCDNH7U4
+kxbqdu8wt9XIUgXI5AtC/vwqKEGLmRQVfyGzXYd6Z+ogprLf3fFukmwUvioBSaKMTOYIC26GABK
qNQcNutIcMdPGqaH1cBUY8fCl4tNnMYjcwKVcRWPA6BIs5EAtGkLVjvQZzA28vFmXFw/9wh+AEM1
qaw1yOd4EPlSZMSFv8RacC/nRWDO/Rnr9rd1SktSqz6dGyxxceE6+ugczq5YczXT6SFNzC5y1Hd1
UVMwjERpLjlXuq7+iEIWRqeqbNcVph91A1HMkRczZK1MOqEiF07bf/gJiG+HHJ25KSZt3PPif2A/
tL0KVmwRtFaj/mjEeLtn8V2Hc/v6wjnB5tVezkYE2wGMdQ5+dnDUqsSitfBCdua2tYcE0jzbG6QQ
O0HjmeZNW1CdZrnF5wRUtgZEKtJnuVzC3RgZu4SudGyIahclAINR1aCb7CKEc4o5/RqaZIsSAqOy
G/rDudw0lG6diQ3WC9Kue+xd0AugWMeD5pr46w2kYzo7xVZs1eVgmWl3ZAxtCKyMnZI6cI5MWh0i
O5NUd4Nhz7DH5ED4yW+w0C7g0KuNkbJ47yBsJ+b1c5G6ptLyvzMMgfpfCqb3bDvYM5EfjwcOdRo1
yfDdGIY3+2pOQB4c9aSTHJ88FvqgoVH1sZWyDRz7Y9S8wswHyZ7kx8qwPf2SzrWtd4Vlb9MYlSgT
flqxHFZIVjDt+gnLsVQmsYlDvTfb1j3G/bT0aHVOTyeNorz8tUxoiJ4KtctfDK7tyLmm74WymPho
5B1zlpViV3LEJQgrA/9IK1oqt2fONmShfwCV2ISNrAftBzstinW8+qHP3jo2XGsJrkBsDE0ZNiAk
ZJ/agkJhOjf2dIaqRt77lT0z257pGkLjiZvU6e9o71HFC7X7BENrJH3X5//0Q16yaQ8xm8QJUosm
50We1at3sCoSiejBIwZqXJZJ8gruPQQ5MD4sXUs0nnlW9k2s1NBrrM/sCXv80zWU4Dzn70fNRZwX
P+Skr1XP1SphIYutwuJdWA8t796p7Xz5er/W1bjX42dcR/MnykMsDoxePlSi4Fp6hYqaBetI49bx
+4NekfXav/3waLyXz8RNUOUdJ0XKvnR7BFa4UYG26BDK7W6Ol0SwMv0ULd81S1C9nMejurUoVj+C
+aL63+hlUS6dWgzVSUDt9yN0baNkl/zZQee5W12NBBahvxPlaMkyZneZ6WcPcf16zj/0tp4Cepxd
56WDXXgKeVvsDmHAu/w/4yv5/bWD+zfxulogxtjNXJkNNXSPyc1GINafiIJ2rDtuy5E78ugplsGk
J8oZRbp3px0mSidkME62GBI8pD6fqK93puhOAuf96RA0oBg6ZwA0bdRaUV5FYqLhHcU/ZEgG4WeR
XqF4dvf9Bh6/pLK1JwZFgAOXTW/ds14SVYoWSBeL88EQlexnSZ70BCUce+X6670GT2AL/bT4+Ixy
vB2NXTgnt3luTyHLC4eF5rWtpOimMOP5GAwN90watfchu/sQNcrN6SctO52QJc1zi3pBEM2Bf27M
sSZKdC3l0kak6rfaE0b+EBVX7+CTgf47eldrIaSBafsuf8IynbliOJB9cTSMH4zXcYB0v7MX5Vzx
2InRMkXHrKETUwOXWibcJSPj5RurMpgNOrj61RmSHtmoTnuSBSHf6fxxBFoCpd24y8jUsAVPuTNU
d/3dJc+VWhacWtVdzrnIPNLqqByKY38bI+IQFd7rofY1lUQRJtj2RLdJoqMMU6DOLA/gVxf2gy5J
0C53MNr6mB/w94TVrMBZkdDrylqWCKhOZ0b4VVg9Wp4X5H7ejgP6AlCPriw2NvexAxNtp/F9o6xj
fz6hcwordgEMZLmaGBjIG/rXSQyi6nSPTJtmdBNJlkcBKnpCHYJuqSFaZTZ9UHyengL4BE23+muy
9kTbvSXyLh0QJ+uWMvhB4WMIx8u8TeWkCSb28r0M1c7gWLqZSuqGRWB+rOgzhEuuiuUsqHiYzUKh
t48bX13Jugho9HYOUgkAq5T5BX1er+X/r3vVAW2j3sGzShYe6SQbnFLZNFlMW2ObfYNrOAd9StaL
0PR1q820hKqML3KHEFKOWK4QQq4jzGDUcMkELolnpIaigfVCorqM+beu86gNTrY0kyvLpS3qTLEF
8Rcxph6pdZud6x7O9mihSPmhlVXiGtHwaJ+TkFCvhyuV8tyEs/WKfkqgB/sqHTcQu0cCJXowsgav
V7HlOiNYkAeotQly80HI92dCjbT3MG45GUPdXrHS/nAsMPt12yGn0Ey+W7NIrDDeRFXwcAVaLbEq
0dGVK63UN6qagGLviizrces1cUMSmuB08G/7nWSTsVUYAGul82LS52wVxUO7gMRxcdKWGLRaHPJN
dEI+dyltFlEWnLW4ylQljag3fZSecxXLxLn8hsUcFwb+7QyLFKXKOSowyBUCYHUfv2PuJp7jctcz
cgoxUhEoQBzLhX75YoO0Sf0AuYWzlVzAnA+pPyK2lbo4LqewdO93HYMYTXXj/Fwar+oeUNu3AgTe
58xyojA6W4bioqpK81XPLc9caBZoeQHQlws8K4hujyXz+TCpcQjOLt03Bfh0SSf3G7fXcSPVlgKk
MkfndaOb3623Ex482BpW0SAnWpiAKkGyVcqBS+HCGuVB+WCyB+p+RViKgLJ1MZG3J9p/zWWsjZ7K
6H8+I+ha3QRi2tyx7vYEDrHjQ59O5BfNaoziBaKrdbDyBUsgQiEKPdchZn8AX+dSeJjwW8SpwcsF
QFGA/EkRMCRA6gP3Q6G7DiF6NO2gqGowM1/cWYWKLYD8JO85rnEEroOnq3ggpwNLjxQ5BcV/OgR5
KBDIWTi/CoHf+liwfvBYtiV1VMo6d5MXwjL7ktH2N/oAy5yHh8Gfo9lSCCZYwUEBGN+IXBOoBIub
hTwB9ADWGSyrGsrHrLzRwjmHYEN/hJhaAyoUH/i953xPBHSrdF0ivPsrHU4mEo/jgywbeYmL22OI
ksIotKgv1AyRVkGkDLuGTy2r3Uu4Jhqu6CkWRlLOUsYoGCWJMWtxsVtGlUwvmUgB/KtEjsYpIfgf
LMqXINN+Vw4yo5+/S40TDVofGbyN3FUuiRCTmGo9WPT6JrFCE4sTdOgVgeVZpwExVZKLj8JZN9VA
Lg/7l4vpH14z6Ph7d1TrF/Qcvy+EqOqDU+hZXYh2ELDzlEi44P3cis3fGL2bLuC1XtnMzo0PHa0e
ZAuQOgf2R94zDnVg9fG1Vb+Ee/rXysylCGREmQYDUbg/h2EWKmyL/09wI7+7X+JYw3ALyxH9A6Xf
20XgdodeB8XDPN2ijWgzV4tG+8tmcAb/RDIhhOnNduxlTe9vjqZtpcWLWBPXNSbAdMo5Z0OhvaQh
PKowKhDGQa1ViLGWLwtw3qw2/0sz/RCrEaqOlOvsmlbJWx1Q0allQSD7MY4IDAOtKctU1iUuyghL
iDfvWbjMs7l8yx46Pz82ogCCAOLwc3IX3RUzIt2hrBXDTsbdO4j/aAxAwxRyUxJywNgFz0uS64lM
lcq+B5/HTfxYm8O6LQHi6q1xgF5hhGwyEeFpkL/gUC+xz4I13IxeJWuBDMKLovlcfCXCdxcIkQU8
Y6B/tsddgmtxsnfZbZkS0/PfTcTXoN6we/BdROjCLivX96z0TmgkPeu5IzUpq8dLo1XSZkN5kduQ
vuSCyudCI8Q26eOW/SR1Fu8gkcjmGLpb18MPZg6UCHiDjZTe9hIabtBuAhw1TgpAMLOLBEuqR39p
dm5PQ4IDl6qiB6zhQjnMROZpy1rsQChapCrqxtUBdjJOtiQP5kF9MH/c6O5Z0Xmq66MQMOdKHkcW
wCHtexd2NbJUk3QV1/KWGUbbL2gpexGMKCMEYD9gJQGYSGCKo6qKaoJOxik1UIfb3KetL5E64X/9
amYHnqHrAE7GOhFSHfwXl9ywHmtdbhPXmINhpW3z0NTF+TvyuPSJm20abRi8dmxvAaAxedJXnpNg
9c81r0sVeOuMDaFhS3i2ce2ycOtQhHAPygylUfQLIE0vvMGSTqxSIpEiqMgfsMI3+d/JI1PcSgU0
+l7XolpZzEQ1G9FFCdONxr85XvwmXLjdgGjoFjs1QeEUDh/GIe9xp0EnoWQRzrjDVBfHkDtqi+V6
kI8fVe+7vL3LucP7Pgtl31DCdxMvc89HfHg5aJYyJRYw6sQ1DxObpOg/Or+nDoXIsom+IYxEiztW
POYVFZwzC7Rkkcrg9Ev7B0xfiFigEmQP0qU/l0gPXVJTXOJr0HK5aotpRM8b6ri/Uf+nmdSq/4oo
ur1wmRP0WfRM72izCPf4XkJwIMZPnrYb0t2pfs+VcAaU3qYE3va6gHz7IN6e82t3A3qlX1D3sfA/
OElWeK3IypTLBrHTLND4GvVeALJ8moPsQMG2kSZnrwTAAESYxspVl5c0saR13c/YZQOYtIZCCTgo
V5gAJrFGXUtn3JnssFnIlGrkJLbRrQhc5+ZtudjeACYR+TYTQHSq8uzWG4w6WB+in0ROS96y65hI
cpcWPYhbQVDyraI62RfCuWyvrH56+4CxZg/2Ba/ZBuSBXmIJota+NvVydoQ4jAQvoJN+V2f4hBQi
oZIX4r6sU5RYoLlE5Xeyiyxop5GEuhh/f2MlhfaT1eN3pcPFJ8Pd+5YAIOszN4VGUNc3avu8hdSJ
wSJcyuKK/0BfqdGvxwlgcv8oKv5N64ChtTiXhWGULPwIh9t5FCyg6NFYDdFFZE2ybcimM6SE4n+n
nZQfxzXK/fbRJs3jXA98TTBpgqYW03eiPRLLDBLTLL2X0mBUeM1iZuK0nBD16CL7NvFYEiYnlGOj
UV5dTKe9spayPZjN/ehj/5jPELrgTI+g0nSZyceZT3NGHQl3CDo1tO4zIRhIxaRSETWuIM7OKbCV
m6LmKV+4gttwSQkBK4A3Vn7/CRYJro4rHv0puk1n8dZlrW7/w3EmXBbVYjGPDOlDrv0diFufgAin
BmCe+vKBpsRnEjLi1t8s3g0LCvNGrI/hi7KNmmC/mjNAPHC2TKEh4pp2gx2gmksne/LW8qAchAAs
Y5sgDfAcZ23DIlFsYJe64SKYG8+w0s4CVqF0Bkn0Ui9eiinzlCS+T4A0CUSjC97KAS9ZQ7ywN4cT
j+wa/TicGCPYNvanBSjkLqbdZCmdd6gnj8v81xD9ooiGfHxi1LWC7ETkIvkbFFN4nKT9uxoN2SgR
Mog3CfhrYaIvNWSH6ZYhJaqmh5Mc9JDeOEqSbdH9vvD56Xx+/dhrxY+sHnOiSqSEYjSS0nDcqj8K
CUedWRRr2yqXX8ewb3pM2U1dX5xUljFueW8/CsH7Sj2/yq5CV1gNWB3Xwo792xy8inhrwsJa2XZq
7OEbn3Onj0drDlYJwSzEIXtv4ZnDm3FRgDitnMigum570DK7u3M8g+W4karPRZkZl9djR5Z3yXdX
mVHKe5elNrAIUfTlsE0HH4hMHPVUIlewXcGvqk7iaXDQhDw7cgzOwo0oE+Fl29OxLKpVMnOu8l7J
dSHDSs1aIMcV3DAsCBLHPXcRf/t+BozwAN/3KsXuqF8W4D9NL+4XC/h+i9XpjDo5G4AKGi3hkC+m
LELmaioLhrAkasu/OSd+PdHaLT0KritDk9d7macq9TvPz73EXiJKTAGBDTVcVyNxKeixHC2jeldR
S0BFMbkKlh3qilIoX+DW/4kf1QBhZjeEWnX1JX4s7zk7I52ug8leazjSMco892n7LlD9EEX2C3Qj
biZmgTk4W3M0br/sH4zvf7hpKg61tTFubN2kjyU8rQ7HFXPxdYjV+s1Z77KWLZ7n0wMajy9ZH8co
ZbvA1ZSWBP0Lc8qcuDBjkyqkNlE8J69L3TWhW/2YjdhX++6wAPxk9ti+GGFFInuGukGvGbJpokwj
fn/YoO73al7Romzf2KyfK7QiNQ/BRXayREMGYrhw+7HYlNTpKu7xsju4RLcosW514Zc/EFMsvPZ8
ZMaIRnVaHbZk8KbTvM44+kB7kviUHvfIDXxW3g/DQiW55lHq/iTYqFRXSkS/t06F1nmHIydCIST7
77s+OVqR05SwXEetw7cLIgYotM3GAv0K1jBzmjcrJdbRRB/l8IrXlWvxWeF8ZM4IUzOxmojsAxjv
86H+5oqVtIZ06CqXBvTFqHO1GypYrM3wyUfMcKH1wIkJ8oReq6mbFnrBhDOA1Osy+7fP2/Yf3g9d
wlyQJ4j3D0sxvs5HBnF4HWBc+Vu9TEgmNSn/uY6HylYPY1a/9KEKm2p2Tt2YYgaYyoWVrbj+BTL3
N/PetMocsW4eVrTIlK4pqbxfTIFxwy7L4PI5qtw7TzUXxbSMB0KxFApRoWQOaOc1hVirO8J8nIRX
FUQ9sjB/de8kg9IxCq2Toii9Y6qXezul3pIBcAIAvfhlUZnRTaKFKXlV/qxg6uG3MJEe1BaHrPKV
uZd5baGBzm+e+yf1+dIzghfdwvFSnRUr0YZJwxEkEERQCcTambAwLb1K7trItwun1JEPPNPptItk
Jy0jY3UC8S7KR1w5c1t6V12v/UcXCblXvH5+corOOlT7fSIhyasgWxA9ics8hSpyhvNo66AXUCPH
k73o0AjS35c20Wi1HecabSeuKqYvyQgYiHoMPry0QxkiN0CRVPoBnWNJOerBIECx8Y9HXybFzTyh
RfM2YVgNN8g2owZ2LgM1H1Fa/+ma71i3oJONeP5CQxXNS6Xe0ZM8dHvDaRiLDaydXF9qEGzd0FiN
NmMX7u3QDR1gcSOI2w/R7Hab0yzjPQoLsN1Heg2GYho2HU1mIdmwG5H37E3w7PkxOWauu2hcUf2a
VldhbW2eOETnVdrNU5Tlp+/DZycuEUdHgumQNDbLXapPwRgsV4DnKb0tqxxgmdIkPoTjJU91pBJb
/7CFe2ZINVdpq3K2qQ8gbE8rLIaIz+RYEi0Z+UNpgH1Kkf27edJG2kkxvr15USwAxiT8diITUn8U
Ccjm/L5I73qy5OWd8wlyzNcTX4Wry+RDW21BQqsfg0/W5Fv52owPUoArAAiwD7Y0Z+RUnp7l5HsM
T+LtglMnq1UOZqUsOmGlHsXc20lAjaey0MeQr9sQ0WCjlPH5MmQk1kfODU6AOzrWJMxea8tvaMBd
0naAH4t00t1CHG/trmvO5c9mIbCeFOUwXoZE9IYcbM67CARZxBH7ZUBRCkSD2tA8cbVlalAKCjoR
+UVzDbQPsKsIYrL32NW0UCpA8vWaX08YfOp03hFWPju/BFjbXBMj1wu3c+J7vyOlOgaCiiozdvAK
xCJvXGc5sYfG3BBR/1MuofWRuPePtmtzNQEf9u6qL3lzWNKpGOqVzLcYUx53L+SiCIKxsDNw+wZM
6aq3TjMP5yheXhNnpIkRVyGg1ObiDrBii6KqZajjWZRelACgMk7J06CpxwiNtvuJjGs4cooIR2FN
u8MWtvcorCK4lzfHdfnrUNT5NtFBvs030DiWTTYyXyjZRlQ3EGuqO/tHV5AvjOyabUq7NLvj9MvQ
agcigAqGFlxpMLpj0MkILZyCijrq7xmCVEuXaWA4rHOLN0kK3tc7lHqiwWJQlOUKxkHRs0jiweRa
/8EuGdJ9Hn4hmkEqdv+XDx3E1+/DEh+vKRiv2gmKExKe5R6evpisod3l+8a+Y8jjDeiwm2HPOnKk
H8BFUPPqSKKeUa6X9AB/RQX3G2LHj212qsezY+snyZSK6I6hg0LooiNDLcUnZnlkr6Vn2tuggIWa
dnSxWz6zymoC5GgT0uNT3L6nt+mfDmEF3VDDlBtO17m2MGmEzhI7oQ1WqzBCqkU2fZxM5NXFSFk8
MdIxbL18ZCjs/qkhgvEiN3qvE88fC21ImGltX1XoJeo5ZRahEFigZneT50CW7ze6BtmSUyhTY4sE
QWEZQQT3a+j1r4Vg5ECBRkqcvJMbjaonSwH5cH68elJfo+1Jj9bwlRrIaSdYrdFRBevfior6FykJ
f1tAk1UZtEr2S8mjWZIDDQ33TAMn90e5cSHY4fZrqsDsKhUFuBjKUfUhzjzIgMx7IjSwesSLOfPU
Y6OQOZpfQoTaPZZPuq6aaRLideVwXMCQ7+mqzJzIig7EJTNjDhbD35+Q4hAoxj2QpGVB3M1vR97t
VU+NGGBIfUVlCHt0M6BQ2Z/xokF3HiAj6A02uZK2N6nqh/DGRR+Dpqkb1ZhbpfDtnxWQ/GpyeYNY
EpDao++V4Wd4DOUE6xTVXPVuw8LtvRDIHR4VQ6dw3KP3BfNZWPgbrYf3F77ZFLOP/mlIfKsRvd3K
pxM28hSofMw2sElutgOEfLTd9KQBVLfVFZ1RzVKEPizyDNg7+a4o1aaglof+4Oqv5aML3JsK6Sf0
eT6ddhmJi5weMHi/ThBapwxX+aiX8Xdx8+LK3L5m+MFA1xqTzqVw9yG2ixn7D6k4u87wkIIrabxt
4jTArfyW4vJ/1JbMKOPX5NgOMPzD0m2pH3NZsaBn1WqKUBIPVJjInVk8ausAk2UsWpRl4DuU2Mie
BN8Wp3tLlLtaUuEwQ4Dm3H3vNJqI1ClCJPKiUcw5JtccbvMZEzbuWhPvshaP5zyjgJ7aTL1Lwut+
lrGYIjGefkkPWCJCsS0CHrhVMLouZ2l5lNhaXLXTrbWP+2nSjClDJvJBMOzzpkJke0HFKqcUIX41
kFzzWkr716i+J+4dzKE76VaT4iH8j0LwJdQcLJ6ttqTBVnk4iK0YzTtZcZZNUaYSwpilBRHS9ip+
5Xfz1qWh5llFKsL7F/VOxAqe42mPjV27xTQ2F1mZ2TQoByzC9oc/YOGJXXoh46NcyaF2QmVqiNjc
vfiF8KprdZLMWWbi4S9EnjXPYhOLfNwFb+hyKm7Dz0OOiHH0H6tJQXAvtmWqzmImJLUWbIFit5Kn
6fVif29AmRzHepEHqgkjcJ5xi2SYZ2SDlqEgVwuvhK/IyoqlWWTbf9xisWq42vGH0drIJqBmf7n4
A7zAMI26idOOWNruLay8ZpNiEUjqmh+VIjJyC8bwmQRiQbiiwCRNtQsFvr+ydiNxe6myMgERC4AS
lS9LPAFD+oDu91CUg2V8Q07BoLA/Ft0PlD1rqAkELKVMRY14PrmF9oFSMibItnvxElgetpLxz+EL
RB5C1PtK+KbHd0iKPrN1pDcgUdL1F4AXZddkFqcvGei+8hmc0QKRgNR4Roya75wvEv7xz3YpptXS
ql1zSuCGvtegsbE0VXNZ5JxblC3uLeyaNTVkqkqDnmSSNSXkYUa63QjVarSVRz6zzOWmRBqmSFM8
10qb6bmAYNHMu1K3xPQHm09DbkjRu+fAjsZrCXl4vQO87cA5Xeezgu9iOPBO7zDb3XuG797tRCxY
nshUrR0JwSVoiYzx5F+ges4ScQShNrd5myrQrhTLZrMlxgdhyHlt1N8X1El0rkbgvk1wh3xvmfsy
g1Q9ohdL2lM8bSoqBkBPEljRdd6zUthgMHiqAdDTUS9qNPP6Ro0qKzGbd7zsidE9zLNgyCgDHJfu
7Au0J4owHuBmb6z10DVjhhlRujAzIzyrg7K07YlvBd/IWzvX30+eGTajlAoSo1C+wl9CtLTrKkLi
EdICAEq/2Sw+GEa8dhzRp45+gznEALWI1+8zfpcaAqvmZXpzJbYfXpqrjQ+jwayQzag0z5sJgQh0
+5hNbd/GJL5QWVag+CtqJ2uzJxMesw4Q09Kk8BwgRWq9vPsDCMGoQlwnQaX7l3LkKjgpRLuxsiyl
TG9uRwPmzbOa+A8mItcuaIKFA8FxsJ4CepCmCwjB00OiRSLsiQb7Fh06aXnopZtBh2KGBZ0tj72F
gE9RoK83sRCCZSQ5iCi/7dPQBIz1vsqpcZVKjaVFaYnhfOuB8uZW70EgEQCLwfANH2vZVBdrlYPH
a4iiCxlsFIr5Kxo9lhVSqsK472OY0lIubeX7Ux2AAwazv9lxoJNc6FF6GPTKFfXOCTJAB+rAmts8
8oc2YgGYPyZhStqVGnmHKX13qt8NGwv56mh7LVvy4wJSIGJv60qJ5IX5b/FjZ6iE6qaBcbCS+zQU
Z2kwoHyymv9NmHACvgByS/wU+Mf+V56pTJH7JclkH8RI/5zpMf9Ns5mIzINPkSM1JISexi+A/LvA
p0QZjXaN6thMcEGqIEirBjyz4QKPjii79WMJsz2I/Y7OdnmZHGPKbMjukpkzgzPTAlmXItfogtcC
WFU3VRnlWxRExHPWtInuNvuljBuro8M7GOsexUYEBsafuX5WBo+6zuhUSNqWZzjWqxhSV0wF2H81
iRXEI7ytho921HGoRfwosPY5wP5tTAzk7iewscObYPVxQ8x8E0zbg0jXsz6u8kHP8qGXfUsEDo7u
QL2X72bG/+7T/uzISsrd2LfkUCLF49Unr+CBT4ehs8r5YD2MWagaln28mrrQCQgxwvrTukUvFNgG
a5QVAZnPa8D4FkQ+MGzgcyYJ9P6XhpzEodsPR+u583grBbi2yQQkOyYM6hyGLgMkyzgICXdX3SDQ
54CngQu9P8gbTEhV61bWbZSiZd/kLPQVANpS3C6JDoGVIpoOlXb1ImLzlvkW86SnltTejQRWCC7j
ic+McYcbL/GaG3wIzuZoYMDZbIBv4RqwVtkrhl6CKpZ00aJxTesmAazHjlqtAeO2YjJOlX4yQy0v
W/Ye48ZaPLi85sn7+sfNsgpwNdJl5qjwdFP0La15+s6iSvWq7ik5kj9BAJ/8w42jS9YSTOe6Oi2e
qchrfEM9LMVHbQLpU39Xi+oegNDFSJHgreT04xQOLQd8jw6urcjfx5sqf/COCzpTzB+0zoMCeih0
swj+InzQhQppo/N1NJUKl8WzzAzOjFEav+AyFxUo+fmGxZBeZxYOYnbX76Fz5A6d6K1FxqCGDqX4
w9S9xwn6a9eflSmIc/Y8t2plt9O3trcCMoXJ3rS2f0To92f37FCK9hbIzJebM6tmtgUovyd9crul
uMiZYlR1tlrVD8xcJzukMIQcUxfsxA/5XgKkyJ48T8ceYxPxScmKFGY7Uu6gDpcDho9WOheEQK9r
l+Tvv3EwYyancEky0aMWGeVatwuuWuYceVi1vIGDDZZKculbz4nrmjHszSlQKblHG0/WsBlWyKtn
AgrxHqEPEHHoGy7tkwgDH6iHBXerILG1zGI6IfiKlyTXyHPq50hsY6L6CQrLaZWtnIlZgO9rches
vWiIu63FqDKERDHyJmiwlfBfOihtErpqH948ycEkUNXlo37/7ndyO+AN3W8dd1t42Uj0PNDm7VX2
xjTgc+uPl89i8/08mtbuyEGD1e1kPxQteY+0iejx6X6M+1dHSsnZtTQqF+gRMdhPpaIRzV3p3yE3
2pFV7aZCHG5Jjvxo50Ee3LhfgH/6MFNq21T3I9nCPeE83zrGgPWK+u6aMGQpqN2SrPco54LuYi7K
T3ZH8lozTDLvYrXu6xgS7TiwTE3M34TLDU5k9A0CGmZBjP69I8DG3eOboCcTTWAN8qOAdewRDw2h
oawZX2SM8QDie3B1SRyykEe8M25xyCgDqxi8k+vWbebTdP16tP3eBNsJ4xcnyIKmE/3XWtI0DGeQ
AZ4jMS/ooJM2gy4KSBiZcDDbc20urSlIIWDAmjLJmaBnCIY9+sXldAlSmiqSPry1geX4ngYTadjO
q7No+EtDpcQmcXDQkQe9XF3eDj7exCBjBTVtEMLQ4/kefgevKnXeU1iSKZzGI3W1tKQLHosL9ZFH
O4ygmjxBJ9LRk9bmonXb6A+RPSzlSrs5ixpqTb65Hr2iRUJLbO5Pe5qrckWWmPpiDzWX3Jxayycj
DuxzEXtDCClnsvsc5nFaGobqDs9ezVZXnjjzBYbBC/Q2Ph0poe8PT57bOkdjV78XyLZLQfAJVD/O
Z0YIZSjxNlF3AR/CrHbP32KaGwjTWZMZ/1leVKEDgW5p/xb9rqAzM5suLs57I8QLrv2/9hEXR1AJ
uo1sd2AdzkwPsZm/PSIFvSlEJD+EfFNI5bEOIyfLX564YUqOuYLKx2IcAqm/byiDYF3ttBNV8EBi
l8/volF5TRC8V4rnx0m7PjQnf4XYjwpdfPP2x4inh1raQTwO0fjrVZW5unCNc10eUCmi4ubckTmv
WTTBfih3iVQ7sIlDY1FgM3XorHMmwkdraDcROKbkfhVHV5VzCOHlNgPC8aicHtOj4BKuAiyYMQdy
CHOvctuTaX/FEsBoAoqu9PytEANTf7ch8Hq/opobmFxYzcD2fEu2/A4TiL53Wrvtew0JcL/NfiAW
Xs3mbefzIqNH9F/xQpULwKTxB/4yjxHr1MRfLgNKddYPzUB+T6ByAvEI1K2lUcB2RcgZPvC/oPyq
KexIO6jiJLQpfHby7/MlXKx2tyP1yv4WeZW59f+BwN1BaeKqtkr+cv7jBCJeylWGOz8GG8uL0QC4
rvhANfNthWCOUOnXacSc66Oiw0IG04wv9oeUFlya0B/VQh9WxAxTDieFzMLtvtc0h4JEvPncU51Q
i7prvZLOSoqycGlC1jxd7+ovgdKnhZ9ucsKSnpFsEqEdF7Is1vPpbYwBIDy3aamPUlUAvjwtGNbK
OJxLpcltrajZfk4QbvAKCHFDDoOHhUO8aptZFT5/ybh2i7mMpWxSgmNKMQ7BPrIbyYVb1jJfTe2t
xxFAIOwGu3qiNWSMEZ1vfT67JaVL8N2KGbvU6HFqWc7YegDXGpwmN0o/3Zz2e1uZAu1HFC6OUDR7
qnDsTWeqO39Wezn3T6JK3RDQAe5cKUG7SzN0AvCJSEf6Vfxz+oA4yEc2MZeM/5/RoEsRYBAa9u3O
vViOD1qwXsjaGj2ycAWGNfkc8Xd/7BtE3MIpFSH2SQPiplgMmWWIiFSOuOV8jO/pJrShaCmhzNqA
NRbM27AM5L/Qmka4qChFABmrBLPX14O6sNW4BbGRPOW0w+5TRMps4xu1iyOHPLegGn2eKeXAmJOe
5jsFO/K7ejHDlYLUrwmTVVhCbnC5eQ7FixMiRlDEC+Zlw9q/gqWH84IP1LEQ6JOTocR/vVDQvcru
TAtoOXrjDDgku6soNbN475yibDcWiA7XUQCEHP/huw+saNiGTGwqZbO3USSuwXQwoOidaEPejcaT
xO9pbsi2e7iiRPfIlkbGwAtbJPKuui9e4LYfReWs1s/4PMRPSL1c8CCMvsmZZ3dARfs7aouYgjcM
xUH+gOLQPJow0c6f6aeIjYTKElG3gs2++bGvR+PYp8QIRGe7KtuvMGHn6xmFR+7PrgD6qbl9pq/N
N+biTSyhZIFKsJMbWHfPwue9Td+lWDGDwzypmtr9yS2RnoLOiaNBbK2UtqpN9WNpv58jajzWHBxl
WwNbta0FCwIRv5uLLEo3ggNnfMZT35Tkroo+/TUXkcIVh5R7cvszm/ShY0ZWioWK3lVwtrUH1pz3
uC/GrCTJqaOdfxMOb7wKElYFPGE/55PPl5YlUgtaDCnutRyVxuJi3P/siaWgXcNgjL6FwSND7+s8
A19katW5XP1R08Bps99gmF7iJjeH5LzqV/MYaxSg8elFZG5JigPku0O3zo57gOeL3Va8WQ1m0NFA
YrdO+6G0k7Dzeq/7/b1vO02SOS1IWU0nfqIOR0TAyqCkfFYShBRXqwX+bl56NcBvqrDX4WE3BSUD
Q8GE7HMgE6KAStgehzV/EY1qRt/b2Dzp7bO8DfCFd5bwShFPkEBseBHAXBJJHpGNykFXsbh2NKuO
RHGRKZ92ZJ6scXydJDMKaZ84MOHujoKmSg0FU4EIqQTIM4Zn4Vl7rmLogJLsoYI6Ym30h8FOHSYc
4xOCtwaRsQTXoDDxiGjb/qCp4yeIzrjd90uof9+aWBb6pKjd2OpVPCxJnZqipWBRWi0OCzC4wP3n
0G7RQBgfCxTaxRg75szOYiBZn65WN8QXuZA1k0xOOEmRhdFIinYzQ12o6v6oHFoOHgOFtk9OTckz
JKoO/AdYW05G7FnGYAsR9AGHKyBvgYFmGhVUENm7lHaEqje6Wpavz6ezcvA5BHwvPA5Qh+XrHzIr
WWj6WPYUvmCzH3awvyMIuQsU8xYwuPPkJ2UFXvT8qVcYamU5fpXoo68Ajb3Pm8WpX339KPto9MM0
TYNH5Nx19ygCqq+6GSpnzrvkSg/bfh48qKgdOvAuFcxjNugFlD6gVqRpa361Us9oR3HvFmqEH2fn
LLBlObkldizrbbhCjIim9v8Ar8ALgrWGnF3rB/WWX4m7Vjf+iKeMjwa+4FgwNh6L/eDg+NRAwI+P
LvLT7jivzxTmR/ugI8hPkxDf3Fn+iLbNrM0l5J+f1CVFIFTxRb42lkqTV9mNVLs7Al/iG49gsnbs
bEjl0hb+78U+rZKvNl4D0v5Xp+yXrE9g2MpEJ6UK9DoUDfu3/pX7RR2DGIQGBSkQjd7d4GnSnR9r
WzepK4QehRUvRloqStU8XyuvS9NkGbt1d8OyllAB6FXXRS+K2Bm6ILkxANZmtEY7ngok12vGD4YZ
kAnsbiyYbQga8iGNkaNtEX0YCLk52MucmYT2U85CRpqsrJHnUe7rM1GGxIWJSuty/d15woPUgXO1
MBfGPYt+rURD0QtMvhdrp3xd7anQQ3+RaROz6YYi7hLhoiyr2Hcv81ZIm342f0jIvY8AYYGQj4S+
VFU78uCr39pGLzjZQ8vtFkfFB785ByHbaAM/MC4Yo3mlGyyAEzilLucllyhIOLWoybWsAbqLN1vu
Q6StB/rg8+Pgl8sxGYYpPZTuLHuJINnuD4tohpbBupna1dhdbZWJfNpyzLh5gZoHG5YhNFyqvmMQ
7kauk4S/WDB+GArWfluPR4oR845Z9YwsiPCnC3A5xmvSG9s3gSFHvmrFPveAadL6mR9AabEMzQw3
OfqKar49iLN4rJj7ryNSwKtw6UGcOjuN1hjQD819trJzOWlCTddiFVllQYF1Xs2yxv9ueBl6dNFO
7K30ppf5IZVh41DNBNk+dMMkwG5nhKFvePrZAZ2sNJw+3szoDkiiCXIdGRFUXVhIWLX8zvb+jFAU
WydJWEXxJG6adMoViMAhGcl7WYKa5gamIoqO8e/H4J9MyneF/jVrr4+QYbd7oxNSU6qgFy1IEILA
FCkBiGZcBPAMECOIU7Ub0Ex0sfoNUX/Y/zuURcNCH8uejsDklHjVyQHAyHZfmfZWfrcYRYydjPMj
Vn2va0ADtR56AlvsP4Afw1PN547tbHMKp/DmPUlf8qGiC7feQxpOYGr18jyNOEXIt1xF2588voV4
rdxHpDdHNfWbAw8X+bYz9p3k4Aem3MTfFK+3pyNJNPQZuTAC1zlABCvzJNk0YIwtCvzPAnUEgkxG
hutA0a/uhn2UjMblwuifesG2RLNfI9vSCPLBXCIIU8Gfgc6citwwXFq+Pegt6IMEKfzRW3E1rDmg
996fMQrlEVTE9Dx2Yvi/mVt8zivxnwJBi/lnnkAQDhQGpbjB353E1euJfalCBBPkbxqIuDKofJpe
Znzj1eUZNgpVSO+nxnPB6S+uRSGJIiiJSn70TEvfHB23MIA0LwboUgLrxwGS8nsL3VqwSh6IAOU2
V9yuTH3qGh1IcD8ghIxChEHbQf+aKz5ZAm4y6rSrHTW9OpGCseZX/JH8sVYI4QW3hB0mUD0YwJ9t
O2JPQjVcB7o9RLa6AqrHid6DyJI4aYvaN01SnffApIgKfmrmanKete4P9r/wwaKi1TZ/O7Q8Gq3i
TS7DIPQm5Mx2yTf+GpJjmRXWcOoTr9hBtjZDoSr6IYCz8vgmidYq9ChFVIzY5pNWo33/nl7vF2iu
EjA9897uEx5fXgpoUOpaIvUJymrQQdvjoQzLLx7HFeHiIDlJipl31YV+s94lJ3lFdp0Qa51/AqhA
zWsdXQGV2Wd4+gUD9APU5a/FHx/NO0xdCqApL5GNi0xWkdiOWdK1tVwGSZOE8lKmh7fiKpfEFF0p
oaNIAFhueutYZdEPuhINi57YzdckbCXFjX2+DMKitfzEjmgWOvHHDBNCr9HsT1AevbHIfVFIe1VL
yIJfDtMB1S8h8m5YTfRAMcww834BLJKD74PZHt/c3P5Xd+UB3YJt6kM6FiXgXimjC9GNudaAKk4+
U3roBs/GXdj3DQCvzr5Bv643AYjbZaie9dGA53TIqkaq4R2snGIoyL1I9MAMhcC82n46ptsIQFgK
0PxlaV8cB5UGeRPakH+gXk4g9n1wiOZLr0jMHK7denDA9Nlj2EitURcCwKonnzNN5UCK1C9sH2d9
3aDhoRsZ3SYpTlvb/Jrwkt+cQO9DWieDgOG58sUFLlssUEnFhV6f2uqb1TQIZ1Yi4cdcNggtJKQH
OSeX61VqCebgxGSw2+I/gmh6mhCJM33TSWX0eCyeGyTmOy5wQyugXBpCSS/rYfQcIxsXs8jvZst5
1B07n0ZlsGavhiy1jRT56ytlztpU1UbS82LHQpuRUZ36nMyqQStWmbM+IiimL+alOKPCmltrmM5X
pEvjRI27m4I5K9qwk17Nx6i4W/rvZe2fvUxf4Dw4Nmv+z4InH6cznxcWh5rFC/ie+mr9A+gJ3tlw
MW5jAJdTAZl4WO7TFLwBxIeWGHa8vHXlNQNg7GvPbf4u/Vnb3VexcObR44vcog3+d7JUqm9b+f0L
h6z981u68Scefsc1+5bW/AZGO6BDqNuZjhl7h8g6GdUWFeCmjZCFXZ60x0xKFYEL8A7JwyGUATar
vKs9bJzNeU4JMrTz5AZ4osxPOTBCIMMNtgl8hjuzBo2c5rbEJq2ezqBuqpLysOBHlpxdyF1XwN/X
zMdZztZNW4LAXbQXTaIrylIM9SPikoWJK96P42eQEyOdS+PTIByExER2G6H9r2qoVer5CVnt3Knp
TQjttVoONQ4aWTji3xWNSHFOb5t9S9JZlCEaDt4pZLTXHr6Pchqj+ONKjvuUe12C+A0vNdLFZ29R
6rLeLfopeyKQtBzDAv3PRvv03JO1lZ3pw37HamJ4D7Fc+QtyDAptuOkulzwAFhaIq71FSRYGKhxC
c332oXYM0xqWF4zr6L9Rc9JikLNdrHhY7FpC5sIiiBZmRS53hdrXXy6eArbRLoV8zKTYtfuLyg9v
KXPvUHfqV0CKlVm/E55zH7Cb2yFSC8EjyNDPIJ07Tq9Cz0DHBvwmCVC0afbfLEGWFXNqvSpKC56e
PUssFEDr1pUPQZcf270X8V0NDIeQcptjKZ18C4YL0p0PdsygwBvTewJxiqS66h0mj+n8dwShhqT8
1bprAGTpPKRp4/RxNPhWzuTHVxQfvYrkk0hXcMMl/ddtSGioSLthvnMpMuql+QIExQq3ZYVxkrqQ
pzxRTs9dR0BgPl5XpV552nNqFHRvRVijdKO8GPrTYeADMiLkqFGQpk1FaYt3rYzAyrRsqFAmTXVG
XxSPmqk/1l7zMrDNCscuw/l8jV260hgQ4KF3ujy/Ivvvb18YVkcheCRRM4k5YwVebbXb4po4mCC5
9oho2MM7fo4iaCNaWTkYv1wFcNeZ3c7NVq+ju/JqA/CAGXhXpVRkB+C/FSA9dVFv8zb93HQxjPYe
A7R59ONnZoed5O94v1SAYCg+NDWvMZbT4ZAoWsiZq1+0oMM95zup/A10jG7/BnPkH3NMni8K0ctI
340tmvYNPw+H8ve4APSCTFAfGk20CxXNlUMPpl5eOFCvphsnnDFyoU/I/6G7k/Hq4O41X2kD2zKw
aRhHd9efb7CcVRWM3E8gLOa5CerPxPe+xKRJKF+LfSYGtHdqIYIApPszMouP4MSGQfsqERrRv6HS
FWeZPvv3IZRLWwiTaA40CcrAnKhdHs2Lf1P8cIgayW2B9qsZwRf/ZuxqRMpaEpfD9dEe4lhjHTzi
bz3nmwVCryvaAE+49fGQjdBbmhprxGb/wTrzemCfQWZkTkz2hjFG5tnNOdBO+TK6YSa3yYaGMUPF
yLSSzsymVv5Yr05Pbkn7+7qLIDz5GoqZs/DqhI6iGaQMEtUs2OplXimQMs6wjyGBCwCRMRhD2aZb
vy+wZ0QuS1++riqpxeCVxAjtpAqjTGFarkOdsqs3FrViG5ogsaZCevu7Ax3lKP9+pj0a7rETHUqv
+OS/KAOMXdujCz4RX9nqKdwSPpXnCmxQgsugJAtew+BcaptEFPoZn+bgv14drrSLNS435X1rRADC
RPmnULrwDDCrfvXkwBhSnTHIwmVeNPo6eOHv2FghMbM7v+zpGoInXIZn7sZ6vejzU5Amdw/fiMom
cMnYeyh0FI2C9uZBW5Lhk199dT8esS3VNc3hxUO1+JDeZwibUB3AlgGFyASR5XCkI14n7k301mkc
ApE0sJrwDphEHognfGrTpaWsaOPzA/oPIOOyQ7HODorrNWWYlUeE11jZnfVj/kjI36bxO5vATjm7
2au0Z/7yvUiCHz7FV6ZMWzIzPu7kQ9mXdwwsiekH8e/hoH/fSJ97qtjkQQG4WThWXtEhuO6B+FAS
Np2ovmXwCZLzNi4wZkB8YjTdpuRlpIwNmww4bj7ndjoPUV6cUh/tX0dDuJKpNCRD8gsqLMSAS0K7
frJAGSS5VqsWjr1V9olcLa+l8yrYZqFLJi4MWUIoc0TUdyqmgEybtndD77IaB2TAiuCfz6HrRlHE
Swm0EZ3/IhJhxMj4Gr0fgkOKeWdhoYV9loD4a9QRSh1rdA9VbQfs/bvyRFR7HjDLG3MR8UGjR3x5
3ovnPadWxqjqgY3yv9lCByz/JS3uodptvuAAZh9dmGqafJrqbzu5zneQNngviMlfMwE+E+axuTcJ
/ioQABXklQKqbDg1Q+KDiBmdRX0Ke4W6Erc5vSAtDh+P68X31CSPw/JdkxG0fFWxyHEZYLWdqE3T
sP/wqxTOLpSulSeO/9O4Lfq3IOtl8AwyGKB5XNgd5kBSMMT8yoMFyo7CqD0B8V2LmpNKHRCMVxbK
TKT4W8+v7Bg/wSq/1W8li38Cp2tLItJQJAFZW5q0nyuhJcNWwuYO7b1a23mkO3/ueMiOjJCGmld/
02s/h6mswV8gLxwr918ON2kL/3OypJfuoshyiS9dWQgHqceBF4bwdODRwyiA1oA/BABSOZ0Lbz8m
qeKvBKg+KZcYxLRArmgfFIszWbgnMUsv4cb+qJGJu3fgU6EG7oJEyoGX4Jy4FEnzsaTs96+DWi0n
JyKb/dSxiE0OZWvCVDYKcXG5K9vMBuFomTLdIb84fdXdLWlqTQWqDBBWsMC+mldB2fYc0K3WmVkH
k+7T/hmlfQgEG4amGXLZNLduMv927ekxtomBp9nA1H5XLgnTWxQ1ACsArr2dCGF3tTs3V4UnzV3z
Z2Ywg3K2qbscgkFLBvrI1DLJ/2+DA8Y+RhCIAhkbepWKjXkLWmh+GkfI+2C90iP8TNWVFbAT1Fph
sLwzGb/23BkkM2fN8Tk848GI3ZZb0COPeT+rdbG4hQb+ooxXKYTAPUOaKI698CpRZOyaKJTDILYQ
x9C2L2lxZv83xzc2IplJz37FsIIELkh6fvwACQMj5M9pwpTWWF//Z5v79SLcIvfRoWLRbpeIlcFe
XaVkHtknAjvzd0vHxApfcoqu1MGrE3uTFGQKIFFjQSm9Wdd2f9tplcHlShieaZfFM4vCUmzmXjoc
V1nuW/Lo1O6isSqIoDjNnIiZhDqVoibxzNOYIKJAnn59VR+TZ5zkD7tWHnyG3CbYfJq8kX0mvfXn
9TR5E5mp8Po/38Mvh1pCpYE2zH8QSB9NnN4o3dywCqVF4V+4VPmacRX7RkHpq5wMWASQ8QiV2JIf
MW13gSiqJzmAz40Zq0YhKUJuTuZVXVoIYZ3GqNY5vHMaDiajBtKZrS+UCFbbR/MUOKWuUb+/ZvSw
YCg5LxtU9f1tvyA5VJJaNja7JAnggRTG2mDmJIhBaphpGx+L+YWZh0WXC1iDee0nnJ2TVi8n4Uju
PyfyFrX+1i1KTfOJCx5nlsbeW8P8bWXiDFAsc6TinPZOrGkhK8uW8B2bxG947+CuTCa6OR6kQBKO
3vNhm/qsFP2Z5ttEKJ0PjVdz2po1SDO8Fnc4s7Q+hqXPnNeTyd4wdDYZE7YXRLLNeqD0AaFnuu9S
dMe0fAdKC9ka+1CHcWI6DWLcVAzm4lGz5AAag9bgxYmnS7mhIay9M5FGadPSrxtiLP4MbQLB6Xze
7ygU0ypV3KoPnMG8/tjsJOuuHgcc+Xh2U5KUGkgj0pjsyl9ioFfCP4xbIIuqvMtbGfGi8+5+crZg
BMddxPcM3GjJKsDVAwMQT9w4WNgC2tgErzSnRihJUED5jprZ34WZ7+w0/PGIGPAxFhg/upLe6x4O
DMsnRs5vzwH0PRDfUNJWbi7YfwgO4X5A8yjIZYUXO0xkBVb2YglNfbUq+PTW+1BuVvR6ZN9Eq1Kq
1i9eCNcjzmOoAz3ZYRNoD4XM93BxdyhmlH0fbj8N28kKG5tefij9ILdwwFoI7mfqvCcvkjKEKNVE
XCQubWBCDhgr32QW9F6RM2bB4gNzn3wvOLpz4+cYJ102hM37cBue/J+gjNWvSbLgd4/vl3OPllS5
BDTJC1SvhqngLtvAek0bsg4ku80ZgQjAIaAQYu60jjFqvnqJgI6wXdHecMJ5VAO/IGkCMTIWdEEK
tZGEzc3na4+eDZBPufd4nDCz/rayuWRSxj5AqtPE/7ZVhBdUlb6GdDqdEflLs/SDO9+iCpIMQokJ
pNqla23vlesIy95Dcp35C29yKz5YCZKZRqWTUEj3rHMTo0tJT+8CJmE0Nftlbd6kLAyEJsVmZVHP
Zz6/Nquw1IV4zZy5jWHvAH8wO8vsMmPSx+V8lk5cAoSbNDbGRPIKONtE0eAtZ1pmpQBaouwOcT1s
PWN31hgkxjbY7aROs+bla4f58uxabmGPq8Qe71qMkEd8JqEfnPH1uUond4kxm5cIvjPsUU4b2tRV
qTOK6BC43hpZxJQpoerPjBeEuZz8x8hTFxcF5f2tsU2xqixaAc8WW2Yu6tWS7tiNC6lMEl6RQ9w7
UJGOrdWMoa2XHtuRVd7721VMaA2yY32QHj/720xdsSugh41H3TY6dPLa8dVcjXBGkZUnvKHa4TEo
cqwS3FAQ8XTx3ow3MQxa8W5ERzlQRPBOqe+Z1ziFFQEnDWp5ESloBFESEpBofgbq3iHtyk2cHBXj
T64Ojsh1uxleYA47W8BtmhgzsGBz6grbvcCcum8uXUoLkWX5mgEcVzd/a0h9+fFPhZbyhy4aIF5F
qUb1UEVTssuRUqapCeuXHv9RpzKGuxvKnoykAo9AdVWlgjhPCdzpoBdumCiFy2CMfZdked4uU4pC
oQQRLx3n8sMD7wiKfrYRluuz5Uq30uAH4HydXJ0dGlKk4pKY2DPUbw19jNQuGRYV0HgaD6m3WnJE
/Uxegec5TLqQstWBnPrs+ax8ZeOeudUcGIIFbjfkoZGgIn6lY7BjOU+48mkRdkYg320eY/tBM9zX
gHt+mCeGSLaHVhFW8uXeOJ3sAICtyRH0Q+Z3oKmlgIz/C9iaEaTp3KVGMm1udtP00f5hmHGVIn2+
v291TTsEAAlE8mgMpdSUA1emoUOYuHYEkTyHhCSwGjei0v3wPvGXLazc40CHXiQS5DtUvOfdDqhG
APS6ZUBgvyKTYippINbzMr+it2GKdPyEluRt7NuBPxMtlQNq0aJ0gqocUG8ZJC4joKhQq6XZiNCt
oet0wfXailCTgqmIYA3UD893hDiTscwMc+GnkoAR4gqu9+1aIduGAYRY9sRZMN3g4vOsssuYhYI7
S1/Eispi85kw6QB7yOavKePLLswmDbpRkn2yVrvQ8/q1He82W64B0n/aYNulAXVfp0maIHGfX9ef
gWEnjNP4pStxHi3rEg8l4VyDA2LpaYoAYuMPY0U/Vl/t0OndTHMu/olQoO32cO3v8Qd2bZYEQBY7
89EvHdwDXo0TvXc+1DN2GHVRnEQmEAneQMdJYLVBszMVAFaxapjnHTCu+eC56i+2z67rAQNo2QA9
fev842ynFLI1gtKqzfpZj1bPP07NBnsAdjONtnS35D1a+GawN5qP2geY1ps+oe6LZUu199HwNHGZ
JeWdRebLylmH6uiRzU3b6GMzDfRTuCGP0ShmPGfKRdK6WgDFHE3RXlVg+XtmOZq0XF93r8AgdZHh
LMBXWU33pRV4hqmUj6twr5AiDd5SfxmRxT3xeFFjVGg4vQpvXbspKy5dEGJGRnjlb/NtIyLZXxT+
E4CXT2Fp+pPgtTLtMXWK7GWlc69gjQYbEbo+FtaDW2UlZJ4+LR9PgVxTI2HnRt4ly4gZUDXJ4bkj
1satLjXSeS+EY8w92buQufbuzWIovXCKI7omRUaYDMuaGU8YV3soh4puAczilqQEtIhYF0XgSw6X
B/AP9dnuOdQL8Xj1iJX9pOI769s/au9rzsobzaUiYI6377Dj9CWpxoBC+T5jKC7T6bCf0xiPKtpK
OOMe3n5hnRkkJo8DMMu8MsWEo9CcVC78dfoFsdxZpEcdOlOFD9GwxbeLV+T0HTTRNl/xgecY9MmY
58zzd7d9X0TMyf1HqDe+Ds1+aQUL2WBEF7yV+nXUHmzY4gpp0Tyq+CYYCfxEidlsrI7162VRd0xL
rpwn/75tAyaGXJnvfEQJcp998jsGtlfirKfTpWxB4ujfkIURBgyUO3ZTqIoNwzyMOeOnBTOyC+W1
gSxIWMcBQnQvq3Q6zBTwcQ5Rrs15GudLNABvDRxMlVtABu9fSnF/NajvgdZiH6H9K9jj9eXOWGFV
vCMU2YXXpnQg8qL1wOpeFdZ66nOxAEKq0g6re0Y2pXyaY5Y3He8OvD2AWK+Zseq3CfIJVsSmoW+O
nr7hczkmmJxXUzHukzzrMnU1KkJlU1Xp9ZcflEpdlOHS9jiYE3qnSpRplh6I0nhBJfK9pvc82evJ
Ndh9p76mPzQbCDcvkQX9n/wTpoA2RPCDHqMXm4xUaMVn1uDQQRXCl4lIKpw37SYo+XNZ2WHQpJVy
iUqzRss+3mlggDARLZc14YuLZQvNviGoha6iVl+qNBGrzrtXUZPIYGBIHXCk1K94wAtltd0uy/Kg
4qRZNiFPHgD4Fh1iazqjwTSr7P6OjUj8HznNUWMc5sFumgx2p1rtbN/RdqUZMWP/jrzcK2UZih7w
+2MufLAepSbgADPmb/j/4TOm3hOry27sCIkwajJaCxLDOLVK1P8t9FtOUA99YO//1WAwqhPmDD6Y
Njq/E4kq1tLnQmeKZAjNg//1DTbxOH6FyZTiatC2nUb0HNi/Bymg71e0q4j2PtpLoubTSkA1MEhi
BY6Bm7bc/OjQpSY+b32AYEfRfpS0pDii9Jegp4HabcY+kopDF15yfKTtLbDy/p2gNBEDQmoAVMwu
J5023qa3OiB7Yi/JqAcPU7SX/O3souZV8+mgohb1evcfpIxRXCVPtBUiIM562mVWHdFncw2+wEB5
wK/MWjwjdS+Uzvg+vD1ORUmeI/wArG7yUmCoOob4WbesKesP4JxjqUmdL5TmgbEqRPNW61KA+DK6
rroU8N43aDEWJQ/Z5jTcMX59v2le1wIF35vLZfhfO2kLx0+LGB/lU1OP36pjehfu89QAJi6w5fYC
PWrQq4KOL/06pkOXZ0F3fsitifousBKUaro6nEGFqLcpF8fQSrLxsli48VYUont4mzysdPNXw0Hj
whdJqd+mHLPiFOPrUfPl8i4k6e53Z3woXtVnC14/8JOLIQw+tC3HI47pApS6u4ARZRM3Rli1Az7K
f66nTqRZnGqipRkTz2VOXxBPvL8AhRGpIb8jvnByevFhMxzIc4xIDbXUa4aVMuDJSlZnfujrDOik
3wHwoNwap63DVOrBkWj8qKKq9XOV2BKwEyT+5hKyYk/X4OM/hQ+EPptO5eAQfBn8N+3EdDnFPP2W
OUjetUWFCj2GVLdXbKqC2PWdu1UN839KbqqwbDeCslqW8qyrjTsrM/uKoOhL/NI0nXwwcJgZt0yn
qoeSIwa1L/rJWtmYrJ9cNeQFDaZ76/4PZfIYqXUtX1UV0Vtl5fsje3Iub55gZ101eXEO3eZC4Cn6
Io+5ECdS9p5EQ2YKSBrjM4JCExpjntPQn4gJri4yqcTU44Rui9Wv3Og+UgmxepHNQ3wd0XzhFmtX
2ll7Bq13a8Yo95kyKSeZ2+77Iz6FaeLqYKWBCja4wfpkgIra1HoghftkaBhjRej9Y1AiUZseHu1w
hS/QpKz3nF/O15iY+sygeoZih2Bn+KC8MrRDZuMjbBlNzzjU3abAJQ91U35E1cnEgrzYN45z8J+R
GrUkxV+leukrYFIv7JgX9A4Q8dfcPlcANx9lZhCF3Fh1tNljs6rXd3cKTOAufmkNGleXpIZ/NVKj
neH16vtm/4vNzNEiyvNw3/wFNZ7JnkSI/OX0jeZg68qd15ZVRghOAr0OaZRd++UdUno+6sOz//sB
rUJ+EUBKe281FHu9g5ysHdpzhNl2NYkGvAsvoQUvJMww61kWnj/DHRONeOPHTRz2p3GdTNr9Zx4T
WiaesEZ+2V4edSjYCf+o7u+vcLbtNwgFLwO1VEeZf59dFhIH7ORWud2hj9yGjAEAaAR27AqoG1+0
OZd/+5O6XPv42BbnoKOHYfMiYK/sNl/WhHJzSVH+COIfXVp6Yi7nGIUe5/JjIS18t6hyeue5XldI
geYhycAwZE6wreqlf6O+mGpZBeSA2aDCbN/h8OUB5X2tOrdwuOg57/CHZrI5Sl2b3tKVyLLdoKg5
lcDX7XP2xgahzTJYSd2T/XVZYknlXxjv6BgLPnRZqrbVmuqbkmqLfw/K07HuVnl6NdbSE1VqjG73
D5Aw/wqkEKVamQsA53RUdYACJTKZf6R2LB5TAkWc1hQ95XbLU7jUYgf83E4juUBaqwIxS401sXUI
VLhNtmk7Y+LP7ap3nPCZ7tTj9JNt2xnPby6+If/K97g6XP8x2V/dScz/aODeItLaUWW+A0KviTwS
duzGc0wVooi6Qb5JF+8BWdepWIcZTZm0W83Kx769n5RSGtjdW25Sphw2btp8FeGTmqCZRb6xzehz
dz9YlX4J7zx23AbnNO4mB5GTp3EVU1KPVfGkaS4WhqOcWB1C/kjpt/BlUZnIVHHj56BWLGpO1qF1
jKWX67r0Hn7d35pUI486TAEpMUZ+OGN1fnam9qGx49BKWijqIZIbiDeBPqLGug94Fb3nOtqUWYnO
nXh12rBrQMma0DlXOvceVpsXXTjeR4XJZNVR3q+4DXFDdtgULnA2eiEfWP8xmv7mnXwEvbik7kN+
rulnyQfIpCdyVgywZj3Ub6nyXuWGwmB0+vl5Sz7pcZ9uzN387S8B6tqui54tsq7dXRplST9QfSRH
R/9Qnqhm/yd5856Pbpdc6H+gCAg15hZixgFOKNijMGPoqUKxUb4YtoH+0NMnStPUN+hZ4vTOMA9u
7qFXg8k3x6iJWTB1VSwbkn3J+Y3d6w93EX3RRuUQHUR3ruwaIkjpEGZrZihwnarAzdOBpu5nwO6V
Dd6JOHtD20pdeaBcJX4B7sWlkgUL3hbpz/mGj8ErXU4UyAh7nAWDZfY97sYRYJIpqHrJnqFcB+h8
IF3tpPO5J4abjIi2psvhIAtEK2UPTH1xM899vKYAZig91BN5i8kessXSn2RJy4VHsOipZNLC2Lo5
bvI3HKNmUvJ1Z7s54xVML+01+kRHf9vJLa9IAwTWckMsd78rm18h+S6IAWLBpd4cd/T4EnPpMCFH
26Do+y7Rq/i0IFisdFt7P0bNluIljeTyFhooD7SGs/wPtwYP/CW3fDGyoAXjbMwDH3CfHojpuAgR
bZoi23lEntCkAd3CuEBHP+iE5zAaIjwmXgQy++bl6MbUZt5HTHhZ/q/mG7PItYnv4Mw3zo3CVQcx
MbHXEOEmH1doGSNh6+a/hGQuquHeWOEp3WA6WP9W/fSU4H4JtDfm42SiazKKfCfhqSQ/vqwCq55D
AmPk8KNU01jua7gFfKqnoGF2JcSM/EMQeTw/x9WlB6nA74pFFeRUzdOK4TW3LMz24acFSKYbI9Zd
L0mbpmnfHhmBfmB/lzwmrxwqheTYPKfk4JTY3aBDN65mTCZrwHhajWR3sY4z+9oGlnIC8BYDZVom
vzudAohafQbbiJ9YRatQ7ygG23IpARhv4MK2r2UtXiW9decabcm0q6XIrRdHwIgvzW9esnXYhHif
P2rX7/kDrVr+Tev4+qe3ivtDNHTpFx4LUauEZyU+BKMGXHJnx8vQF9PwYj3tD3iQN3jt8l/1Xnho
8Qsq5+LKtqHiktE0iZQBbwn/0ReNlXfyUvOUexj9zwWDhwxBdgZitXXeot9Bo1yTPbtEUJRDSzCd
PEePOcRrDNv5aqXxgndq/+i4PBedXyC35/dicrlowC1Kqzoy54VccKAnJh6ensiPBJp8hirwWUKr
jQST4VvXLkeIqd4clzu2VuB1Am2S6Bx4KXQxF/HSdrnLf9kPKYzxqnRXHxfIJSJTOp2+MoXZXF6T
H3NE/AvLoECoVf6G3hudWX1ZL4/kwVsFJUBt4bQusl1aUPcF7UKpuo3+pBeQoTjFvR1VXMh4uxxq
Cfu5Zsko9FwFmowq9PKtbOCI6lBJTRvYxa1ILXrJ6aM966Zl8F+8dQ5LdoyscJFI2TMP9cC2PJHX
DBJNL/efuIBlVrIzc7MBYr3ikABkvkiJFiVnHT/HwQzsbCjE4kzBTSBNm6H/tGb+dXvKzGSoOytt
2knK290gMw96ZTh1KEsn6s7eZMdVPPXdFBqJMJBkR7AO4amAK5Jm4rV8lDfKiI1Jy9tkskLrGpOW
NY9qvMWPnI6jg4hIy4R/aUIrCBeHli0aQpxhaIFSwBojlDegu7FIttAsgF3UJ6YaAgVrW5TD0C6q
MclkBFSR3OdWFWd4ZYD9PrQFEERP3gGSkFC5YImfLC1Uaw3Wj0E6b3T84qhrwFGk81Lrk5skUGj8
6vyNCXdpd5a68i0WKrVjhKtXIC67eYa0PiA7Uja4/lUsfuVmO5AFQb6316duu/gI3jNj5zW8WXNf
koSd+Bue/e0Fd2ULFnGBlOwmpWIovKRhHuO4G0nj7qZasNLQDsOofB61aeaMnnS+1i2q3pvFuKt+
sXK/qRSSYYdezeIEyV5HEbkkv/8Je8b9GvYjrCvOfjcaNzrUnd/3HBRGJDOWmCM/Yh1t/9XChDVi
Qi74p7MDQzA0T1VaeO3sdvhdeEwzAuLfgYyv1sjxO1xnmjdAo4qAuo33IwI5XxDRWxzzb4wMYcm7
+IzMBAs1T+KgHb697FogUpftpkEKCiDuwkt2Pzpd1CGg83Y43rdB3rGYeNgbTeZosD3AtY1GD4O3
UR4eFR1SSugjPw3/mr4V6FCIJWb41NbN6DMGUCR0KG8Nq/qJoUh/I+Z1QOw6w6SE9BNJ6hyXz+ys
pa+E5r4erPWOxPWWVwskSCfpk0DCysisKzw0978dDz/3w7PoZiWt9F9RpSud+4IYpYUwmOGXjzDL
Z1z+uqes+cn14fUEyRaw9stzDJ5HBHBkMPmFs/kA+WFX7+74ywaKF4shOcr9p561ca8LpiU4++d1
IMzwZ1AqU6nKljCrK4dSSMUxAuREkTpeH/nJsjkZtEFg3xhgfqBaif30njdp5CZhIxEABtTMz+Og
pAPyXgMitePOKIDvcJlW8TFAcxwzSz7sCv1a1LaQUtGfWWI+6027GRepb+FmMV7L7JDxpeNjZIiB
iJc214pVtkaBHdRzV/kqDpBkKzXTrnon80g+gC76k3POfSGBPFT96Qzp9WqccrdU5dV+PGgIOVmJ
lkFqciXh3lR3KXyEDUkTwv7Wd9lrivFUTpyflt/jRKr/AGtbx26YitCYaI+50KCNaLcrQt7QQLst
McGqgsm0qRmCpf4Ikh5i8gtiBb77ShlISZX6+kofRlcT3S98U3MXZK0rm4h9MbyJpC1TPGQokwt/
PHT8It+ExZ3bTshyMUSnHAYoJp8iY8o8O0VPvR/C9a8swlzIJPHwsmV/UySbooYBAxjTTc3XIKxh
qhd2DLjqgQqU/kWb6qeBRAFdJJ+eBt6TXCVsqU7vTriynC5dpKnynce3ymblRp1OyY506JpFAfA8
Zxnh4jbu0+0Dsn4Fwj7mQxEjjZf1FMTb3KpCg27uLlipqQ+BgdUoTI4xd5jR3f0wTtJ8YOTRM/5y
bCMTs9HrX6pV3a/FqMbAYciJAXRerRPKC6ygCiK4vKhMxYq3Jb56dBFL4D+VPp0fqyvXBwEmVaOQ
RyVu/qtuqDtKhiL1HChHe+WLZCxM2mrnapJhq6Pb7bDIyls80CsnoMksB3Du0AuEbYnQt8STtcZV
ZJS3BwPnNFbB/RYL6KjfZdjKMJpKVacL+FrbQM8WiP/RInGsofCHhLvdiuNOqFY7DaNMmA2iLVTt
+o8f1tuPK2Ery3yntWr52BwU6+pl5ZbI2YhiSXQgpNkmHiHdH/siQq2xReTWf2vzujmV1TTKU1Us
Z/GZ29sBqYuRLC2AiMPr5nv9lRloYUvP9+1LK5V5Jvifei8XdsPpGzFdBqemR674JlBhjg0WAxub
erCeIyIDLd4TBSBcT4GPc+Jz5x0ZkjuIhqTlOUTmbnwLG4eC8ldW/mf9jVSaqAylcBAR2TCo1Inl
JkwAKoC/qu/TXArm+lWKccAXGJv+TTliFMGNDLM5irO9MZFYNSYu7AektbCYxomvkuBajfhPQVz2
rpWHevWq+O0gZEy4AjqWIdQXVHtIqIsqAyACAMlH6/UBlxH2HHyQvNNUeOm7z0RgaBchBn3/F0hE
uYKXkTeHNSahVvCZjy+bKmL7nTCbpURwFYmyUfztcD7m7OJXuFI5Yz9vhfv1ruk7HTUKo2PEQqiX
TYEcaqxcH0uVlbYj0hUBQvO0dLEoamZi2I3jad57oLd/DEb1ax/iHFYAUbGShsrAPaDyAFagnI5A
DDmQ+2drDlhCzMrL1Ahhf9zYhru7Hp4Z6PgHlhIP62f+7XXswRu3pBVxeJX5yCEc6hRM2+y+QmO2
JQMVtmyn8JRlNCIKVWhhmalVA4rFP7y3YAe1+qbP677+GQvLZe1RzFbDsZnaWWKoKLN+B13MLWS+
4D778C2YSfKbOitF1fGep/Vnjxz9DC7htzJyRzN0dsqwEDRLPsuv2/7BdaA9t3SSRwPQbKzrSuGO
OD/oP3Z7b109LXDUV9OepGfYczZKjRvZiNHqsUtukYeee1oJTEhgQHGfmThUYpFRwp9nE5j5YDTR
t48NXL/Hw/qO+fNxa04/t8/tDyJNdi31qP5aoluqDD5y8sO06h7vpeFmd3nv+BHaFRAbrGN2VLub
rx/wwedLdqLbxFm5uqdGwxNgsIy5aDgvJKbEsbZ1VUPAEyBRs3E23Pyf6uCy8p0INEkgjI6eMuFk
FpHlUrFCCPmsU6x7wtRpN+L5mkjxbUiezqyKx89B9M5MKgXNOjIwaxwqrHZkIvTlLMEoytlCgkhx
jfCN0JvZBz2118hvkOA8Q3sdbzTtoRre9+ZCuSRoC5IIjDkRk93/y/0mELKkzWFZU6vueDsaj2Ct
g+Rqcrfk4Rc38jZD2c74dr6yQ7baqEuSEV1xvxImjqJhO0jVdcgTbBl7so8itZF7l1HlF/fzqg1o
Fl2cGhFLxJqnW+j3pCn1n9mdDM85B/lKhAJGOHRyijDBT5VQ3xApvFOiXLa8CJJSGLo2pjIWywVt
Okcg8Sh+jqRmg6Jw/tkz3DIp7diB6PFeKIcGGgpyHNW4UNdDJeNxX9OC5RyTh7cALISzZi9eAEtq
0k2K+v2FUNCQAXBMvA0Pvp/b2UvdTZDCsweFIdcSUDxbcmWHDms7xFcFAgLHylWwFl5qU0zku5Gp
3/xglzYTByAcFZaZjOWhOeAIjEZbA3VaRduXsGWBVXR33Ia9jLkDMRGzKBHL82EPAsocH3MwtdYw
JHSWNwY+K0WE90q2Vmsf8y4ue505qCEqyiBUkpY2PQUj+g5nRSgJUkMMOgtloSjtS6oaWUdNY8DJ
2KLRlVNfGtDQ8zRTXJbfCZQ5JJt6ENSbuZYPeWwqhI9g4p65FIfPt9KaKW5rujEOU/3GAg1g5/W6
ijJbCw/nliJvkhr4F2aTF905jXfPeE+SfxTkYzcax4wB++Td1EZbGAHUXCy9U+N2n9WWzrgqYqYA
CgwaZ40jZqXb2gkaaWPm9vWVrGX829R6Zg5n2lsaWxoRlJjGdv8SXfqbtNaL5ChiKhR3iZA8FG3+
bEl+IlToIRR/sMuJk8QQkm02xskfSat92xo7NWieRCO3xnQB2UgcLJUQO/oUOkHVWo7yTq9TVV1e
5cudoHBmciIC6G124GfB0G4hAZc9ZnoVxWWBs6mwM+TwG+XumQgAlHsX9TU//WQuLD78+YUxU6GG
1TyECmXJzonqMgE8uYDB8Nnt4aedkXeiwCsBG6fNgzsQmTAAzKROUlisYblDYlE1+lqQRb9McDyU
j6XDWaH8oaVhWrjlFhfXkB/MEPEAJm/GzqtwO2TEaQjYxAFU1ymVCtqAElZxJMfCvKTQdwT7xqgr
AFd42D8CnTHAweCzYIQzOMmylWDSotmxrwDdhtK3DwirjYWNyJnLC02Wo6sI73smmmFADktJoKBq
TwnQ7/Ue77DTgzy03GpebKkeUbp86bs1EODiqL2rSu7YTgJCSvg3NnTPcFR27TYfLZrddDMzeMHZ
Zlbxw1Jz/IoNHmhX8C2dfF5rJ71aqOkYsgYXfcE+eagJ+chpWpOmmh2/6SrmMuGVwgdMp4Ey5J4f
nFLpJi/nHOOBHiflrDZXaGAEkODFoVO8EJJJbDbktScBKhtge0hITE9Vc9gL5mgEokTP8kWynDTc
vB+yemTHjvbOaHuT1IlCchZXGPESLKgngfgh0gHjvG58tY5MvMLFGueDb73a7Pnq+xx64rPcaWTf
b8bfqa/3zUVxk8dQKV+SVXDPQT06RCTtgZlbSC2FT/jTIUlHPxObrNOZy8m6Ct5ioJg6m7RglEHA
Dj12Ez1ZW6N1TkYQ3R00waMw3a+ZS6Zdz0/Se9LzbGEu7MzJ5PiBs6YzSsc4cl8/8cRkvUy5+vqW
cMswu8T8BQ7+bFoGWTDR66iJw76ErXq+Y6qVoJ8tT/3AQiKC2IzE9q2I1y+BvzX8bBPmrSOXGpjW
ucfjkVvDjxmLECJMesJd0g88RrkPZidOa5B1I9ayrexi0ZLHLWrgQARaXaQJt8xHguVe060T7Op9
LPX032WXiTYkh7gZBqZ+7nWUkULCYm1cI7pCbOhxZ7htQrMTbLC5PGfBgavxkJCyxAMZ45Fj1f78
fjqTyj9hzRkIl2JHzU+TSpWx/Yhw6ZlOgtMsOfVbrLucv1k998PKSxM63cS4o3FGOaL3TmgOkB1k
kl1IWXOAnHkH6Pc481Phoi3vuTmIg1Byo2soE6jZuTMWVdbZ/4LSbJRpQc2LiH6CAefc3xAeyl48
3JTIB0+JOak91mGwaPoj7ckTJvhwBGA6RNK9BdT/w4/sfsFoUotGZxlVlzY2UPBhH1Fc0EMjNvT5
Me/Z8TToIcCkD1zjSU1o++fPRajNtjchu6V50b1uN2RPHlxbGsYGEjW0GZIRG2GpNhiyXYIy7y5B
2XwnqCEoYdo5QDYw09sSCUlcGzuGG90I3iPjxoJl4YyOOKeb99A9MG+4TSsOTzI10LbHIx2vMDv8
A6nLW5c+SB3JOS9o0QsKEP4C9ik45Pfr8X2YpbGZDrsBctJXg0VlJgj4UnyntQ/gX+9Nuff/yN2r
AP51Vu11bu+dn1F7slmf56bV/KS442e0MRbChBm8hI8ISDlQ0E0P6S6A/SGA5nzafM0UYzDZtrsr
wYZ/SUi2igV36YMJehfVl3LEW8fAxqBIewIkziAVkZg75/CjIQEEXd6cn8TPrEybme1AcOT0YVgF
XB2DiRR8tvGX6CtT9ORbB6/7o0llwS9baxyHbeHqRuzusMSNTEGX5sxXfuq/zLCVf4pEoLoCFdJV
LsWQ1wk8YS65CxPKIOOTsW+tkwrJODPP1OLbc/Ark1g5PIo6ozx6V8cCXqwxEeEn9r6fFLfjga3B
bSarFUU27nVe5W9/sumg9kHGVJuRF4jx6YxulTao3PViTfs5QdBQU/Mydh/kUfj28DXbZYcUa18D
VQUBW7t1NrMOdCx2PqcnOflXHThgSlb9pHWQ+mwWV3760/gDxDJusCfl/mSHR7qascBe8/sgT73m
QDeEtjUE48AYjR9zCjry0DoN1tjy8XTabEeQB6Pn0FmYiQFkXuNC1XpSGk9YTDldC9P0xX0IimTb
4cj1CXw+QEx9VsBDDR77H/gs3qGfZZlzJpMRUbohMPjqkL6DrF7M1dLrEk9D2DWA+X65Dj19MiIB
zV8/4NMF8ARo0EdgwchJoHGUVD2Ha2ssBbce0EaPA2slPjELuphmZv+i+Cqh5VDKUPBMtdZWfD0t
BLfzYNGoUUnvaJRZz5AV8H9GBdRE952gzX5iqk9Dmj0h6WPy5/XY6QGFSPbJ4Lr4r1kXyW+dTMXL
cUdDpEZcxgT0zjG4dwhQlWBEbtiz//ioYevNwW66RxSmuZ5zkFmE9DRN7uXGBEStoZ/bWZt4EwDL
W1VpuGSCNN9SZQgRD6MpmGSgthqF4Rv2btQihTT4x4a0jIReIPq5rcnuuVw4O0fsS4eXww7DBhUM
2emBpglvXGGdfq+/Kqep0lmEYBCP+G1fKJ/aCKT6hxLlmJifV67xqiX7xLHUsWckbI1jM4ta88L8
07xIO/5dyq/ZRNyDe8zkmNc4AiDphMK70JH5IxG5A58O3bONHfdgTga1VNQykHSF1XRBB4phNF9W
aU8j4SXXQytoB2BUr6iyep9Hkt8UY9RlHTKBeBmnt+KNR+YvXeLnANSTsP86EMgWLNPjKEc9Suw2
ylt5I0PG6H58H6jDNvsvhxpSD9rPyCRk/C83kVu+EpdT4jglKoMN6S6+JbY3WojwUykF9MtF4a9v
MZ17JovvDHoqlopTDBvbz1LpTCbVYUsW8SCNaTuZhpYnpCQdqlKU8Po6mPuJVZOIxMjeZNVIhhZU
0f2LREJwQhTHMSD1/RAxxD+65MG/0kTGeuD0xu0A1ARgZWzUR+t9+kTwiZ63ve6XEAo9pjgmuNNK
xdrPGkBPxdBDmhY/pMp9GEPDBBJYKtI+6r1FrDKyr7uJQAm2yEDnVhnqi+OzoplDfs+hxq0Gebk+
jj/E5rNjunrzV+uVCZPVzALQga/UVeNrNSVOJ1H+8BFkmyvdY9XJGAPeRf99kgQVkZ8dtmTSwZwV
lx9ExnX463ipMXSi9H+pUn11ctrn+8XZUNh0y8xTaeM8Z0knvszovTP2zRF+NBLvf/CCHmP6p+X+
jl2oxtyPum9NO657BXW+BX6BIDkvhgY2tZPShMAwEzry3xFBQh3PgSUvkgrIbxSDfU9n17xPfd2Y
dGwdQCjWkZjgIdangRrpwypqsGEY5mvs1AHttkqog2fJxj6O0wPodIDIv+JioF2JCMUAx1SsO/Ok
+r6U+5rSenhflk5ths6FHcunx7YBem4b3D2No65miOLY/AgK2l/IF9qh4MlxfT6gWrGk6CzOf2+S
gKGYlrUqRRKUSzIUDymFdjyyTg8wQVl2amDQ81GsMLKHApmE7Z8JZrYNXlNyQfjgDrZQI+14QGTD
o5Pbc6jN2cobjhj+8wvnaWhbRGONj+rYLQoJuasojp0HtXECGj/yHPVD4Ma36LjwpwquVfTbuShX
sKllPIKTRTcYlNLMCu1pNPMM3Vm4Hj4vcElHUL5t3R8wS3YcuRRJClVdEDEcJFcdCZLwjDp7Ti4e
kNiumHtej0RLiAU7Xx3FAMxeeEppb5IxDsW+EWx4SE/hsxqerjxlAJyHc5idLIGZbYOODjGzxnh2
C7UCiUR9PYfRA9CsLB8ts5pQK1+VtJiDD44rsQYi99CNMagVQxl3Jk77NaEd5JgbCkpn6m+KRL/1
bcXql1SC1E8sR1jQERYz60P1A9x/pWXhHbk9BP2Kfsovc3muq4vOQ19GeKliwRzbpdva70gqsaKU
ErIni+Ljx4nYHtlMPiyU9+WABLuGcJOiyP8OYhWGDx8Z1TEXbh/RUUgjYpJrGqbvc4AdCCAv+FX3
nsfUL81EwwwIN3qEI3i+IQK5kRn1TYuPIA/0LPIRmDSdoeO0J1X+HX0lzf+4UsusVKSQ6LIVRzG0
eI4mLUvIld+q1KPoXCskimQnCRxsACs4iMMN5ufhLSAvzlNKS4EAmSJZE376cnXjZ5CpjnpBkF+P
7Sfku8CHpEmVTBBMBIWTYm1I7Mbqg558ZXz6or+dVBnd29lUP/YB+IMCFrG/yn6qJxsbJMibnNbu
/L9zIwZhqiTcZDn+w+B2UnPCCrZPaE+JCBAe00pZqRdNRN2f7NFRsCsHxwM4Djey1Cj6LCtUisvw
kb30G56VM16zS6c2vxffIcqL9zr8qrvE917Y88aXJB5mwi3qazaYRzBA7UP450W42DkXxEGjO6e7
DCTlQtt0wEeznlR4r4jRXi5WrQsTIHgD+nQdqCB7iUk3EqVN6jMCUU60ytgX761ihjrXqqHAETdK
++mxNuRkChKSok/f8Lht7im0Jd2LHpPIq6M5j6hXOnzBkjb60GyOzWdYftE4JVKF99oTRdGoTXvC
ljRRBq5TAo050WcVEL1XU+MuEgfPUWiYbGpLVULFPAoeZSA1TDMuKocksepL9Yo+9FMMaUa3LpCG
D+s8pwNmCE7Hj2XKs5jm00KLwo3z+QQR+e7VUqcbV1/ahHVU+9E1RNmdOcrn69E6QF6yIyaXqdKQ
XqDs7RfDgiwdVBKyUzBslt8GjUzRip/kyJKxUz4Ecjiq4qxGRMR8MUX2GexIg1ISapk8d0dDoVF0
HoRszYUH/Qxlmb2r9VeR/A5NKL6RPoWYFWgfBLHbZasrnBxDI/HadVO/90hSXNjeKT638dijyK2G
9iyHiRJEAxbG3pt1WppI+Xat//zh1uI8diz6I9rwQ0TVUfxAoRHnyomL4ZHKnn15w5oT3x+Xe+y8
8TfHRPDobcPBL1S0CbbwYDX0779yV1vbbMMsA/CMu9S2WOo/PLv3pFRXaGTqkRHawxtOYMkg+iUP
xxYCu46lnoiAz8lAtL55dvX4JTSMDZzvryO3SsYymwZq7ddptnkM0ZWLbaFHyA6ROiT75l5AyS7+
f9JSh3VD3DMKPaOm/nhmNMSiSHAo+MLF8QHiAhHx4Z3sKvUs7saKCjKb4Ba4t0wewesAkAfTCbnf
Y3D0PaIeqinSQxRZAKk1eubj9+MlszJE52WuDxHWPuAC6NmywPD0LQS6Cml/128HZ864at46o/t+
nQxu9uOKbtnmAEHMCEY5cb1xL+dwQLm88WvOXPSj2eiTF8w52CTDmDQIVWycci+DfjyjESesh4KE
kfrSsM9s4BT3dcBFwEPeLSuXug+p+ESmKz0a/ekWVgsOqJ71o2ccK/hVy52fLhKYmbOenxJbrEa4
jWhNwpBRtTNrfv0ueLUGSkickim3cfAtYJkNhpt67C1Dd6PzDcHHMxX7LiUCzTu5P6Paytul6Yu1
XHVsTCCQymb4HHFAf3D0jnpvzPkK6RRl0fheywK8ktxXlvVIGl92sX+iqC8D6Djf8g4BfrHFFsX1
lvnDXtLqct7D+ZGqIXEdVcV2zONqv6J5jZ22Ya5j3YIp8glPmb1tlNV5mBs+RxDZYN3g31Z5gEIA
VpdjjzKn7moQvA6nREFgqs32NSa+UXwFbsZVJefCmJvxelqSpi+bvqm33tr0HAi5X23oxh8dKUIL
LxIA4QVNO2jLyqTD1awaEkjXaURW6J15MH/IuCj150/+lj3fG0nCyyF7c2Pf/3M9cfsGu7tiuh6S
cefbiYCDOjMn91ESyg2oemp982q5T2nUePRzkAXB0KX8uZafpN7CM7hEzMUwmoz944Ux9/Bo5+ja
/q/BlcUM5pfYHhdqFjJMF6xKsH1NwKyAiKhkeVn/fhrfuP7hRLwnn03pc5Oo0zsSAexFm8otEtnN
M4eCq0NPpcGnZR8Z8tz/xaEsXSVUQW49j7MCZsygciHY8s+pG/MixPZJtzMxWYVWgcSFSg+YvSgJ
OP1NRSx9uDq+fn4mgmef/LlH4dW+CebJebM9LUyBg3b/34+bh6cuHsThNHAQyPkRJFvce+qu6TuI
dTzpHtIx3WgnDxnYv+RTJSw+lWDd3pf67zfIr/f5G/qkvTVxMdWc9bdDVY8vxG5V8+D0iP1EGEHY
6S6eFUeWc5hXvBxHB+x0jKV+z5wz0qa2BesGVB1kE4RKznsV+e8pUa5MufPoScIRc0mm14kplFVQ
ViSt8XJhLT/J9DaVDirXkYR5xukxbNfBSucscJzfPpG0E+bIEZJauJUGchn8PFKFgr0ckDrfZ2QF
w1NAJXhsJD0H25g484vZD5pxrUoEjVs2igl96kzI8qfewWPTrrvKFPv7LQuCRXIKkRCIqyrHvORz
3MhLCIr2ck/BiQcAx3rmojHFNwtkIWbyHq2snd74399cLbMlnr5tICUcG9IsXZ3V8xY9H2OJiow5
ah6Ek0AaozmXaHNbkQHMusrfmcKUiwMhAdBYDLNSrStQZ1oCcNcWg27SN3UYoUS7m4D2/DKL0cUP
NuU8e68SfCmf4tojGn0fNtFwsJ+A4jTRroApYekP3BGE2KB8Vp77jRyGt6TQJ5I15+K/YHNml5CS
+RN4w035sE16j+gSikxy45+EBnNUPJBeNgLsqaYiYlUtKLVY1jUkv5PU8Gx4JfLUIogI4daA3xWZ
YYGk3q8PMe/5UXgWceorKDSplieIpVXB/VdTKMvkmqs3OSJLX1TI/1z0nEw8CFgBSj5QVKAbR1DM
QsTcY3tlY/MXHXY1of58Eh7NoXmXzP2fg7F6hfTSETxuOcO1sOo9JtVqGLIhNOEs2IRd8uODsRaS
rsA5owlMgqVzeBGChcC0Bbxb3rV3dgl6P/iOBHXzGQABtl0eAqH9RNV6S3JwJdXxxxU0DyyqS4cb
2CTT3Ycrkem1hHgbI2uBfvg03H8GjKkBzeDdu8Po/ibTzE1oNlFVukqRGbTn6cvKaUg8EHpxzt0S
hM13RXflUzKngNOe74XxhwlowBCoKdC7HoaESBNSYGFPhc7U5Adc77MyjOXBF0xSMV055Adk8twk
UhXSgZGJ4CNbwUjhZv98+bIV2wMEms6m+va8EgFEkZrcc7mZjFFGPvlIcy5rO5/gBjHcdnLQLuGh
mQDTRnNI065qLcp/7QkTSdYNLbZH62fcwzdvFakRP3HTtZkfH/XP2zOa54Usnkrsxndpi7ge3noK
PxZOEsMbg2f25ivAWOCVDMkyK7NEpQgiOGgZkcnX+mbJz4x5EowZjTkzO2q9YrBlxGwpfwoDC7Ui
NewAZvEUePR0oslMKHMh7ZbfVaLps3gbS319sr1DkMhCwj6ZqSUV902iqaemsWW4JJKe2ALOay3P
brAIET0l3/U7lMVhRRXK9n0YWRUSjyb19LlmRvrCPQqD1C64zyuZK8Iv4JS+0mqiZN/EeTLszHzQ
kzozjBJgmTrw0cnbPUZfH+Jj60Q5CEf5mD+oGvmHIiAs9W12Zp4zLrJm0jkkb0soPycUuU+Y0/2v
UCgRu9nFd/ayatQhBXoQx6sFv79EFVWoNH1WzgjSx5I1/AmpzBPkwmy3wHMUaN00XMfpD1CPJ9Oa
xk82mTvh1yAJtzWZNtf5OTzj6+IGZZUqfrEjldW7zodHQSOAAo7H/CErdY3u96LZuo12//INITFF
JvUJngL4G0L0S8DYxBPwuzdktk9kuJTDvI9JnyMKAEUOtuoFUWvF1MxJ1usv3XWlJezc84LsAF0G
aA4VQOni6ePJ+Un3fAtSDfCFCQe/pYUI2jCSrKaNsWpbmRLCdnlf3i8VgsYDvi0GlI0u15ptCAzt
oA21txZEslwcUqxe7V3ZutX5RIwyXlQt0Pv2nd0dO8zZaXDdYo+6N++Z/5tr2Iy6b1uUnpsphBtD
dH1QDmTSOscu4flDqN3ERKpMoseHXCKwe50N5i5n2oD3JH6R1JpN6UE1nyHZJRdtQd8h54f6kzTO
7QBbHGL8MbPuZy4b+H40R1PovzZvudXI2RyToDhCHwIlqgNVKJ3JaycTbuMrryKlINacq8/foG2T
XmeEjwOLujaJYzDttIfQ7GWv8AGfAIWzP+87JFA8Rv5IM9um3tzRlB97ey7HGXcGW2THNO0os4FO
T0GlqvV1FImVKzs0ArrLR3oYLaF0mJyqrkTYY91KMSG2fQ7iFXsE3FP/QPHGUB2G8KO1Ug9/Wu+n
j0UBL/7YWgWVvSsvPmYVshxULtStGNT2j/cE6gRRA4Lzv8XAd89VEkms9zTGc6ZzssLN37uoS5yF
NcGXY2IBPxROZVMK1XPgJNoXo9LmkX1Qv40MOOC146kJ+rg0qkKLKDazvgqnsWeFOVt9aoFLumor
z4fr6CCmO9Lqoqnhm79jfdI7PgKTA26wIljfahHNydrxc7+LWrHBsOLDx7lV76giuU4uc/iybHwg
ySYvev4NYc7Lij8Tqs5cQ0R8Ds8pKIptjsNJuRNe0yuYhgiC4rdsNsIhubp1EGbyYt4AstkEy3Wu
PodP0ECqn/qQjcZ+C/CaQr0zNwDHvHEPOWt38853MUueUj560859qguiA0T5rOG0kGmWClAMM2YX
kO+5n1lLWW7GOyMxyxwkGIi/xSUxcc/UhWMo/NYfSQNpDYpmaoIMkNweyBOhEW53L9VS2YZsrOST
ojB7yuTrrAVsFFoeXzy/JDL/jrTpzQSJw6TByZgnfE6JECVzn7zHpu6FocYT08e36fmlEWES0tap
EW4tIGKYPy0ykqw+JxGJmGNR/E5kx0lE2xE7wZNOSO4f02ZViUPrXxzdEqQNEgY1k+iwXyw5EeVk
MkdeGoMDxuqKBhxh8pRdv1HJalnb7d1cxAsg3tfSXXJq0DBAjYywJhb3eFoFGBhoVXyzs4SgABkF
ofWa5++grohtsIPvMrkZKIJ8T82lBYu4Hs7n2uahtRq906Bk7aPn7ZsmE4LGEYwN1EOBmUQA9med
yReCVbXGQ4IFUOVrl96jTPkjAlozWX7jrUSwX0ez0XOJtp0mn1M7M2/9vBiGzmqZHS5nY0KgQypT
bJsw9+0qxeBWoSNHcESq+DFbzS0f5j/yoAKwAyNZT5vVFhsGJt3gdrSYiWSwTCEc+79TEH+35oB3
P05rKT359H+aeZWfVuf5Xqu9potFgXAbrEzHuU3k1x9W2WbmGvNs03gJC2wl0/R2xSpjeVJ1QvuL
4zvMjFYRxkBmC3gvXI4YVpennZNZJjvna2yd7KD/NgM1Rs1aqHdlgzRAGZ6nHprYhBAza5BRP2b8
V0VGHowpHNlU3mgkILai9sXQ7PLT0tbOtgvTkano/iA3tmNeisB2hUORmn5/yfmJ2nqZUUwH5IBt
Q5SMmWEGGoxBglDdFm+vUCFbFD1eD0JhTuBhpSGVTgH5U6QgqLmOjtCzGJREDxbXkPoXc7bzZfUI
wE4SpdEMFE1kXzQfgCl2T39sWjoUMB6RHSOyOvJ77gS5x8Oc8QAMFAmkhpnTvPSyA1aeM8AFTbns
m9W6DOrArqOCj/lbMprmTvguqRbEwLBgjZfFRdZLOEOxZWK9aB+WPzXA7oQTz9MuEAr+Xyq1ynqv
OT2UVD1B826xXfOiXm83pSs68cWGiinYf1L9yPi9M3TfF+frwKXLJZaDYgAT+wv22JxOulu9pFGr
z7pkU44C+jdjwP/6IRKDdmE4xDMnDYq46dzKntNSZbVY5GpbsBJL/o9VuoyRQBtEOjsKtZbsY9z3
fOW40qFuMOIHenPisfJY70YkXmciJuphDlITarKCnro/SSZ2yoL4SDahzJ86Z+R9wNvphpgziI1G
HII//9LTpA3zXAulghv6O19HQYdxizuu0IV+HkS6lEb4Q807Fsel7vRDD5h34v6UdbJoD2RCGjxa
KG8lHD9zpVZ1kdJ7EzaHx7Xgbq3TOgLPAT6hJex515gsucaJqXYNC2BK8Cl0cIBCyZ2vsZ1XHbuP
OOdPQh5cj3OJJ3AqbEGpefb+ihXHi0/l2dRd0h+wj9Y4/PZ//mJ0hMSU4M3VRzbGPDheljfo6CCG
nG8pE6tyH+umyqZnnwjvxH5WhVB8O8MQPCnaRNNqOth4kRdrR6VgGQ+gHCuPcDo36C1aW/nsStWy
Jsb8swED9R/l8kTBjNuLuYnVKiUKuxEMcr7qSlp5fBxsaVJywUAljBpAzRu8nnDQOagO0+YHkH8K
8OX+w9CIkmt2GITLVgqdtRsRCbGiGPidJ0mXa4wXWGu8Y7sDp2q5f6P8qIN8ln8v+TGyNv0Dpq6X
LkckqGZc17VHZvKOdgmGC59B75KtvocNL+yv89AQzk7PYVeJ9rHwlV9kNbBm3u2tRYVorb1GuofS
di8gn/Ipe2zETcq4rpiDCS1AIGkUBBOUuwpVIOJuWGaGYGHSUA+9Mxu09PK4pEeyxrpJMqHK44w6
V9lA1GO+oYCrH3tBf/+k6xNS7O47g3OlW1osj/+aH+ohMP96uJtcJmR3W2qLDTXheW+Cr/rg2O+O
YTE8V7JOLOsBsjBhyzp/+cze8uc0RAdjodUPBjMneOq9Yb7o13p+VVMm5sXUPxdxE2Khl/fN143x
HQnk1Sv/ESxu75eXfPe8qeAbPIyJq6T6MJiN8wfMesJp33abtxpzYB+FwnEvAWJ91fquoQbgxTZn
QE7fNIb7ahq36t4Wlt6KyFKU1RAn30gXcAAh0n6IYD76WFOhbATmxqxZ5ZbKq+Jk7HTkrr0mTfQx
qI/xFt7ZmiJrSdap2KRD98SBXU72L+IZSutfpX20ZBOUxBBquQa7lV56eIFQME7l5b/34uW9qCXV
nEeZYIWyJQenSdSyxBqgarswShjwjw4/xKfxOxmbDFxHYi4sjSj8P2JNLu3i6DXCI1UiFnV/sV3s
L+d66ku47FwSnfXyZhBkW2mK4mFIkyCjBuOvYAGeuB9m+rE3E4ixxrYcEizyxz17z28cmopZWzf5
nOb7PWz4MrxIio4F1QUq712FNg0+qblS0rn1NzLCg7JXLCSPO0tMOotcDq/QajmIF9RfWRlANSp0
VGafQnQI4VpF4OtitAby1/GTZTLY7wejFOaQB9Wro9RF11fL6jkimfT4m9R1SOdZcQlsu/PiKZdh
+sxp3cKbvjqZwg/Z/uoRq32OISwGRvmYkhJILkLInXRAQozCRr8lqo5hHQLf+6ZSssS9cV0AgaRT
lzTrrnXFY0Q1OPbfXozQdqvqUoIBG2yeLCXNMGiqRtRw9cX5V1Q5YvshXP05MfyoN6DE4J0hKuLF
4QPIi2ET204KKKwkjPxWMSgtZiAnjCxiHmpMW5HRxxCvdEZnafRn14UPGilvj5l8SIDuY+5oaTsi
dRZzRljBPSDChEnNN77vVFwO8Flo0OwUd2Hr93Mp4Wt1Cqu5kJh2z4tpjWuGtm4uiaeiLykEtFIl
7kUXWTiGkh2NlnMLTELz/GUi/Np/a9O0DY17ns3mxbC0UkTfNSxtIXW8NvuaTxOiY4ZkQw0qufQ0
j1kaup81WOfVDIGV/YU4dXhc6DL2uC/PWbxvPf7iK6eq15lESdqykkCuCaLVyEETXQpOe2b9uceY
/su4dn6E+Zkk5grqXIkwNRSaBabKEZqHV2+XprCtTQMwOMU6q6OlcvrgztAnnZVV4kmpNQokQo0m
5S0fDX9pWHa8ew8nleFrmwDYsvoEtlB3zUbfyu+K/T+va/s9ZfRjvg93IUFDFwh4ecTQ7d17duMj
fSMv0U15DEN8ie4EeLGqtZ5QVUGKEwPI5lnZTTC7NY7yfcdqRh8rlrJcl8l08u3PmZOw/msTegEY
WNVAky2FF4F/sWf2v1d2qzfkXii+u+yQmv1JxUndlGoqvhgAktdbFh9XpDOe2BEScXhr0gk0JAXl
aQKd/S4oPxyhkUdk/JqVFCX7nfi8sst56y5+HB0Hnw8arViX0K61XsUWLwYa/OpUpPD7TKl8e7QJ
egddL4oXehUFyTgu7V40Z+gWa0iNeeseiZnmB9l3lxSFBJr0XwbzLeGOnnbDybS9UHRPltsHBna7
GKqIGe0yFXWfo7JBwZIR7NrJTItOpCihywZ3a3RsS9HGCeQPrwEAHKdw6li1sDtxgT9luG1MwoX8
351BdW+2XejvozpiSFAXHK1N0WFvt0AL/6HLIHDPWIHU4WdiNSA1cZod240TPbGtlikbDrQTVr5C
9X+iKquITX0oQ+81kBB8mAA7cz0/APG11vMvgcze/fAQ9971bnAwgGSI0qiyXukzhqt7BJ6NJzgA
xWwt2qMR+zoY2ekB6jHO0apQ9sonuhQfjXLtmSaYnhLvszG/LTHhDx3ORNp4TBvzdwxSqhdP4aYP
q6Yk45SYcSMYC96ZncRKUpA6O1EVEhV67yfhBKm77qbbmGo8DfqaP8ldnl80BOeUQdui0dLn134x
CKcY5xxpIES3u2v0fdddGfhcrRg3dPW57oEKtIbYp+VD17wn+YDUaXHwBjT4biPlVBGqLxfNdhtp
gMnl4juZ2DfSHyVMMelQQLgrvOz55f1YwpWSTa/RzXa2zW9S0cZa1vuEfoFhf0amEOsAQEQXcSpJ
/8au9BLeEFSrskgrhtU5qSrIxXrdtradxVPgUvYPwBYMOk16vMaIIXDuZdmADTCNX/6QNdR3MAq3
ykfkS3Hx0DvcTEGt4/MzXcME9BVj+NNaFpOhLIekA5yT9MKddlWTmP9AyOLrKXomyOzlSNLyLvSn
fWsHLyUXgCfFcTVBBvvCCP3FFKJzqSq5tNakV33jCmd4D7qMQ4yWVub24AjdQ30roeyOzXURPIJq
LyOXWSCNEbd7xPPm0RL4ySm3oZtvPNQKMr1F5qnlPPGHoTEOWBmFmP8A8OfF8E8L/uJWpGvCZikX
62gLz8jAvZO0aew08yRAtHYSyd8NgRjV7WBNd0K08SnS5d50JFG3Y6XpuTJjqbo32L3K1xos4uEH
qu32f7s01ND/h9zFrjWgqSOWs2XliyRIuRypkMfsGy5lFjKm77v81JdNdeR5u7djMnZomsup/k2+
hdisamYdojaxXdTkkgf72rPET5JVXEkwc06AQAIdinl3rkm3ipW3OOTRRuk6QqhuS/+mke5UATs5
xRmEsoSOQlcRnrcbD9PohKbeZWgbtjqLAjNo3pSYlTRV24sEZcSy89dJw5hcOLYT0vVHuuldR6L/
fx28IH9PBnqrQtI2mCR2cfcZBZ9/cFdFNaeXAUmy36gl6VemGbDSNsz5YawpyGmZ/KBhwjAn5zXB
mlSULimHIBYbavSdXD7hyw4tvzs2aNATPFCWOUiAuwVRUnAfARo8YikZsSw0gFU5VoIeWNZs4mX8
TKnfRegr2ggUNCIRQfk4/bAmQVw/27QhkuCIHgzAcK7cDl2UQqf2bVvBh0voFSjroEouNpBUD9m2
ZNKf51vtO22uXytgmXOf4Vl/Nlw3onm4h4J5q1GQXvQMStZMthcz/y1vECHhoD+LG4vf5YfvUaOw
t1xqJ/K7jSsxvcPLRovyPh6lHjlnA3u3pwxKSdCuiMU/87xAk417I6tu90OZSxkj/6SHklC6nxBI
udi12YLmcxqMJYlmSy4s0LIE7MTdZRkFvbiDt7ViN+rvT+HexK0TtJ8tQCwAUtImmlQVrYEMtYAN
qQnZQEo46jvkfWpwXNVSp33HJk/LiCHoumDTBIuGJoNdxJ2gb0jJUsC6mAg2uMnopk1dayHURuv1
9p5RvNVoyUmhVKaoPc58GeLYul3WvdAoHtweFn1wL6oWvOzYsAgAIIQoqgMcInmHlK+8L1Hpt9mo
pXFhAY6lxGmVqQ59Fkf5Q/oT8HZwvjw06DAqLrlQCWdgzDoxcJwzkDyuc+VQRHGTJ22INIl8icPa
VkLVi07ASD7gHW6bO0H490mtm0+36N9WdXUAT3oPHXhPoyBUo918QRErWPNbVsvGXN/re/c/y/UJ
4BnkDPysokTay0/zp2iCaJMGQPvtVhgLqjV9SJTktX4mWIX5vQVRY9BDlH/+fyAGxdP1rk1i2fIC
A5chdC3mK5XgcF4T88V770BXJtl3ghzhcrnoSZh8MgHFFAkZbrqUrZwTYsQTqIrmrqFhiFGvX70a
H2dWf6ZO6+4tMFA1n+rdbOJoWhlwqG8O/LF+qnblQUBCht/yYhAzD3JR60YLOOFUCknO9AqmSg1E
EFd189IgglqB3x9boMBQuhbxXVk2vIXC0LoIAlSOBAyONIvuabHA10VElbOkMgYRminWgfTge6lk
VkHbCRju4fFP8dsd1kepEndlPGK+UDSOvgixwGFKjYmXq7R/vRLWVIRb65Os9vwcn3yai7h48ENK
2rp2Ms5fghJu1wTTREG/fXYQMeM5vx/OGhucxoqNaoF9JouC0vwtEUQdJXH5SS9cU0vHBuD9BcGq
Hr4gnAsBwnuHXA01LbhHfnN382xN7sLTWJ191MUO981FVwWiHF1S1q9MtUJgpONxgCtE8yLjhOxg
eoh0H7lr9F5hSA8zsoK5e07aGqpTWwKS9Q39sSkRQHpYTcRHLVITvyBFwG1fJmnxNiO+SEsWdxYZ
cU4FB3QBYAa7XeiME9GRmyjgdcjnvTLeuumkFUpFmklDbqC5tTM7aWjs7b2b1XFTh4rShD6exZ32
vro4+qkScFfy1diCXaYykG48JDzAP0Mqrjjf09m43JMttqWP2NronDjnSVkkje99psDHk89MNnSU
c+Zv7gzgGpqvVPYQ7shRGYWwE0wh4KfS+wt57sO+Bp0HJd0JCY9Ex4mF3ijQQNzOSTdZlXJrXhAz
J4bKbwKqX2910nf/DjhSRGF7v2lMzeuuN7HSQrMCmzVzb12YU0QTuzS4kD0O+cGqciWdX01XtdB4
DUvFBJdq+zC1FyVQ3fs4KCb3U09eurhcExU76D2Z7x/tWMqn98ydbaXw/pj78Qitp82jZ2SOZSKC
ibIuVwL1OCHpjfeJ1YLM0Pa+Q88LbbqbEQjWAhEKyw36tUFFlkJhdQnAf46U/QJhOaCtaD2GZ8P1
KV7BJfxUwEjmme3Va+CRQrE48jGNIukE/eJ3hItN/0yLz2/4PEvH8aW0DkfujhRfStmaYjoekaBx
MWSECgAhVvq++aytd9H19dJME2BFT77RzDwaImaJFl6aAXbWhSl34F/zmgH+pQrPxTt/dOJpzgP+
1if5EtAtoEdihGHr3J6GKiD5RxvHqkxwre+YMxQzZ3ArKoKYLN9Rzyq6EF2CdtkqDnycp/Ii+QMt
aQgGe5DEPOmZyOLuM6Fuj8rkY24fwPoFKK6PrNl/n5AMCNY3chaNajFqWA81NxnQIyfwYfEEUTqQ
XZhi10CLqv+zYrW51dcuW0wp8wv5opJkZl4Nhmktqp7SfEOLE4Ol0r18N7IvsOVIXwbJy6WhMHn2
5aekOfJtBa493cudTF6nxAhXCacS76eC3bbKLxivb2oioFHFFhqI+JwlkG6ExEV6Zg+j9vQdHOtT
1mZ4hD34rzOyXO610Qx+vJuzJx+Ud/V/fXy4EZ/dQeKtDd6zxR7uaOI/uNvyCeeKL6qVaGB8YnhP
/Ld/n83XXVD1umaVX3gkxoW6Eg9rqBC43uIsU2LdymtVQi8PCQ614EnU3LSSI8xnEImELH10Avur
GR3ad7Dai7gZuwOv8woxMNQ3i9JBV9JLewnoFrv40wyW9v3TmA0e0Pbqko6+U1q4hR+JioKzHbX5
2oGM0yUKf91W/nV1KokHSQWQlpy5EX9taeynnOgayREUYMu45j0fGlOD6t7Dj0TTSMecct0GO7Jb
ABmwA5oR5s18m7gwtwNNLCJMSmG5Hgm/lbo6CfYlbLdMYAro7gPhcUl2vJ+IL4GSMgFcUxg2Tuup
IPHuekt9Erirp1FdsW9a4zi+RigOD2l2oOwHQzSf4MsimbwiMxfGxw+hnco5uIqQGpTPjxNIalcQ
DMo3OVPwnOusajg8+QE4jh69deUTYh706vovvkZQadj4/+z4gc351Fs59EGapW2tzu0O/ZSeiVF5
35QMBiBq3PJKoOZQIqXxSf8d3r93j+gfz0ldZ4MjzvpotIN0sNUW2R0GeYmisClA+ek9SFU2UKDh
9Uk+R24/7RMZKglVzXVV9PZVWvYnZ+smgjp85ZAITKBU2NGWTb/OQmOgVMsB5r8rQIKCMZrwmsPp
eNuPruoI0nXwRHvZYZj3oZ+bC5YTAKRLM7QRzjJN13wSaLxkQuYUKbhOXaDLniMn06f/3y/wNTxp
jBaFfq3zZyPdBxDaOJi140iJaXrAMrg1I82SjESCXlYx0ecqyjqAteEprNkbiIXBDO+XADa3rdRp
BQroflT4y2y4RbSxluf6m+2lWY9twZqL3GFQsOYhDGdGR5Wi4hJew62vG9Czo1rWaeol8OeOFwoN
O+Mj59K/u7xoYWMWPrsRUaeq0rsf86GvDGFkjfhPlTFhA6cYp0eyrlzqYqCLdkdqlDl1eQ+ydnSt
xWX7V6b7aN8ERoMgEcSCudI2IEBYQmNk5B50v/C+gg3bJWHy3dd1N38jrDXrFbR+97RoyW6BHP+Z
Cd9WsFkZzSbdumqzSaHRBm+ctQ6LRECB3hvdt0tQAVY+BKWG4tSWN3wJs8TP2C1ayVXHHgDIQK7J
qHhyaayA7IeNeUsx4CcMJbvWGhY0K3nJSZanE31NEu+pvd8vDUjSRgymuTyOkGNGSNVZr5RrywKU
bhCiYuW+KotH/xQTpSEj7hgB3VL2Y4wSWg4Z+PcSWcRo85r1ULLBVPUHXZ+dcYP2Lz8LduLdQWaA
FQ2z6dB9JCbHzjjO1Ei4LTe8+/Nk2DGnhDupC4qvYbNslKA4kd/BQ8Dl3kFSQ2ksv8sxanWP70gR
5IdMv931NRWXHFwXFsYkROKq1V3yp6ct6IJDLeC/y8imIki6fyMhnork8+NRLKCv8Q+Z2mF4FBEC
P9ggfc4+jTL2Y0Ea9Bzeuyjo6QlhTBD2gtTS4CbWlDdLJwgAGu1R1WqCYffp7bmqLJQYO6riJi0r
kPeAzyIJdRImA+/DVKTrX35sAhyHfISp3W5u00aZXrYvscO8PCAnxGChw1ylNvlpVhiKjePqrczT
ZY7XiYzyUmyHXMVEgyL8PJ4Ub3Un/M+7vrKqWFbOxW4ofci4Ky91oQeOUrAwkmMl20H0oufqiYQ8
zgiLngkLU6dtOScxlVqoHwLYXl4gNZ8XTSvLgCrGQVyaKr8Wy3kEvrrjVClUn2qLJ17zo+nJtwZc
5tEDkbCrlRjyMycuSLFiYxyBNz19emrlBMeUA4pQ2MC4rYuA/DBG5/8/X/c+0NXOkQeVV3FxQSQZ
VR8+uFlyCdhLOxoe+hYkBHkhXSo6lMFwZ9hTE8R3lKtbPzdSUeQy+uQlYokTr717PN3qZETGxAEX
PUXNpNy8I+0gIP8kgfx9oxk1WEm3zRJ1nw2xiuwUYvxZWDHG2fdBZMo62ISIpdYDCTpWTCLUqAu3
HthWuxpE9X1TqSsu+L0uj9rK8BWNi4JJSDc+U2Gl3ku1w9u4WQFBEsgHocOdMFijWQ+6lFYDCHl0
jFMPmoHE8oODYk/2Zc5FJGffYS+8vjxR3Aaz41G+KaiiFnRXS9WQ7c4FUYV6z7LWnv72GhJxs+Nx
GHDG4TsEWPSmmzNjCdyEwYzRxPYm9HC37D2UuIrWxnAqDLe5UlLqyPWiZzA10jiY/X9HBXfprTTJ
8giNjWwBZQLPj5zZlJMCkCkHzTmUtWvY5j0vjJCk9I07xtVlszbMuj67dtgFFk2rnPNcA8Qyhq+Y
mYuGC4y+bBb3EpcOSzWCg1R0gVSWOQbH8HlXYDlLdJXsndvzbKI31JrY5Y5ZXrwjIjZ/5RPeRi8v
H0QBfKuDAGFavN05tqkcRNQ0jRkPA6fMoXJXnISrseqcn13eTbNcgZQUFcQreJ/X9LRDNJtWu4a2
fozBP/9wPqRsVnLHwXA33+veq8NF5y0GpM92T40xoR7r8T0EDA+ssRV16gQRbQqnHBK5pNX2xnqQ
eWJGTdT5Lcsoo4qdXcn7jSazOxJZ1aygjF+QAW7wTNtOJeoBzpP74N3yrzAt8iJgWo8DtiemoQaM
LVhNjvDr4FXNcniSfeqIxL3rMqKTJun9wVYfmPLsMH0p3wTYwEkNXgxyqemCnXfUdIwvxFkBxtr5
vUkRLlFA7S4TrJIAWgOnAkBghK0T8DDiArO5bmkNFjcxlx9wxX+JzYt8FddDwaOW6D3uUScfyCgo
XwQfE/U2AKHErBz97lMTQ7gEL/wkFvKSE4eO8GcfQdvmJQ0IwgOXmmpUAaQhcxTDecfGAOQOCGJA
DChEOWbkCJvpp4N3ymJpv1zQhKAmP2R4kqw4wZ9X/RZ0jgut9P6Zr2NLgAgSUlEKKreyWpVDRsSm
AnfZMvcUWyxXQ2ZIBNcz4IGqE/WQZkYubVCPFCY71xkmBkLYaJODHBizLDRxv/fvJEdaW7yb2kFE
PB8MiyePGXiO4q34vmkNczAHKC2MDcLDqDrHuPP7vc73ec3v1zFQPgqqh57kT6G+54qyCX6Gw25y
aP4Sra8jBhOWYx2VyFn1mkDrtJSpLudrUqr6TZCIniwMoKmSgGXsExrsRhZcaapTJDol8CaZvcRK
8kHr3+EWSFFxG81pKHwjJWwsmZH2Zmb1wlkDbWKXWAHvEf/AZWeNvRmIhXqcN0oXzWFpn18NmGrv
kjjztnPENzTMKsgb96q7kXfTrvIQdODrcPczh5KgtuAxZWXk8ZtTonWRPT8Oj2WrVmem7Hr/4LtF
+b+s2wfKjDV2qdQbyi/ROOblfVAhC9KKu5HZ+w/SsIxecxRGUw0pL7sNKDi0HfI89ppil1C3u4WE
hN8P2JcOvw68/R+oWVB71zUKiH7Bm10h2GpLg2HmSg/03XthLHD7auk5U/VmOr9UfAv/snr3cNFd
M0jT4VopRTdpyOoLMQBNLAAUJE/5LVxOSoBSsZqioTa1b3jDGGI1FYenc5XZPESdSEUbRnJ3Uqqo
nYV0zdCee6wOZ5VPFHzNs1ehSqTErsOV0e3DNoJ66r2dBvNtGmTRRUpP0VXWAq024zyFXeuQBE4s
iiYw7TRx2d6/bxvi+aMyIb7vF3Knp5UqNb3QIR7KO2EVlrL1CcQolW0aPBOYfALPDXTIkvf+POWt
RsR4JeIf8JypWGtVdyDFyB5LpMgdlu9HMBqHburoYFYa/c2SCrVdJWlIBX0BZuAwgBSgTIlOsUQ2
nG3dSuO95lp+nV7ZHRx0c9/rHLnO3+YJPbWLXfQbUWQBkKFcpYj15zlpkie6KJHmHOAbTH9PMdM/
6UKt4mzlyNEXntX0QXT4Ak4pZ3iTXgcHA3qBkINM6/2g89hoW18ExtIpsSM0VaAFik/5ZTY0XzlU
07pdwTo/6KNPP/xCgtRK1KsdxmOFAgmp/C2n/sZfZKlIO17vc3iVqLPbwl7A+kLvsDSvPRMGJNMZ
SmQ+Ks4b3mcPuc9CgGhJZVaN8qdSG6NMO5/qK84dSzS3Sq/pZVyafRqP2rNeZcxIYzNe3LJbNiWa
YbNdLOLi4nD9T0OCAM9S38rMHWnWMIGP7kJ9p5t58qTLSepsaDDg8oNm7HZekWj5kzFHxNwTJSl6
tvMvyBny5HfYMKuOMATkeMwjcAPPZwl0jEhmQRB0YqlvH6H/aVs2B16+brIyWejCG+AE9p26UdXw
Eg1Abzm+dErHIzFzX9A+9bIBNgLQNOZo24Hogxn1/+k8O39EsEVJe57DyaC2aasfY9fuIdAbUf1e
lAj8W0AU/Zb/I/KxRfPrtFQlw8azccuMUcnCh6f+LjL+JBsrAHPN+zv+gLISCPxsR4xygUfrqVTm
3m+MZG+jLe5Z3TZVmyaAiW1BIxaBF6YtNq1PZtRVYSv4FUkTTzNL+BrwZf2muAMM8xhZna5Mnk+h
1d5Imjrpp8wHL7PQQhG0BP7BPIRnQa0U58/J6eDd3CJ3DPfED743jyvWtpICMiJE0CbjfU2j3wXK
aNX+aytkxuO4vq+pKlFHvHVb4FX58OFA9cArW6yl+bKeKORloYAOoh4WNQiih/Aee8H+Iuank7Ax
C6kzXHSIGeykdAixbqmcNGFXdYlz/Sie9A8ekwvLM7IJ+M6Q8QUL3PoFggK7+JFedVdh7IcB1dKB
hrB1LI/HMJFyO88iGaMmIA+/IUl8WJX3pwYU0wDLrNAZ3+F30KhRW8QjtzG8BsDi8GCaezn18Lym
WkeqiaFPymCPRtp3XU8kyRAmBvbMJ2sCOwVKbPPhBtYXfFwNT5JfnEcFYGpTPIY0TeU1ed9EAX1K
nFwbBnbOi6ylB8fk0f6o7p8PXKZw+x87VWvWhraQVWPQ/x3KT70bsDxRh3fJ8Y11mT8ofy/QVD4k
pActgmef4VTZNmzKU0weyNrCp9B65OyTFqq5bZ4hhtUsbNV+9Oeo7hSZOR0CjFuK/vpOnmZu5PyC
lHEnwWybmc4pHOlVpjXa9RHtCBuAPyjiTydu52PamOciKzPFmwLerbZ7CJLcXVRx8iQGNOF/XDvn
nex8hgy98rmfDiU1m+7fIBCekAYY/uf03ImtPH56rAVoRmDBTtGAI5K5ig60tcJhhX2CfFNN6Vo0
1NnrvY6K0Hm8jzZ4+cy5m3hVESn/6m+VB9xn7udE64ZFYgcdIItVw47ViwEgTSfpFqoh/Bs+OcwS
5wA5FB42b75rwHcal3UlG+xgkHbwK+3kZ7l+GdXhiafmQZSTjUwcRrI5aE2Tvx5p24BThDLN8suE
PvX8QNnL2ZjH/Zg3GDc0gEzczEVbt412AVhBpE3878WBVZ3yG1HnGcQ8sh9ssscREghH9+cP4bXs
vBpffoDsVvHCqly4qXaOQidTbk1DM60/09IFW08Nf0a9Lb7p18SFBEDb92+3pOvGMNR19im80gTy
oG2SElErukFiuSNA/To99JAqNG4WwJgZeCCRMitHaHw2opnjoqEM5jU+cnL2j3g47eA9upM0EDXW
ja17mHGRV5MWUPoSWXPueDlOo3L28kE3tsMJ3QhRKikCHnxXEnI5gGGtak/jZZCmDa4iiCgcnd8Q
v4NPETe4WcBBp9/3odJwW4UoC4dtZmsen1OcYwKZPn1lUPoRlBNp2UpMl+1RdRpXSifIVIfg7Sxq
rgoL+MpO9P3IDHofRsecEcRWy3pEF2+o02ieNNe54ByXLfr3Or7NRhlwF8AVbkB9ly6vZe8tYlYy
iuFVfp0daL+fridSfPJ51iVSuLa1DAlN9J8GYbIT97tg98v3Z85RJ8lm0VRJZcCfD9KN7nhOgavX
Mqb4EscmQgfLGdf3sPyFN4RajRaJWbN0u66CUkFKsikIpDjuBQB4xxgVTg3EACiyQSeXbil51auV
8rw1G/uRoj12v+zpNbGPeI1Enw6N5Gr18jGjZnpgZC2TNlKSpbhgYgLb9zCRizUHS0MLyDzdZ4qA
Wc8g8u43QXU0MIy4rsQm1Yovoq4go9p5lnreV0rE2uUZJmWPZ4hl5hTnubSzLzPXA79DtSBK4b0D
ekXZkc6XpD89HGLWDoakuJpJeChbyXpqLfuzzfr/olPvVPfeKHT7O1StC6buQyuHC35h4kj83dha
rcdYYukjZulK/LEc1ZZ5dMIUdCY6kITUm3ZRV7lRnIHbL5zurni9uno/9m68m115aIEwlgB4rf00
SYku2QWv1k5Jj5Po/tV8sZW174R+plzC4LA5bLoOcy55bI/jZTmmOOwBp3ATqZ1uP9X4ydX+mf3a
MhwWX8gRQj4lQollmso/KErqKOIePBycejj51D/LHCff4Xaj9Y7xDfiXwLdAzEfzdYPUnn1TJKdQ
SqrZnHj5dr7457j/IqoI1eGaB+qiGHF89jwYOA4Uyqvjl+Ssp/o2okuV2fjc07GZldV/1lyq4kDR
1b063y3RLrBKlf9iAVHX0kFNQflGXsE/sC78+gX/r9Jt+A4Ayaw351h7MpQdbHQkCDuZtlpqP0JH
o4WLQrZ1NvCPdg72QbH1xxBttn2P9z2eOESRfPsfaEKStiiUCQDybnmlA+NU7SgdgRWYsn0cfYiH
G6i8KPHZuk1kYoyYvT5HRaEBaYX7EoIgO8vihRpc/ei2gFAoXuEuje/pxkFZ3q2sCkIFwR1nlWxz
XZkm/ZHdYsGnhs3ViAaMx+07QDEUVOPhaQ2jph3MjnGS0dGLio2sug8hxFSYmW7CODLlvD6yXeil
dOCL976zNuYjGWQhQVgNOHLuppcZ5YpDRWvQ8Z05No803tH1Aru2RDTYpu2a6Cb+zSv7zsnJFdJ/
I+8mkzudiU6CHj0qeP25ii6jCwZ+EbYMPh+TSCbeb5Gy0h7ms0/vCOQfZ1ZdyBNvWr+TG5vpKpQY
urj+450RsWRKwylDFjuIJhcNHB8/O8Ibdy2qh+5rNUH6AKxNZ16MFXG5b/a8CJlq1RIY4nJfGbYH
cwetr6BrxON9FLMyN+5SxLSyb7FPQPktmAdnbT7YcjbFAeCMQznNWqQZdRglimBnJQ4KxZwwXuuu
irxGdXg8g10PNnbqA2mu7vYj6XBcG8CALBRmnazqHXi/ivnaThyo9WHlYluW4Q9SoY1dOxzSzziI
0pgiO+UKjbK1lbDlB/+sk819+EsG9l/lfGq1PI4rj9DnLUqTXO4TXSkxa1fZpSsC+WzYGKdomisl
ZglmLy4lvNOCnUZ08G4ogK1sTX6/4HBQLj04ZQHULnsFvv3FrDO3gIJ0o05GL7m/Dzy+t2wUfX4z
sRcGbhkLKR2dkpuI1Z+EBjX91LaaxGNMcuO9wX5h3TmPT9uNRclM3w+kaMh5FZF2ntE8vBOelc0q
AWG4XLLEkWjLuvaYCH0D3i26xCubngtYC8nrdVrvVWceonE1oryEXXvgDVIOyRvFKw0g6KX/05Wx
UKA97YCAuxhwgeCu1ogUqZxxjUlbe9qRQI/mqxcQhTyGByV8NafQpHxPbQ0SuzprmxbaVynr6MJk
NEpg0ai6hzhG1UfleYu7zs8TW9pLox+M4wy1w25Qsj2GzvOhsBUvbdU+uSBQqmdYnyz/1272Tt4c
4K09t+smpoc78MYpRJ9FuZvuRYIMDbj/EzZPILuN96fDno6ugZHUEr8cINbjGRM690BzgKdmP1Rp
wV0WBH7m45d2M8jMjuo+yUOiaE1G8jdcciCF7sUBMqx0GbaPAKp2ViZIcf5VcMg9AtJ6mrNL62WP
JAvDioBZdSHrgqWQ6vxaCongy+fpMIo8KT/a0dhpq4DRYT6+FZY1skehjCJqtZYFOKzm1zJUB9T4
TdmSfpeEn90qdpRMHphmaK4QnNZm4vOj5lpst0ACxlxLYgc9QOHcHB8lTwouO3kpszsEp/DPYGSX
hoZj1S2uIUo2lQcSWXaTXiOPwUOuKPhakdRCoKYms4QPSvA854R2/roZdzOaKH35KDJs0WsloCt1
tEsyg4Y6+UaUYx5d7ekUP+nxgbXeEJhweMvFzsQO4BBdc2gnMNaVGitD5HcGytjq+mjnmdXOJkhe
Htu5exV+0+Lkg/WcClWM2x+BRKcc9GSYGx/BFD2CSHyzCldPAGYi+GI7DAPhvkdCHCHOQ3GBDRHs
j96vFQwG6/UZFs/3K43TmRtBPQbUOl8p9Bn0rH9ScHospQZhv/llbYbbaOt05ogG0TU0pka9F1yL
shesVMgMiMw+peCf26TkSg3qyNeOqYzikheh9DIygs80H+u+QF5qFeBp4L9G10UiznSWCCX/T4IS
iDV3WYMo5phkWoA9LY1x95omsPGnfzz6/SR2E6RtOhNggy1bFZQGtTWt3bVkAlSGRCnMOZUOSufV
Eg0Rsia8ThxaIh+wLnUabeN43LNqeCKfwG1pbm4yGzk2AymmNJDqMSaOHWPI9Ue4hePllPTqgZ03
3WjHJ4836nLSnj9KGqG5MO3fDIvbTItJpshcYYACIi6yS1cMHiv3qTH0TpVWxO4YJVB46MT0fW9t
zhlbPcsifsAXEMFYnjxMvwgsIy16i0BwTL73QV2FRdXtehdLMjMXgqqLcU4z/zM+QTLbop8gcfiq
qn+38Ay653uXWKMQ/BwCn9Ik1FAmd79b1u/viVM+Hkg6k/fnuJlXzebej5mhYg7HfIR99XT6KULY
ZMv3+vJ97xZbD2MuYYYGy6beY8mIHo5jolb5YAjoZWq9HzZsX6VNON0peZeoSr6laEP7BrwKu+lQ
WzIIAb0vf022nOf6Pq4fibZVA3Ib6UxgF4eH2kcc38fkL+jTASGxN+uQaP4jG04uJzv7dMhq9X0D
jUO7dXfehSiTVrorGubpuriXiYx0NT2z0Qlj3XiyCMFPwoccWbgPjhc04GZZDk3YPDcarxWb3gei
33+b9c/KoXTSCyZiZf2dDBEbHxvdVuu+8DCyDhsRp8xOdOGy39TQr5vuxoIV4XVpzpycVowy82iV
1DRgpD2PNuGwtXOx8lNkHy2Z0J2CB7/bmOkSZFke77BQBOwnx/n+jCAw1StifxDTgWKFZMV9At2X
U3teOJy15NEnkY+4CiRw9zRk8YwNE2+hXKeK2uujoG+kjjcho6DbN1/BfkwgTiz2YUqc7eTBlZsq
CL+rPB+IbA5sN526bZnvPYsZBNatKi2FkyafAheVNAVEd8G/AVh7fyHaIp1EhiTQ3jKr8HeeJ8j3
Hq+CZ36La+z1kGsgJlzew71Rwlo1FaXjjbDWW3EoJbz8/J2XjXLF+R+nQuklK4/vph8NkaRXVAKR
8jy85OYnWplarWhnzfN9PmY3qW/2/MlhsKtuhnF6dVEs6sA9dKn7mQUDjSrci3ysbWPgNNf3UQXu
DIFc7BQIvfXjMQLaR9XCRszBUV4ohiOLPUD+GJhocjt0uQFfFL50EMvpvlv3cNKbGMgGfEmIXKtU
q0uMMo5Ritqek5XeUqsmh3O1UBPng8EZijvoXJt9/EN8ewvKHGVLQWIbhHK4bSoxMCt9UgNbu67U
SSnkRJkKKS9BUXs4obVNLvRrAgaR5i/FLFIRPjoyi4yAsWgbxU4Rd1JjFH+y0ZA7r40/CqlONkHg
CjmTyeNNVO2wbKCsjGha8SIXMFNc0/WZDcaCh76QtZPyVye/aR0I+Bblr8dra0uQEIUwES93yEz/
8f01JChD2L5yWoDqYT8/88IFA6dFyZxNoGeX4CqYe6w94pTrAqAyo8YYxcDraiAK5/un5L6fnSk1
uJYesMZOxVklTRVAYuYILjcVzKY8pmfmt6J7gGSivv4kjRVSuU1WGeNLE/428UBuxRwj49V/2cf8
FoFzRDSgDjqvQ7rKnUgEkNfPR0Gmohs8/Cc+jpzxhnRQzRjTBpVamPC/v48VL+13uw3aaiM8d/fU
ae8OIBKNDw2mAQAHltV8hcQYBOw19Emlbwbpkt8/MWqYXcJ9m+3MYSgeFe7ObKsTqVWq5BvC5PW+
dPsyDoR3BguPER/whyY9gCMi0MeE1A+RahH4pzkhZIx9ak3fXW326Y3QRQTgkKmsWBDQ87GBZxF5
gYzgGllemAWbfoTMDRfK6LImk8mdqke4z+7kpuQJQIJns/QRL57xy0MTyWJ9yTHQ2jMWXQ90UmeO
Rbm00VHKzEppWv5cCGUmoNJKrP93ggiRn4OWoXyO2+FSDD+ivJudbdRAVvwX2h9fJsL4yMd5Bg/l
wi5c6NzzjxJ4Kj9UBQNb8UB/8I3d4P/DuAsX3LCTYE2Zx1wEIhYn3OuyjeKiw1yMwqvUBQazyte3
/bc4aPaCn01tqqBte3xfeiSgxXjwx49F1iwQkhkNTGJflw2O9fQD1MRZds+fN8LkQuyy2buVTQ+7
dY0FgRdwSBT2Wpk8Mjnn6ikOLkhVaNTthcK3kO/eYOFPKuNFZJtxZuMpANJjxwjFcMnFY5ibdAgp
fA/RXqfbOF+2TMMru7t7WQWlC72S4GVtbJHg7fVWp+EUXhkQPbC2YUgY4b7W+T57ZdZChOEjC8ns
7jqrLjH4n8/sEZcWn4T/+MEhgmg7q54GAuOUpR0+C/7fIRqJ1SYWeYwihemx/LAMAytvl71v24Vn
rNHOIE01/YbXUIsiT0m4oys/W4c1j4mYNSxi6G9vsohAp6TtcTlxbZC8zt89uNBCPjmiTpKKZalx
anIk4eEGfB2Heg4ZXZm/660AW+qXeHYkRgdoRt0yk4HBah5QPuibEUeRbU2pYIRC7zLRKWEqOQHh
C7ujA5mwTpEY/gtfkqmm330d/AlMLnT+giBDU3x/mmyc/n5pY8j9sTEeZN152aMFhwLugn/ItG50
StWo8UnLQHIMfBdUhl5JzL2f43rtq+nMYsZ8tfKcttJm2hGV5Rmj3GoVNxFrm2B24YuZH6+kyYRV
cDUVk7Xo4mNeLSG0wwcdQ9RqW58r3LUO+VAuD4Qvop7gidfXcWX/za6GmjnzqshPakvSfgKxUZQZ
c2kzslt8q5qH3am898neZuMS9TDPSfjsiX8oHuPV1wVA98KkqxaNCEXVUtqnKezgmOLpkZjlIZdw
RdbkNbHXfkCNOQzszwMsQaD4KL0BCGjxYP0dj7U7HMBwS7J/vL6DJH5cPjZySP/i29Y+JKW6x93R
SBkxOmEq8AuKZahKnJzCsbo5i0z2epAFA3Bxz1bcplRzebJ8tsmH3RUzRCLYdm7JhggSsYPwzxCo
XfqVrVkiVPlzMQqA+t6qe1f0ZHXLbYWji1MzUIL5vUY3aWNJkgZ1vz3UY4QjalUwPK51yDMzpxyr
kfWdv6MRiz5h9vitCwhAGzoFQsVra7JQ8rsg9t3Gz4QT/oi3MKED9yRLMTNm4IFOxVZKmG0ABkHv
O2eVEj7b5qV/0fCnrP5A5yNuSUfkKRVe9VkpXNm5xPssfu8wtg4+6VnYBJAW6WW+z1emrxqyDY35
X5SW7kyX76T0+6XOLCJGNZswVJ5LRm6ntVUXMuI9kntYtOubH52jY80v1SRYstY8/6RXts85HoC1
RHkwyxN/RB4TnVYUEDZshjVTViUScRzT6A3DicQPxbibVPFJ8oc8+M5widqwNZGMF376uNxv9oVr
GjXsK5CESWUVxUYinADEEccT1sxdf8kDQJVnTftqXpyROOJyrQkXnSEq5MJv2HPvP1oJP+CNn7c7
UF1mj0DoLdmtc6rEpbnETTgQq7fwO5tr2avNkbsUd/URkEdKgneT9OshHTJ3cQuSPPc2IXUFhgZZ
taVImY6dMsewFIw96NGNco625IJV/67anrf4Yy+e5fQKa10MC+Jf4iOC7eDv1g4HQC6XJLyt5og4
veZVq7M5VSm5+6zPS+etkhT35GkkVaE9As5WJczMVKlenQg21eXpb3RNdFPhMOI2tDNxy1a5LID5
Gb2M7wf7ToyaF0hp7NLDp5lmqwgGtBiV35tHKz088585LcKfNz5O5mZXA8qEE8uVMuaEA1gdXEHO
Re1HrcLYeb42fHqIMpd38/CTFXaZR0zWV5DgQpqDbG+9BHyqbzpLjOwEpToOZ/3t8rtFKbtd5Auw
INF5SbPAMUISJqjtkrme32I5xXkJndumpx2imHIMky+ddjfFGWLw01EClf9xuUkFUC70+fjw4lLo
+ycM9J+CVxGfw0jexxgW2vjc1uVPTt4kO6xTGeZsp74rKhoCP8KXlQcaVxHn+n+4cNwrVH4SAxpK
W9jDBNFLiPEjt/A8AHLjea88SVU3o3ixgplu5bhMxFBts8hXWu1p2+AI+PrtOFdOjbcmzZlgAnx8
2NQ2ZdiZoFSnGbvFHuRsW6hwkSda6Ue93a34ngGW6STOo+gGXLMfTF3hrmI+0lFERxyvCGwGkicR
DvD4rmLAKWwyhx8jv96EM7hAcqRNbP/bURtYrn1LADw0/qHN0LTXU9wrYz39oAuhpG2Kk11HdHt/
KDx+8V1XDBm3oPxnThu7WwIstiiH7JYxfYPoNv174XJYLCqcPiuIE8x80lDHwfsaczQfU/ETNEcz
tvsz35pA8al0BIzYCbBao8ZDEN8bOuOACEfe2yYCoJfdDy0Ja7MDMBbsc8TWVNUn6xIfryS/y8oP
1fDtXxk9nmUlDUa1b3FjgMwpk6Zjr1BffVMc8koFYJexEeWkgAKIVuENTqZTE5LD8ZLeGhb/36iQ
Wc9bLirpmTg7P6b70SCMQoIi4XU7riNp5dI1gE7EV0LliCsoqnopbBQG8NyjzxsBBGD7dO9PsCRo
djPBneDWQ3qvF2diwwd3zXQngghDbTFF2x9XXdQ19XbCKVYqfN2JPuNqQKWOOGgBxL0w4iAGb/3I
zALRmZGb4LlBgmPzC9zK/AsePXxLCLZy+gbTcWVyszSfWIcUqdqJhwi1ls2xo5wJuMMDloO+wWDe
T0VSjtBLthXS6u+krSYIMxAoKjnf8SKmwfXmNx7fAPkjAagwvPeusq5PPgJ+wvBIImMQ8Zzs2UlO
DWvQqKBuZfKLx9H5KHiPcNIzPyPWEIYnTP7GmpANaQ0r1qGZib0ARe3Up8QqG8XKUejaeww6ZNkY
OFugMh9lRSd0e24J2tu8hfvuFm6cPCYGt2LBlN4h0TzswotD6FMe+rfoPC8akaAYRKp7DwpTXPD4
RoNzVIKrhx45weBHJ7HAzTfMR9m2sLMd/ylimAEeiIYjUb7q6uRaqo5zQoAT4UI+Ng4QQN+KeC+Z
bJx23DlOGIOitzgB1/LC3ggLcCZi7UyZY5Jwq6AD65u+mnSn9/iAzOM6av9chtz6qhP0TJET3IFU
GFcDdn34B179CG5P0PN8wDL3XglvyKphnMEc513i4g0AZoUl0rKUPOeAnRqhta50+1a0kHcbUnQ3
SgS+ZFPXPfs7a6DSyYH05aA/tyGVWGisyIBwoQ/TJQasw3yAR0rKwJNV1+oKYPc7+9oKnowK1Qws
6wk2hubYr1Yf+qW0DQOpX/q7axzf0awPcRqUiStpVmGSThOTqMEniiAitnu1K5rnt+oHswjelB+D
SvARV7vMOKNNOAfsiILS1rTxfKCtYBQ78QxaEm/GViHvsIfplpym0pNbmmUfm5KPQtDGG/Ab7CBz
ENNw31NuV0EPaQ9YHPrsCtLRrZbHvidjfpP8GXoGHpsaK2ZkVLl3mAEZYgzt8fy21CoXUf2NHxth
cAZajyPfMb4k+IRJiqVwUCdPft2g4FqSd9lQEgwe1PW4s9idO2rVSt5vzcpfnvhDLEKE0rRjFE3w
6qsWU/AsoHIAJIn5n2Nih2mdROS1Lhizf46PBxAVotx2fGXKWL1/PyXl1SCrNssKJlCGPzgt4aEw
SMoQs4ufz9Ht7dI0GTJxpzsViMYJVbSNJotb4ivQ/vHtRIW0ip4wAEp4RiDJkUkgj7H6Pt9QfhrL
gSbeWFJgMbRq2E5eEQOMkLo1qc0b9F+lKQM2kKBdiePFlyMoW/uLaWOHsONTQ7NDke+sadoWALxL
wain/4eYWGZ8GNYNhlRvLp0kyGRoPRCHY9i7goWAThvb3GPhIjPIwJNz2bQy9YV6yweySbzsUNP7
1/YIVobEQKlsutDqSmC6fHUaBiJRQRkM2GmPdqMtART4CAtRw3U65NkfBtu4pLxb2HYkChVEH3bc
2+/xWe14ddwnq1XXI3dCQeXPvAQPR5F69VL/uJCahijojEpinXmJauRdbEByZPecgH9LztgabrQl
jfVi4kZNaezIaY/448kubLQ7D3rMUzvWkZkXDcSVSWU7vGULfsWOC/fkXOYLn4jpgMtJ1tjDwKCI
MCkeN80LMvhYtWq+zOriqBwi1cYWeiyeUbaBIkLKOAIM6uo/oMz8KNqj3SlirVnWPeBpVVayXe7/
/Rl8Oi1ZWG14uhtI4VXRM49QYl22UntgYEesxxVWnVFn8Iu+2QWId6Pp2qEDW/G5jY4rNZ13ZCVY
iKd9iwTDSz0i7LLAz37j/X5fYQmQJArCQQCvpXRrqIAn1mLu+E41NVvxavciqrfvKVfXv0Y+VBzJ
qFYV7DmIYnH5Go9lL/HWSBorYW61MHxFwA6N/fGkltVqnUWho4M8aJqp4AFAeTiDzx4Uv5koriom
ev+8psB6uHCAO9rIaiR+4A5yz3gRP6U7gJRxROgRmG3OpsnnmaTLaR38h2BQXYMPmGe80mQuVnrx
ZkbHoqc1JzQmFRlENUKp73xJA9iNE0jY4hrjV/eHMEVdutdnq0NR1eFJeqmvdwp8V5UVMxpnuM6D
TOE160i5Fbed60jRABKMvRwZiGJShAwfesuFvPMRVNM+VD6x5DRL9Y48dNvW7J88VoHbpqCjzlTu
XwkKDkTKsQdsVYSZHBodmKR/AUZluNUIdcY0vnSopL/rXDcC1bvV79N713e6vI2YU2JcaKoT5cSd
/wV9npGgYBBLgvbcArdfwnQaalLiS/uWIe02FU8wh9ypKw4OqwfoR4QYQ15FfQX0nIN9fh7aNChM
cePhdhFomBySvBlxFC/Lkhb+A0JAIrW93+nIW+YQjCS1Xr6zRzsllOJcOIJDxrqpxNGhZhGKlu+n
M5Rx3DekH/5vNyuHkLjsZvxxVhZrbEE+8ZY1Lnf5yWP6o+CGWf+guZtOreNqAxuM+XzBcoDYlJL+
y/pY1Q5wtsroAmBuqCv+DsufyRs9mbCh6St7Vl8gP7fGjmt1G8LrF4jIoJxz3TBLz3EkZGz/qdmb
kiKGsx5uJ1en9/wuLjl/FDHEJ4O0JGlM0DA1mTPevr3ZjXsBE0NZv0E9sl8B7wjV1wZ61Wokn96o
gUJ2FKe7uJ89Au8rZm+Zh1JKmhl+CtamiDSMyP+eMcmnGf24zkQL4QYvFozejnlZffYgmB2tnC9U
HoFct0cudLEJs2uJE4thsNZR5Ie8kDnZaBusvzzYLNCmqT8btIV3K9aI5lDsFjtX/+YubAZxUwLp
RG2a79tgDeY2LbllFESaGKvjc88DSsKkvBYGDY0SirWk+wqC316iB1+CpYfFrevgQ/CXvbWwrbum
BEZOPz0UI+8amiCfBM8A7iypVCeeyh+UZJAlWdgP55G5mYFCEuKhTrxNm59VVq2PQgTCapRXY0Tn
o1KHtIE1xyZEo2GbnRsYBnX5tNT3nbVDZUaLzFadwyunCY1j+sYVuyhehm7sopSWhcwSWIrQc476
/zQpH3k93cRsuFxEs8mfrOeCRmqDF9D4Iz4pz5SyRfuZuk3x4qB4V9o6VOobKCVZZlk+WMJ3R7J3
vxCIw/CUwu/wxCL7ErnZ4TGOYO6suBMIU5zD7/WvNMcUfLj6KpdizIwhEFGPF2pcsAmxygK8YtLF
f+mJJYqQzSKoxaAQApYOew54pEvYj44aGqOU7RnepXL/ffdmNc4NcFMYSoo5JvFa1EWqx47d98jv
CErEFdU7WwayrwtW4Ww192FKzmxhgH1SksSFYTPI234sBdQEkFyKZGwvNKIBkkngl4reAv4O7Ot1
T8mrPfgdW48jFcjUDzoSIyA89kAdtFiXsvP9LEEuyfGVvvQYMK48RAiaTSx/gj+ZWL2SfIRDD0Qi
apDSfDtzT04C9tVPMlPvJSq4KKT0JxGda2M5tjfl6AXdV9/B29d+JMm+58T0avNtPgH5LBvBmoLt
2A9UhOMCOanskh0yshaLqx+DGgOJ18tl17NXto6oJemdv3XKFMK5t8P1EF3N8/qsFKPLa/2epc4r
PxTWmqzPKzVe65ra36gjFWU+aNIhTkDgcamd2QMqt0Upxu320bLshLuC6sDGVJ7TejqblPz1NN/X
/zs8+pO2dhA4gXDj5j58edY7lVXpCtIl40PrVGsR1Zl5LiJdQcVvxDDne53cKFZQKhxFvTZOuwcH
Rg7vWgpF8y8p+eSpzv+pywEh2oG9b7YSodC34Hqv1YShP78xMTshA1mk5XhrjF6HcvhdcW8xhAm3
8PisWKCw9kG6ainmOpnCbqGwHq6M02252pHE9E8xm38JNas4My2hY9D/zIxIR3X+6d80N8cZqBqe
FlOz8uLoaKQyxZ0nWzDRUUpZwVidQdUw+QTnd9HfWk52Tqr8M/VYhUSFRaht8H4QUg/4nDS0t8J0
+0s/vTQqDyB+uGh0FIGUJNX8af88wDbzgwId4r25zLyw3brUtbTtzZfHS7tDgzhZqh6oRBpGXoU3
UISlrfJebwY8MgmSZg3/GGpElJ1E3WdJGSkzmVZM7vuxUKe05bOGTZ5y9hZch+hhRsY+QqOQ0YJp
mJLpO/NbS8ykqyuRNuWrtjeofInNXanduUF05ZfOKsF7KS9GZ1Y4RexYlHt1e8fd2t2wYvOz60P3
m9SRv1kCQ4iKryAwiNYN0PgB3XdTVBxgxmkxBXMk1m2bBohKTR5DsVFw5lgcpgE1TKQl5VVAgGSA
2n+SumskWk9wQGLfSWvdjC3ZSjXmCvFCOcbRpr/7m2QztAAQH12daTYwBM1LZZMaGtZW8I+iH88A
ZyatRihjhYi+mv8rz7lgK/vCuBYz3XMs/LDISnrc3unrpsPzqSe76kTzA2OTLOPyHaJ+bSCm9ZfC
2Ym4kA+O6hseEImhPlUrTXSL8NKP3GD5m4eAWUS+T1LDielf/M1Te4LFf4bsmsmXC5GtR1QiIuuy
sLPvhH6KnEGCtOja8buailvHUft2ApIBnBv8jyjtPKM9Crz9zXjDEeaOTnCw1Ezk2o4NrZfkwq1/
JVlfEiSzLKznD6pJSSjrBXEX+fo4BLwfjl1Y4WQAoViVInHLGqoz6Ctfzp8yt9lOhGRovGX+IeWm
MAU8IgmC0DlMcGAl5JAOz0mw9V587pzyh7HRJnazxiT1eCVt6c/6udd8nLmJ+ZCpJu8zIAc/z+zS
0AyWWhDcUCiui69IGdMCzgI+IHe6wIzbpS6zoG7PlWAzzwyjYJ5lm2EF6U7JIFPzXe9GEqt90+oU
b1rNVlGUSN9gwXCtYyQUSjP89WuRDEql+HsWN/exDl2UdFKZgR+TcrSnskxFe/EDD6y8ycLsMuEz
a98Gr+DfKMUivPyi4VdP6s76Ds2Hsto669VinpryXZn4A9ywz7VPzMvT+3QAEYEjgKSrx+DtRTG/
G/90/jJM+kqxQAV/tbXcF+bR2dLFt29E4TMJ5tlPZk9XSpMz39stU14gSoVtI0m8RSAVE7s9N576
nJK5hxWJPtfJK0YRT6Si4LWRBlTdOWr5+mPgqrcgSgc9Xk08sa8kP0U5BG21NF7HGXQLBoBlZeXM
oCrXJBDb/w5sbXevho5089eU1RKm/OkrtPSlaRIVQa7pvtveMbxy42v1DSfpROZHNIlM8CKD03kt
bLYrhjUwAtM9cb3I4iJTQC7P4Go7gM0XOIJzzKaNc9jyfqHvBIVfm6QbT5w8Y57w6KvK//A0HoIF
pyLdlHq8sd14W2Hmao6CXisQaN9GKnViu2/bV/SRSrmiLFeqncxtPzYQURcsg2oBlTRqOpaPa115
uxsa5+6Djoz9C0MSciHcCzCAYQpvSiQq6X0Yiw8I5R8OIG46Bq57ETS+/diVo0KVI/H3Twceonik
4dU8xMFaMcqPwLtXL+UKXYqgiwGy1cO7a+u1CVoO4s4rzpu/+yn2ZWMGNPfJfrQJ3h7Spzub1Shh
oiepALiFfWZffqf/Jb6H3bgboF5Du48BfdBqIkNgSCaxxj7ae8AZ2s6Uks+49KIB29hWLOqGgvqf
/g1S+ZdnFLLqKBP7i5zX+5Fl0vFOyg87lnC9aJ7/Bzivi9GqCIJdiLmrk3lyL7aYpKG+Vr5UUqkN
zi6SgwIuatnuA8oEHXPwoAcMzeWPbos9tUY/xmxUe8b/HYBWZqjhc7kBq+On9fK3Sot8qJIFXsAj
Di6LCN5exi2COkG0sfr6JiQYYVdLhjBsr6z6LFSxCGyiLVRkNxLfhWaeG3hJB82TV6gDqrv+cJNq
s1IuTh7WSuIfMUejV9KMVZYi2cLgAaNYqTNWamKIaKpC6MqRlmDom1//XHMRMlMDaEFgkGYRQMzj
ccqKgrj1i7hG+lJzwCnXxpQryleajcKVp4N4QdXWRJODwMlud5fW727tBFBRYtql55i0xiUq03Jf
Sdr4JufaETpKlIIPP+YtSKS+AtPFGcPmXUZ9owtdkjuJumr6MLXnMYkZGT3mdLxmxD+kRpByCC1a
7uMSgvULGOHvUNLPPIrH1tPjBzn9XRB5t3ffWEqPaB/1YSwGyQXmPVMj+sw05b4PLCnQcBmCwFW9
N+00e7HqPt841R+ICX/hxC35BMyOUajT6k8pyHiGvYdamVHq1gGS95aEEYk6RUY3MF5OTyhyt4i9
spRWDqQy5szYilqGS/XBJV7n2YO8znn/k+8cKmJGLcJOKldAOnUZDU9KTq51e3nI8dPm0XPIvX3Q
7bGklsnJQjI8vQGe8j/rWP6DE6nObHhUpFfA/u+hXjQGi1/ZzPUAn1lZZQUHkPWstvx32bEWZ/a/
URdf6HErRS2tih49/vCp7PZAZM9+XwolcGjQWgPqzQrBHoPbHWVpzSvHYp9dVty7igZC+Wj4uuwu
JVfXYuo7U6Tmrcgm5gjCAXAEtwSJ1qOmcui8Ccjy+u3jjU4sQKIvYP/cypTv55YkQlfgMyj06j67
+84I6Kix4hxTjNvaJ+CmutBBTAbCtyUX97DQM/QelmA6/LPvM3diGv4LG/9EKJNpJO2XfWFapoyH
qm2JgFvMnUVeWR8lWYl/5Bgeja9nIZ+pVYdr7HKQzCfRLFx9K86ckGXzeGseQ9fzJ0xWrjhOcAZM
zIV4/OZv58v5YRHWvbO4PlFHKqAA58ldTJ1oTX0P2fiXAnUizeihcDXvn2O2XFMM1Rg656PWRNLe
esniz4yyqwK94GQ5HDQHP69lB0zhcPDmqxGJ10KPG+FweYmBgbgWB1qipZeUr7gLxbCqk46LPJ31
fIcX2sARpPwXI/rV26Q2ys3uALJ8R4rW3OXW1IQK7rMlFhUt/G39sBRDAQnzV+IICPQrx15Wyp77
dpR+GvESolDvbGCM4TtdIAN5sseMx8TpuTg7oHmTk/hKpEfwqklPqTqvC2S+ue9Iu8yEoq/Bp7tF
8tTmeuYsoXkpt7lSUQuPV3nGoUe3H0PFT8QLq2a8R4ENtLVFdX1KjBIm0S9Zq0ZjGAS3asObYcD1
YUlIzLv6cYcCtS5paMHsCIapvzSlWMveIE3oALVxNEdLE2GcnWDHhrRid29F8WJRSfXqLiX/sAZw
yNoDkzXshAKQuy1NR39Jng6US88Hr+63joXwqZ5uc2okMrQtDpVLFLZk2+RFZnLGMl6TaCgPwqM5
+DAri1UPbLY8gxgtERm3VGQ3Zv68Ib5IZ+8PjTEVuJnPc3F9OSZdj0WdVEDi41Pj+DXhZ/kve8tT
FchJHS+WBd6PYZdvPWNJyad6aW/U4/cEz3vPLQyUV4OTNJhcF8f2BlGlLWrxJaYBj/TIXV9YPSeZ
KTR3BZlQ3BsuBJyIAloLZeitTO3bDpP0AMRdAFqNNvNAKYR1g3/tP30VtdSA6+OYZ+QNV/7ATf/T
N4xVcjWRaBfZoB8tQ5sCdfAjwKaLIcsSW0Zh0jSBcmGVVqTbCyccplY53E/gIG2MMd0OedNTonJJ
a5ptJTy+8yGlZn3qGf3YKcWtVfaGn0pgvLUhsjNPGyrg9xScODshTRDcCbAWWlT1oY13YDZToYPm
NN3U97WL6gUzr+M1thCpHU144rJubS3kbRWykjDT235rfJFxw2tM3ehjLl/XhIJgv5tI7dqFsLMb
xAB6xZ2/kiXKtHNm5o9B66SZ5fZrWhtXHdPwWHW85Ot9lmkTI4LkjtEEgJUMBhFfRfwawzWAZfWQ
XQN09tf2I9ReahZpoJUI9I7lLKUX3vLJIr+FNmRUMsOyrHpP52T+1nVR/CEdAFQuhICa2kFSn6cI
GzhjBO7imtcMS2O3nGq57/LYNzLcDKt67to6cw3f+aDL5ZLHRlPRnQNvv1ol24zkhL1vSJBV+jnW
xdrlpwIjnvh/s7EqiiHNlEvulXUBuHcBlGaPwD/JT/NN6NVdiQwayl7hooEx7W9zRFee7PXxDGnG
FXdzEPtdTLuzHgHOM3tOO3t4ZNuFMMaKMi7FmHRg/aYxs1eu2inVhykzWKFIMopEQ9T37tOR6zcB
omJHkobXhhYBXqpCfjznW3h/EzMJpqr5CxVf/bMZeHMgh8zkvOdHkjgIkMTMyFfb79V43aguwqzV
ZGPnZ2nwAZT/FlKJ0gZaML7VKAHlV2ubUIIWM+E7aIqBB8KJxz9DC2r0xwgBKhhlDTTecTSs0yU4
CZ007cXlrllJGRKMTHWXtjEGLVCOEc/HliwKiTKtIeSRbRZy5UU0furihvHlV0rzqOmBi9T1+WcY
ldCWm1JfmAe0nsBc4/M5igQG79GNWmzfN2RnTaHdBPVlcynh5j/bdMQCQ3wzm5hySsRfANT4KsE3
OWIPsCPNHXShk+2k6DByarQ6qO/dQbfBrK+lcsrseaxHqKnd8YygMKykDhqPHXSDeji2k27SQE4v
/+S/eBlRpzrj+X3tmNbVJNowVVGjmZ8Wy7+dF+/XtffN/JIPchWu/2r3ZZi9HhBJJaqWl8SS6d2t
PMsWn/FzXuKrc/QHPwkl1Ce+ko27HfG1BsNd8UY9VF3h4ag2rWFRMJbQLWjF3D1Cft3Cm3nN4tkC
Ia9XsrcB+S1RxET995RXXtogmHDAOTwMKu0AB/HaO8yxAHTC1URUi8HHkLotL45vjMv3j/yzJwdR
F7XyvyAdg8JiwVboCQNynmGhkdQL9FIP3xYvL6FsZC+SyyniM/LWE4O/TcjY9LNjVOZ7rr5Rk/JR
Yj3V7bQeOpfQ/dm4i66PTr4FJgWXLOH8L+GiNm2LgfTZXl3+5VIOotRueEuD1CbiklS0IIfcBbKg
n/PAN7JEvfNtdCHPrr85PTEj4hmDAh2DbaDUkxqkHcUJ5g30d9Fm9Tv56PWptyejllorp1Ijnyqp
kkExeACAbOCUwSpJ4DGZPLKoBPL64yGPVqu8HeZUrC3VRH3CZ7qm5PLInxscXqVNcugtdIbjdcTz
1XNAU9e+137n7Lk7wSI2SAWj4Ms5KVHrMWEWV0psXG/Dp6tGOA2Zi6/GiGrP/BfQ1xzUBqUxMDgt
+HvdZorIsSGJ+/CW6bzLgMLB0oBengxpF/InoHUQ6SgMQLoLeuJwmvwUePZUomFmkVVHHP9NQgCk
F5dh/imVgg3QSsDOaUZmkOneypQjD3O5L/JvITfcP6lUDnjR/sBzv8fACCWZAxrz8KsREGz4kFg1
dc4mSOgIES6vB5h7x1hfastGPPMFWhD/AX8DIJ3pc19Zf9qPv7ybEYWyrvOV4kb9WqLyRqftMW0F
L+g9Oq9SiPAGeS3fZ0iu4BnyUbpg0vcwr9zsafdS5HLhExh9Uj7k/WWjDHrU6gmGPBjgIP9vJ15H
C9nUiLbmcFhAZTV6pxVMNzq9jrPBW3XVmslVf9exj7XSbMuLnfSpOkE9zgGCXoLh52Uy4BfQIxAt
KhksDDPSUo0qsKEaYK1BEfU40IkT2vp43Usl6kZdgUFTOMwX4o1pTAKztyxHfJlQPeSl9Y1zHgYm
UgnedG7ew1nVam4EeUFtUUNTmUPeaqvZodzg6vDvPMwZEd5ynAKwxnU6YkNIaGNHwq78WgFwSSkM
QhZ2BmBZXQI/QL5QO6kzJF3STWFDboAy1RMoEqRBlcg0yAE3bMXo/dmkTAH8f1IgWNaLn4W54aeh
bCvLIvCBPXeOijxXdNFneuhnu1oSw+PO2L0doJChph8+Lf3AqfWakp5NDdmL3tV+j8A+daXsaq3a
R7SRdyKFXQdlV4ANfktAemj/MJV39AxEzrZo5OHXTaYakF9XDgQLaVurnlU0xwYTXskqvR9FppZF
K6XeyJOAPavDWGUp3xmqBjI7V5y3TF+smjbqdCDVh+FBuW5rMwX+XJK2fl8+geofKe+fYTSi5wZT
ITXWYo6ZfkuKJ2i1uql+1TzK2OsBci3gLjo+fdoa2YiFkVhfJJeFiRtXBScz6MhHzsrJGrrnMhk8
+VLfb7FoDu/OuMgMG14/UHgss9/kNV3C/kG/MGj9h8k0bCvLuHqeu7ke9g/vSVbY6FgJT1M+mbCl
NUhqVuirraNy4zxrGL9488bmOePx1CSUVBXiTHDFUwKsnMvSfAxqUfWsRnVSRH7ncxdknvXUqI20
cp+6O0of+/bxpLNIRVtmGVQenJlpq3NH+uO8OISMjgHjzReUbLeaJnZXwzktcGhSYXOZQM5Nlki0
1UTGYEKG3zC1lsOL6hcevzMK7AJ7PjzX5sbFLekwUgePo/oS1xt5Mih81Yl2wnoYIu3kSaK5IIYC
Ts2Swi3uaL4MA9nTNCIPNlvcV8jdfHiIH6KXqew/q+6sTItVTBYzf+X65nEVcEqu1DY+TBdHoMRr
t43odVDLS4MXktOZxKsxP3OyexRu9TVTUxgqn/nePP6TzGkUQ1o8+qEcBWQifq3Lzuq5ufxsNo5D
xlokr9i/X/+VZ9+JE+Vkf/YlvPwfqSumMI5/r6YOxBz7HiqSQ0htcEbNPXI8gWTRO/TM7C+B4KlV
obHKy0oAxwYjMSv3vnqvxtSfvzDqucyPT88xUmEIEmoxktIwWpxkX7c5qY3Ahr4tgNNwO9egByNM
GDfe3Fb1ZJEE1uNJglSU977WRPnLVJhVcyq+XO3F/bYK6dDTPk5ir/mncjZxO1oXHVYH1bxOk0OK
AEnRd7E2wluLkzNljXatZVxLHEddyonVy4+DdThn8dWYznrM4U/rcFjaOchTgxlLE8Xy5opBQEmS
z46jwHPTm/oqbE/qUavolCjUPGx8dh0W4cyydwfrjBfXGIr7OoB0kslIfKl/pUL0SKkdv/rFk0bp
7L4hkzyCYC1OpskvKJKQcDElRlrM+fKte87Psr+AHypHodTTpfpN2nfoCytB0o13ewbFSimlWMXV
BdRuS8Ful1QplQytQlvQ4dAVEqG8/Fv2Bo2dQr6QdvzqEfYvuv3Kd9npsIwSe9Cqqhj/2gHPlfaW
MmEVmbx+bRfMPzl00zuzESj49H+o6RHBKTA8y3/fya2brmnSxtjH66tv/CrLT9vO4K1zVhCYKi6w
5JGqL6mEQPzqT2Ae0rMrCZFOAeu9T1hPRQSVl2QGrpQEw5JZC7pk8jka7ujvGHXC7KsTiL0/eV4n
TzlndFC56+Wigk4iMW8eF3q64HUIocf2VRY9f7H8NstUqMmsF/51vAtcYxx0xLw2GUDrNJdSLixG
o8fXGk+ZNoBbXjaZvZ0Sf1lVZL5/JPONcIZxHz0TRog/dUIsx/51ISea97qPotuSdKi+P/hbe4/A
6jxY82FHCaMkBJaRpLILWNneaQx80ENg6HPHuVz2LpLYWgCJB5EPNpt7iSS2X6vLN7WnMrHFJ0nR
oLuBOYiM6unBcojKB8hS86mMSnovebysJgZhxvXjSCiEv9AXubPkR9YK3H2KWeF+8Zvf0DYa9p27
RaN48I+hW+P23SvzrqCNqIRNHnPc5IqlEMKymj01qgn8xprVB/QyZVFflvguC3JfOsFdCQVhFPy7
2R5vdBwyspWLTn5vR83ZexpVr6nj8fW+9o9MleOcUUfRL1hhPeV5rcM/syERKV96Yd6q+4opVBu8
DFNAYyUc/Wo0J69p43RPi9BnSQCEs97JCOC1s2Qp9jLLePAncohathufJBzZuEbzvAcCpVQ7kfsF
8qDPCsYwtcjWbh9lbAzggxV6WcELzYxxsIosETrlNeFB7xB/FgqqrxBi64vxSNjYc63UV/uPB/T5
wvj+mV8a6RjmOKld/MkRbo9iXt/t/piJ6w3qnYxG4PoL+kA/ArW0MTiqNcqN4vkuE1MuQpwNso7s
dxn5kJ/W/y0t+q8DU1PdLhd9PmUUPJdqel9T1OYy+5AzADgs9kTSK8bqPXu/22+ug5RhC8cYJ3fR
h2AMdMMfJSuPwAO+LfB74xQllrrLFKx/++xz2O7qbtjkfXmtIM+HH3iQJE1k3oKut7Axdg5nIc/z
JvUinFai0O6Of/rkFjS/dXPb+hYdKhHVWK6VebRDFEgmpVG0sFd9ktidvBWdkHL0eD8sqo/Z2xFa
vvTLVW0V9RwbCZ1ELicFxAAerhNyPQcKEVE4Jpf3A1izYqD0OT+jyvdEIXBlSDqgknPw1NzPatMa
I5hnBPdBuh3j8WafaqpYyBFMCN/TleGQC0vcbD0hkkUE4x/rod4MIl10rXbSGax3N5TrgYm9YiuS
XIMzLQb2TtDA+leOg8KARkZ0eBVubc7rvl35Qs+xp1rjma14eIRs60cZ4SchWu1G/BDpO7h9r8Ji
f4LzvTBqQirqjejq4h73fyioiSuBYVcYLx5SjTfEz1Rkd1Er1IVHFz+B74AuDimmye4qOK6Wgr9g
W73f6ZTytuc3iviFpLos944LVbFugXR5SUL22t9F4zFrl46c84NYULXL9jh8EYliPUKPfa4PKE92
uoz5glSeLnB7Db1U3FG9BDkHC6AwTx4VFvjm3FP9D+SBNaEvhN1D7W/Q0Kjo7EwzNDy7ENLgdneQ
MrkmF8SjfxH0cSsr2PVAKkQTGGQg5p47qglIWH6bWOeOM9Ww/cin/spE6aLWkM3k2zR7pOjpzbmF
wbFIqu4jxq6zjaos7UpPLlV56KbjmgFqQIWi38W27mLFJ8xXjd8Cvi6CwLbAWWmTRtgQ6DIYK64+
TTB74Xne3B8p+hgRVTgZSwtw51+WmTJFHCsHZwhsaXjZHEbAk3nE10DntuOCStXkj4bBdnQJtyPS
/EH/3tc/5HddVQxq6mP74A+J3KWdr5yTAPX2VRgxQeHTTWzBOKvtUe8POmzJ7ThmwKaBY9Gi4xAg
cAV42Gq7Hy3HKygs8kgazc7UtLbvtYZQIdxAgpedjdMmc7BqoJbq6/ya5L39sHdMXfuBohO6mTFX
jFDhmjV1/9buQT8Tlacmkwpeqags4PJFahMY5YWgestRgkT6oVFn70Dd5STL3CcjEd5gWMHUt7MO
tDknHCrdlSiXewDAHFyCKDYUliduG0wS4p6QofNDk6dquBswn37E3VMorQNOQ8rr0JGt3PgRtTeT
1sTJktAyWiO5KPnZtwfhFMxZXPwyXYs+1ZJuLHh1d5I5kcQHXaC13siISMljIlSjiy6P+h8hzxyB
2SbxpaPZNfhu6KH6Ux87e7ls7ANOyTo39B3DPuh6EKDoSqmTnYGElc3GR/RQnhPYQiiBSxk6HExo
xOztOR/XqWOow+Km1d+xroHbIp8tlQzkaOx86sdZ0KlxQcRL48L2jz9n07omqNd4i2PCdFiCvClz
3bMxrX06qF4h6uOif40muN/wF1sLhUbiY+Hc8W34Vu4ZKxRyM7qgQ02333w5gcZ+LCWtPwtIVBhh
E3zWB7qVUydGVX8a2gZ0YBgyLa6vlwT87BBIQkEGdzngNur9YCNXmq0eW6iTbesTu2F2i4B4zUJT
ZXatFkCl5dfKkQValYqvrVys1vZ8kSWJyL3ufgDre/IHjLmAgVRQgSiLC6XvLKqutEtNNnRbjxUI
FJQQELxWAWvXeb+MkO7RLfMyqPwMtQ9QdZZG3cV/I5hEn1251dA3lpUoarOp+MfduoSGlp04hgUe
D1dGR2BeIitv1yPk6pKFW+BN/N0WhiN5QEby/ZhHQ/eUFBjrlqzalznHl5XCLagAuKkIBEPpuJqw
IE5zzfINllvG42Bvx7EoIvAfqbGA07gj/A2O3oqDk0k6LwCtbysASr6lgihxQ8wSUCNFCOQScy/n
3RprEGHBumduiBQJmDxCuUMg0OWfYtCegFxH4XNFGX8D1VDek7sicpnwfA2qZUniTp+UtwYWmr86
2AlnSnZ/9Ct/6rrWiN0fomAZzn1YYyyMekPTjoFbyXDmdnhJwYMEJj0d2OwbRKPkY/O9OnraJS74
3LSegER3ciz0adbyiAi1T07mrda+WJXJV9hUVn69CjZdgAidFUM9njOg4A2vPgAxMOwCYHLDQkvj
JooABRDZciY+vgI9kjkzxSToqo9QJCkw0B5R2AsdNW+fg+S0jDh96auMTqg7NPmZ9yWmvHJbXLzD
hj8h+SLTwEwOsIeBAPvfrMVgLxazgSs/NaTfulrBMCEFQSGmnZBzqHpDUpXLfy7oCacZlj2twqxO
4qI0DE3DaEx3Zdllz0UHbFNUdRBnmp3MXDHK2ZlDoPQK3R5a3Ii2qFdhMBehO8yVjH8uxOZT6j3i
szoz3vm15sgAI+6UwshFAaZpaZXWX1uJ8v6IjPtZIpKk8Rkmq8LaSVmbWkxq8jxz6tLKKFxI4+rX
NZRjPR7h2H3KZ2dRYz/s8ey/n/6tEPJAIb0awnyOL3btTztRN2a0vtzmR37DMcm1iW/38faZaVJ3
CS34Cx0FDa/NbWJSNManKR+XSdep+964KdPdsrRH5kERn0WfXWbWzgBEjgmx1UPskcIWWHVXVLks
yS5npVGuq0wBIXv/DIsRZAVEeybtz8l5pb9At3ggXCyCFPI8u9AQpCxiUbqnqIVXYngTRYDEkK0f
IRJgseufdPbeX/DAx45v1XhaiObwoCYHO38Im7lBXIHewTOt339vTZVOqhhy2E3mUk8dPNt38QFi
QhsqGE0HCvzTpN6b1Oko9J84jUMFy79/Rlx6ZskrDMk0nQZUXGnxAqtwWKfJelMwCWFX55/ZCZ4t
fYqbkG8dEUxVUWphvpyYvKz7PQvipVBtIme8ZWg08cl1qXEAlZ0PAfhaL/cbKfMdjuvrvpW8n1Qf
3Wwmx+XO/4K75JXh1czcXrxsoFkYPoP59S+aHkDGN3p7JYYZPhNiuz3HFtM7SWFzMaVxlgCSdhU1
vGn5KfjS5UOtIn4wCXwaH6pbDGd+5Crqldy96IoZ6Q50IJEemeuVVCJYo6ifz5FvPIUTWCBKgBN4
k361/2EIfUSAMU+lzJauqrbQcqXCMMgy2nwsOh5xsHzfgEJxO8D4SEdzjnFBVkU41jUo1koAMt6U
FpQxzFegtG7v1h/7BCx79jrAsoHIQOPhaqeB+ggufvXA7N5SvZMpZ2lGjamqmUzAPIRoTRxuBWkb
cNuN9NDG1hCLt+m5wv0jA0v+XFX5LrkbNo5xuoajjX+ZI9qtOWRW+J6AQBQYq/eezq7DEuWED1uX
n3ZLrTfKP5sS/AT0gFXyjnRgxTM//PeHS78j0mvsysTjh0kyVjgPyqs2ExmdvRuPMnPhQSsSZRAj
bAWeqDHPseAn4kP0K30jLvfrZaVxAkiILJy/4NsLo4fkWJbSPRguTIq5gRs5q7sePGy9R+rojLbJ
prE6LK9M9C++m3X6ChM6H5ak/f6G5FY2kCZ3qOHLC9Cw2dbETb1vVGFjMXTU6dsvQ7jlz6w3eCuJ
+HTn2vIdNhzTDS3T0NfjRucRqnGmBW5YZ5QBiz84stj7LC6kDKz0n8nQy0ocxHr14Q5XYXa876Oi
IXiQFp7UMaRTdnC9FGxoHCazAfMmRVQ8qFYaJc3S5/KHg5w1JXvuuJT4UO76HHE+8YF9kq0WpPUF
SbfjcRB8tJDswllwpnggmdTatvqFPGSwZbBwxPKIC9Zb6joPBtd/ozl8yzotbNMjxSCgynT3gVKr
AsfpojBV/fmdl8GxjHqq91XtUEjHSVSEChjjymNS8CKQxtghmaXxSopJHBGtTsRk1CTn1G2s9lZ/
+7dGkS09tP4fgxia5GcTHlFx1hJSOGd6j0GVAogiWUwS13wQLe8KwRnrobdFsJN9DWSBYcnVMip8
0Y8GHu13sfiZsKMNRL2yOa1XMKr4J4GohJzCUgWsTSpEzN45cVH/nwahUp3kyqDfSUQWtsNCa4vU
E4fAUGwm2+pA2uaGzO5YtodpG46fpKHXi8WA63CiUhMTA6ZVMSlrSKCFo1KAGZTiYBiwVAQ4x6kp
I0/rKZpPuXpcPOr4Pd23pTck18AILJxuW8U1x25G17vyf/SgQLO8CdQY2DoEY5fYGVLikPHas52H
eg6jWiy+WAats1POYgpGf0lbVei2lqgWqekcEGpKEglVb/+5WEU4f/trFUERyp0UcUxsRw/kHN3A
GOE70GWg01nPhW3diLfGnA1YAmPrgqPROg4IcCR85eQKVxttIe54xBxuBI27MLM40k2C2ohLE5yb
co2DCghn1SMFS3EafNs8eOivoAA4wx96T+GjGOyX4mIjk7YUnVDHk4guWnpPOuOqm1fD8Wo/dcXd
MO1yPHaziGaIjH73Rev1FdTkct93yOYmxSew4BmJnMuvOvmoO3XHK+mPxFF5me6ubrXwetvm5ZyV
s51xlGNo8rz+CKiX18Kackm7XOwmwRJKMAAq2ga0kfaYrwFwaAKYiM4bA65LTWTPANsUkmdE0LFx
Ztd2DIweDUfq5a/QNrmROgFP4QqtDZB31oIeT8N4Y4PSNIgU1F37f7hOjozXM8QA5poZO+O1/r1+
yl6a9CJBuYEQ3qGGtqLQfQqgHfeMPoR/G0xqRD1DXQZ7jArpH4pNHcZlT82qLpvUbAp3TOTLazvb
mScA5v2qjOZNA6yrRj4R91lXvldQ5kr1o0sZd0VJN80TJoyLm/rjQK9sY5LEPBgdTHhCD8cqBxCZ
nv2jNCFe/cnatNtlf918amYrXw/IxcertxmpfbdyPsOUsLbJt7Lly3PK7S/0wlqlawbh+BEAbwPf
i9FfIyzJfqR/vw5zJHyibDKO6OVMnNLFAk8C1QmHATbK3l+eeEHRCeXXWSBBQnMZRkMgC9+wtXZu
T/VyKnBcLpunM5ME0Ie6IziEBUEl46U1Bv+IkYALtXs8knzjk1YtUTHsYeqj8FHzTHaF/1Hl80Dz
hbdTPqa+8gIERf/o6dmpgR4zLoSOMxM57QE57E5lVAfSNe7W2GKWQQRBwim9ZPXAUUU3By3UGDbT
11OBPnAEJ5ENUObbJjBtNE8MdNrXrQS9hIj4pFVyPtoue8sGOzEzOokOWk7qaNPukTI9pyTDKxAL
vNIUUTrLQ/6TNft/Th+rPNq6Z/SZeQHPZA50OXtUp0T+CVgPETrI6X4VSXd1+M67AEY6gTAwZhiE
JpZ9jtKx1jl2Ij+TJIMZ5Lpzp1L1JO7BgDScI0d9pnJgXdaDnnp0HtUZtj53SiqfK7+1y5Gq0o7w
rdeSrBKX7a/pdbDXDY0YbFBoDNgCZ5lNqwSjgqrr/khQCygITviMzA03KVT5kXvEzIRqWCKEM9E+
rzu5Rd4Y+gLikWbOgkR5hM06oPcq6I2CclJQ7kOxJHIzW5VemVv4VEmBvaCjban1+bporrOfu2UP
LDkzcdyRi7H7VtuRhNHKAEJf+ry4vYLKBteesO9gXOMP98el8aFJjuXD+ezjs5frIwVg5vbJZRXt
kEwtS45w0cQlf1J4RQ0uRVFIWnLYG7olSrt6CUNYnGql9z5P6JwiFvH7d7S/KUEi+QJBm13UOPsA
sbpQvtr/i2YjBkE99kK27lhvfedsOQRVOCI9k4jTiQLnqq/grcL6uD/o3iLqHfbCaLxdytGklbam
nfuMCNnAApIZXDc1lO2acR8Fep+cBlytMDR6o+blStUwbLaNBrzZ15o99GZs2pP6p+nsxXYKld5r
5sTt6ug6ruMCjKPzDzRD9Jpe9PS4UY4tkaCL+pghldrGfTgArFM2UuLWmE2/2ti85Nkhe0GyFbbY
5W/OFkczZeYEMUztWSalmml3kEcfzccpNG/LP4wXOfgARQwIU291/PVECEsbVj4Gag7HDSi1oY0n
DvqSTZNt114zrgp8MCDVugf6PjEMwlYthHHx3KxnPOA85LPZczRmY0jWE+JMfm75yxrGq6SJCd98
s2aY5rmjXq69x4iBf2bPx14bnGpYY4zAowG1CouKWIQs+C5AS6rD3aEpBGksHNsm3oMiiXMwUihk
lH2pedm1q5jD+fL79T+qfrvo5Fmr9sx6QlWSNu5VFn+UmqjCdRvh1+7kUxN/1pw8hr1o1mtlhPiJ
suMN8fOsqGx/0wgEomlE2J+vUokrce67bHWrOX1RIDyC7baBmQRj6lHFw3bO93ArYlZqDdKxYgW/
EgieTuyTFOuXDpbOR514OH2Y8DcT6RMhrn/X6naZeFYiBH4JWDRFp3HHH06utYQKSELMHRmrUKbo
P5VkaIZ2FRE0sbk2+KiIh/ITyr/2cYYFRhDtNJ8u7vtVau7xQ+M35zNHWH3zcoNyjtmaZLdgQFZv
/sKmtPK9kLNz4vfP92S0EuKue8CblvKQytg6eUrc6HmvISsxAlavHjvQLf08q1LWEDTyt1DrVKbO
KVQbZa9x764R7nkRJ+fJgI38HkJ4JRdH4m5e3SduutW0OLwI9dAxqBIRHa/El3Baak7TK2ymAkXU
h5zJ3jAX9Pza3vKLQnvxKWUeiOGzl6tpJtTgh6w/VpDLMl74bRsMzTIJnGYhstsI7B5cL8BrVaAj
OeA0aClGBQM7Qrbew/E7xy8hIBkI8rA5ULdALezIuz0PCOTv6GE1zLcB05VYDb02ePeyyrFw7Pgp
ifAyogyrSxK9SO3/PFuOzPmXYgjX9ZuLoPVvTOGiGLZzuZTjHYl6RDQbHJE9Kd2uKrGyPuICOjdy
mX8ceZGK7jPjAiiALjnf0mdr0AnSCuTKNSsPKaHv38WBSw4BQTGVs3Beq53BoCAfgVqUTPBf6v8W
QvGZYP2JuXYfvTUizujNoqHt2lFJ40jv6Y95WpyNWnLz3W927i/LNk/DEPowbmGqdb3r1Gw89s3i
u0Gp5oIgRrNMDp4ffclGNH4uLhUJKV+uV+n1fCwE7OA/EYb4jEOmAccTvxHC9cfSOlbbCVrXWUcm
+NJqM5q3dYyLQ5u4J9JOXKWTDf8ZNTc4gCyzkKbZhkfEPcxmoR+vsnhbjEWZvAcTKTt6SG+UzM13
RHeF3DmsV+ao3tJ5WJww+oBieYt36BCjxP2w9FDbA++KXmKn6Jfm3HOT79oXZjwIno9yD74gS83v
kS6FgKp+Ydt1WjEKV0CVc6SjAz1ew5fc2gtCDAwPjhxsaAse8EzibtHWnh01psoKAkFfrOI8QTWe
UaWFZJwsD8tD766M+kOH727KvP44+rAR7VdCHfZ65Tut4Sb2TsiuD9MT7rt97by2HOTXwlsG677d
ZVuodW8nFseu4kh5f2CVXgLbKyZPU2YWiS5Mz6MIACfmffCM+h+dPp3rB4JaeCu8/WUCvxgRmIlN
1L5bMGBtk/unzOcuAtxhnJN2Wn8oiIkeaC/1r16tGa/W9S0r44UpDEG2aNEN/GBU0LsQUD35BXVL
Zc5+THg/o0fIDG3JdZyuwOshd2B6OB1RwTCmQewuvWOrMNs+oi/QzG6oqJDtMONb65cm81nFNfYV
gZjIeEeSA7eRg+Swb1Bi+YdfsYP9/CnT5cFb/3GhtyVRXfnKIP8Hf23z/AHSONA9VQ+pe6E+zVt0
S3o3NALX70SwCOstc8QeVMbMja2w0CluPhSHo5ORNFUZ76bIx4okeuX6/VjnGUMX2cU9dSQtN+/5
kWarYyiOmuR5Z78PpjCr3vUz6P+w19ygfEZO1/Kgevfeosrdh6CsdIcUMD5dbXn3gCY801R4w2Dp
5NvW+VO8RoUJXRRoXnwutiK4hfMI1Zbo0n/xBGgrOYhuPKe9uA5e39cR8UhGGD3Q2//8Sby/5HtF
nawJtcd9BOxPUxTv50TMmCc1c7h8kYllboFPOE37JZO2ofDp1ff2sLFXgNaJXJ4wqiANzl8DLMxT
9CYmL+wpo8ozu0LfhU4tEIKs+4qHaJ+4XS+/wHCIZpz98Z0BQU2yrDmfx2pypkMZKNt9u1ZMf/Ct
3CxwkPODuq8RnimBL40CiwUSyQcxbgM0bMaQ4zHELFmshOvlSDuEMOHVtYAtsv1ceR5EqyhLP1pI
jNrjznOHvNAW5xsEPn0SgTbuaLb0dbsASmeLBmDBRbBGk2gB/2mk1I2+Rh7/wnDqGfSc0r/zyZRr
6dZBTwwmmUdILq5cmd9LHkBbqPqV/a9qDh2389p44EtvkSrHQRoKlTuzxPS4VtFq5tzpaQnXd/Eg
0A8yysWtmDa4AGr42cKwdACW3szMnH9OKLA9Zbdb4huytxVoW102ZNfJXToCsSQx1CJUGNvlKzEe
llY+wmFrpWiAKTNuSJdAt31GL3YSJgEj9O7WjdblDtXyYRjnKT8xsmYglVVz3WVXcG+eeibY9BYh
ogyECDRrvDSkOdbqjGLrOOAkf3Rr/YbGeYl9q7yN5O2ymbxazTvAZUUCbVAZY8fz78N92lQgeA3Q
/TzToVLWgojZcjn/zdBm3IJgTPpLqv/BsiEvQiNgDEhQ7w5bHScGm591SPApbmV67qLqvKbjCsz0
FvzU09eZck8C9dvDW1Z1otTkUw70f2EWIWFNhE8A/ltvT6r1NE+8ArWXjHCKj2ut03tAI7+rVLrB
7BxidmmAFOnxH9QG0JH72hEq0PYoV6ug4QoLq4bo8tvtAdZxiCDSn9BceFEVvmfqmaE0MFy8NlHy
588e/4xEoOF+Sn13v4QysZWVtaqSCfq2kNI9Cc+d9ooG9TXs6QjnTvMmtR7BFfRVJe75BprqHzBc
/ciY1mGpfCPvKE+1Bj4E4CQSxfEHDMh3vgUVv9+XPFU3EtjR3tHj4GuAs29bQJb4KoQLGP2vK1sW
MNTo416pJ+nz8UK+4bPjAimt8viIs/J1XuJhXs7TnFlokDSmYVz+0X1TgvtspBRTFNfiw28e35go
4qTDrTNW+W2uuyvSE9mMpGXC+aTtZ/ued8xXcOy+llyOA+Q4dU1dOJgybJY/8Pgi1rwXEW9GAI99
TTgFQxX3aOZNLA5no5JdrOC9S6I25hksYCMXiOPuwfmLwmgMAe5KOb/+64Vtn+62plReK4Omx1Bn
2E/NNm6CP5I/RZIN+WepZCAoBzHf/MuY2IaQKaiekB8NDqpgWRfRsgG6A7pY/GcUErjO8CeiRWaG
y/GtoGmMPOn62M55KB8SLCsF80EaM+Rs/Qm7b68VDAWY2WFtgeqkbrHcAqSfj5aC1grMObobOi2Y
d5s4FHLunRJVePfY8YnfxrnRS597DVNIBOA+AuuAeuIfB3DxiNvDNjCYY3pK3ycDWkF8JqHOaCs1
8lnA4t5SE9kpCuNgdgukyMF1Nlw9Nu0hw1+Iq9aN5bBF2r+60oHuR4BI2BKnGqKhrU74Y0LDL/VC
wdBSAFOGC4CrqX7gmPKhpiZxXIPJXAXw2R/rTCnzEAjzwMTG1YhyZ2Gly/vD3nDy5yDIQEK8NfU6
bFrnUytJYhLrjx8nU/fLPpMYbLVSENNU0dEudcnlqlE9HfkVrrVluiVNCpZXFFPtj4NgMd2s/0l3
e3CJxjm1EaUhigib7CmoqqyFClhA+UOCEP2PvrtwNOnMX95oB6kXNdlwqCpyybvsTbKQae/jTlLm
4PjGGdPBxkR/6NwOlgCqsiQ2fn11wyEhA3ptxvf3RqcyjnQQDfD8WKT0mGuMMT1esaJZIpz7s3Jg
tgJ358ES6NlYW2Wv9BqxDf5e502JwTZ1RnS+wwgbinVBcs3omT6oBKEsA53PDFRQFKsrwlZKyBkF
/ref4Bx7hxCT7LZRF0ATrl3XdQwRnxtrVxTiyeNiE4N7aySI5rU4AcNMmFbgAzaFAbyO4I0veuSo
bS6K9Bd08/v2gCiQN2MgMlPzzWR0UYT1DySXXbZIRfSLB2KFKSMGlizv9tBkEnOpNFzoqTlWAM0P
m8HCUcmHsgnb6QAw3QFxVA5+vW7XpC6+C2EVS6Pvn7jMtY7oA4aOy5l+YpD0em5GWx/xxSKOIt5A
figmjIijhpCkiyzvpKUV9Lz7P721NS5M4ea9y2jm8WCMZdqowmlIKXDxgj3AHdtkHCTFuPkhUpSp
k5rm7ynbXsaE0kN/vC28ST+uohKw6UzegLAY1UHzzlVABR8Cwbmo44JSZUGXpWdXNP4rdD4tpr+Z
bNrIX9qHYyEC8z0PME5Sf0fX61YnGg3S1Y/ATZBPQGg1imPvGCR4KxvCPQwtd4++8sND7oocQUtL
vKm3rZ6Ae1+epdKkBj/UtoiT04bzvWRzbXJUTkRleZFCIZI2Fv55mFfaB0nQNZNoFmGeseyIw9QX
gFNkD9yiYI14D5cUV/L+yo3wl6hD8mtlZyVr+YzdiZRs044EE0eOGaWPmQyxDaRFxBKbtygkwqql
AQmdjvp3pfcK3gYFoWTS9kkBu4e/13Wo+j+NLTlQd4t4pxDmLEAVvX5sEDcjgZnmanNJp8KQcStR
IfYxmfmPGXD01VPdrJXtjPBGvJDhbU7SGSPRTTcGP3EFpNFbSsIz97cAAN2k2pBlZLNPItGxvO1/
4qcunja1ghUHBurnGlbTZqYB511MTJqd97E50JoYDxtxE5kT6JYS+nAY71ZzMQ8x9JMyLGWYwTMI
vp3gJpYtVMKIfTVHgjB0AFoxPZCtA9ujDUbxhY0U1FwtUlaM6zoDlvRMplLG7cVi+XXFlTxNWKq3
83fOlTeUvtMsNRx2VwNEXLGqNaCgSSr3zl0z8uUsAjHLaF+FSKR7yk0NIPwGoaJ/EHaJDhwdHuTc
jk+r2AKzGsziqqFfzeV0a99kkarwBiXONGzS79Fx/dSbBApBGVZbR86Aq0amTsYbWQn+zc0ol3w7
0+WOudhYEPAlyiH2kle3KOLbfhQJFaOGuiAufgrcqzOEFk4xOyBJJWUYx3R3sOvJi0O7NXM8zNSe
VlxwhhXPNWWaA7oKVxEohfMnBC14iu+oeMwehgU5TBlRjUy5aLdFnCyMfF/gQrA9vtQnUivnGazz
YyURQXl0cOrO395gtdCwy8ubKkls8P6sWljhEXZxn8teEadHkjTtFR1Ig5kyweIyfgRAkez/7P47
UCe2Eqic+13zdy/cRp8I8sJBdXNwVFbLUuE1XRwg3FTRNgYlDovJGYrYZbSLk8ovEp3D1W6EoydX
L+2Y9QZi3kWNlCjpLZDb49tWiPxDcDklKMQBa91K8ijfffp9lq+OaWUWNL91pny0DyA9IT93tOq+
IpsoIb1U3osuaiXZyscB2vxhxOZbvQAe+lqCLfyb3EHsL5dCzoDZlM8I+MYol/UuPe1G/yn9quqo
uwBurNARu0C+GQtqlYqYnD5b5fy2E+i7u59g/sQMwg+ehloIvNuuBPwtmQEHJ14H1xKHj0tUS71/
gcFNVyGrV86Q/VSWE+CbhHZVpL+lkQE4z6IIEkimVOYyPElmLCKsM+heliCD+4XH15p/aGZIOgBS
+BGB0IAwuwTNf1eEMJjfp2R8WL6nLvWcaFZEeWWh2eCvITgDkjR2S/yP4Z64NDyssSQvwdY55/EO
Wc6stMmudb2DPR5juLtZFjpA8UiE7JwmL8JuzSh4qHSVV/xL/apPVTa4YiP5oRX9kyThRYUVNL3V
6wYZ/zFTAjB+i0lvPl1gPBGspj8k6YgQvWVXGAcBCuio7VIAwXFBqfG8MTAA4oOe329uLQl0/9rc
T1ZVQPiGXANzf4mGPSmtEalzvp0jIrcW3IUbH1/8/XnQTtE9hXvsL4DGVs4pjzAYvHjuEQLwT3Yh
48ntDA5T+574TbAKhkfu73se3jAKZGcyNcYH0OIds0S51k+65pUWVPqm1GdLN+zh4EjiGfyBlxdy
h1zBAdLr3Wbo9gxSLinb7bCzhEJRthcq83jUp4y95Q8yf4BWb0voEWTlZiU9NtTw528ysPZGopmm
8JGmejc0aplRYy7PLJJCwpQz5Fe6R7lkqp67ZeMf/xl0kf0MEJ8k+TXTGWRa9bMmqfZHqIjHLwXO
iFMz7QgBZh/NzYmc3s6zHhduekRR5n32crSK8GhNJxKIOV55v8WmpAKREfsI9v/OFDvr6ujgIuZK
Dga7nIBTxuEeGIFRFVWdqbMLugnnfNsDnmdlePIuXeGCH1ylsj+5nMP2jozHj/YSnu+rOkryHcSx
Gfy9rZQAl3iYdDk7f/0QHh9+uTkSH7nRpx4zJl99SR1iZwmaJV3TE6IRZtRvXnxRH83VCUe2y/ba
zhj616TuhedhkAaJGcy0dsuW+jbFzH6oPg2TbSYt56DzQ7mSccPt2ynAYAiHEfog3spaM7shidA9
ky3UJI2llTreBL+t0yLcW0UVKlZqECnlLK1VrQE7D10anemDrxwa1UNgPYL3a3ZN8zV8fSHgtMtc
G0b0iMrDCv+THNgEloe4fsIHj3AqWB6KlwrnQavj9ewmJ3cci6TkxeeQczZFjgHovd4ufKuHKjMC
6QAskKc6tzW1flZKgoXp7zZzlSBWk0nSqyc59rBaCW6+c/uxd+hKZOpk4ZUr6UdCX9nVrpIsql75
65anQjcFmXGwVBCKLmfngo22NK3BAlbD+li9D1zPasnWZcBfp9KCYqTkKWijm2yuSOqlHSc10lAg
zkem3Ux7fJrHa5tJckZNcamjsQz1j8ElQ1Pc5hE9kGOlJCVhw8OQQCbMhNY73obO8jEkODdBypTJ
p3ixj5kGCsbPR+Dwf4EhCgWMLBabYVK8N99l7xkWyJEXcRVF4is6D89IHA2JY7d4u8qk0qFZ12Ti
NAfw6ASf4QjpJ4LryYRV/Hw2W0U+C3q5vAgu01vMOPo2qsEMaWRtP+nPdrWmGw76f0DKJLEPDUl6
4QiVA1/rkdDWu+XeM81fh3GxZPjOa+AYHg82ncygp0I+CME3xK9vgwKz8xoMxtaM1HLZjBFAb03m
qmMbTus/H9PsRmK8Ey3RixRQhn6MhTE4yyLQd9Zeuqm1T8GayboZgEPuf/u4fyEqMS30qSb3adYl
mNzIG/oNBulduYdKFrBKdtp4aVYNXDypw/uKTpLggH1gvN1zRR87cghfwWIbcZruIUk5ttIFH2rV
Rqg4MpRd62+pYGIVvK+Ji8UsGQ7aR82PE71+DpsAvOqt49H6HzvM9afBr6t6bul/KGb+LJVLLZ5c
WJ4hHgba678LZljvDnY9s5PdP8X1EMeW8Gb22CY698Hb4hab7KHaNs/6iLQ88OzRYL2jzZc35FUc
ckoVGfLhMhhiebZooC7Bi8nrMniS/BNjxrdfhUktYQnC878RPZmri1wpSsAb8Re9i6y4Te+zkG61
/PvGLvnUKGKYgbHvXdqHjHIbCvedT3u4ssoAHv24tvg6CJ62Y7KjXo14dP9Y7dRPrTgUrN8Ogta6
JOKVtD/UxhysFFBcLFrV5wYIuyyqXAMqe5PJ0tUIN8ZBBVNHZZE+P1deNtHLNYgXPTbdQPplJNMq
vSjUMAHh6CbaZfEanIG2r1Fupn5/PQff5+cr92LqXcKaKnO0ggXTnxnpGdJ3szO155fD9kBqimfp
07Z81OSq/eLvKuDYT4niOCb0P0M9mdtQSAsyvNxySPBfzGUO114KXjz6N9ueq6cFCi3nqVfCgGQa
VCoR29FWlfPAHJU6BE0hYMfCF/QuN8mWQ3NdtW8wcJlIViIoj52Mrb15rUdoXeXbzprJXZRC82yr
UYTZ4seqefEf2f1KOEMzvsGQKgSGZ+v3ZBulsVVwKrDfK9Y0hocT+YOj+yFttHD/Vs4LXq/EA9gd
njiS5ON36Djuru9kHCOInr1IO45NTfWrGUf3IQxlbPWkkhVhowHk2CHj64i33p3S6IoCB1wlMLox
Jyh++TDfuOfYjtfSusuQZdNT7FnTVS2tENCNvEEDxYJSiFULSw5QKd6W55TcQfbw38RHGsRPwBQB
S0M6vLb4JqdOUrMaIP4tKJuDjpiHV7pJz1RA4Imxe3FoeuM5Xmf6T5RqP+tmBORmbJuBF+tvfoFp
bGuiAfLq5ts3hlW+ySVYw4vBTnbI4yXwbxDoMlR6XKb6HcIkcGuur/eKzrwIeeu/S00MkYuQ6Y9+
4zk6vpr52tSv3mW7h8Mm9T6SS2P5kkBqO61PTzfXa5QV+4v9sZSXLkx63tSjZK2X5BNRC6Ig/rL6
MHjfHIuMjBIUNGortbmFoG5Dnf/8va307iupdrTmX5wtTOsHo+ZO0Bg3IHtt601qsJZiehiFyZoS
OW2lo3ewg72C30Gxyjqa6ttE3HFNzddwUeBzoUZZamqqBHUgkTB6SfzlCeJL2MnPCWUfS+fJBHTf
RgfFbLNBbVBHNMWSogIzolbFzO6sNbAw1q6aCtnNDAdwmN3a+phQIQ7RQsf/mBLg/kYmH2qnNbNq
Yl5zKutJtkj4IKPjXUSYraEg1RE2XcDBdqFM4hTGNpeiD91pDbG/8FAr6zZ9EMYZEKV4P4RWwYkn
8Rspeo15+zGZ0LU+nyCWbiYhlSQI71rzva454iD3AU8vHNB+8M9tPywebqY++1t0pOoC276G6NwS
P9WtLBgZ60DGyHBbFFNTckW9dAePWXBNtnISSlidaKxqO3135ZHXbxrkS45JX7SA/8cQfXR7JBQ9
zNeeup1RHVMSSlT8mGlZak4QSWMX31dLIhQsULPln3H1yv4DvrhWRpvOKJ7kELqmo4+ZKEnUuAOh
fWJLKvkgSp+UMRjzyWFJqUf72U+CBP1jcSpYOJqYt2yMPD7xjsT/W0qMHaGO/uNdr7P2pHzYJvuQ
pEktJaUv+z+BMNgMNblyP+o9X7WIeKA2ZJCLNopaik63bk1SD9cCvt6rc9Uo7efI8RrYyJKqqycC
RGAmXGtfnygBbRIVaQwDDBUi18vD3Roub37aC7Qd6vJYOOLtgs36UhVrSk+qQQiASTYVG7MDtpdL
9dL9SSaHuJg9nw5GjOVwlJKs5oRUsKtInFg0xaRvr67qdU71dRluewpceVBaFGowKimyPFJCY8hs
fjucDf5VwcSDT6Xaalqr1QIxz7/H+QtEkC4Nkutkhw+cJezBwJErQcTG1Sh8/LYiRdYHN6VcqwLx
J9R8VCJcZ+XXUja85f7YoeO1ioQrEiFgjFVmQkgu35wIkZ+EsdmFiB/cQvUdciHDPyeJKet/9W0/
RoDiBmIwgKBLZAYxIWf85ANPv2DMb1AzkCG2tWJoU5gt5x8THdA/5AKNRWjJy0u77RYbeOTlwja1
rJV3fivVOk8yppg13gVgxCH7toF3eIq/3nQ+rQNczf8zGpVavtQccvjg7W3Acg8T+86fr+V28HhR
VdjTAKJ5Xc2f+WLwtbgWQOjSqZ3rO03RCup/MFqWc47+zDOPvrTAzy7cgkWoyDtO1JH+N/Ity/dt
hKJJZaWnFUbQT6WB/1vUPjpPZWacnvcILv7GDjUEJvuWecyD5oGchpq+VRTt41ss211xcv3eBGW1
brsijfUNeqPFsuRA06ejjXesmxaBty6Mt6wD5bXHW4tziaKR/tGPuOEcw7IsrHkNGGl+S9eG7Ght
R+b6CLEVuStmAcfMKH0Npi2J6mXDPMVWNFSf8sAXsYk4EtPOY851QbYPm4ktmNww2BPq3XuE/3FZ
G6l/tlBs7thU74pafGfKC+/A68R9iD9ERYKdirqlLJelrvtIeg1WsVsmz1nWm85E4pYbmZEDNdY2
Tc+uyQ/gI7nJYrHp3SBKy3UN6BFEvHZ1/5I6GFky23Iu9LtvWwl64r4DRiadQ3idRu7Vpe4JdLUA
smPStjLSD0b4HV6YISRCBLjhNThFFDEno2GkaiKsjRxMESMZBmcYzcjPCtJSTNZaufqHi3S6WbP9
QOkHcn+vB3l2eme75EHhIsyYC78Uiz3z8GyKrm5Xi8d4BwMm6OK6w9eaBj2qBMHltG3Z8mXXAYXQ
zhO5ZB5NU0QzUAvBY3mQBW6WJdTZZrgJbcKfsyqPGMyRwzG4Pw47i4cKfsMU4C6IwUmcnBRpZy7d
H6fB/VJscj6mv6aGk+CwR74jV/ZmQ7cb0WPw+lJFNPgfd1V0HF0Jw8aiJEVXP0N711r1c587/l93
2YEOqbhEu456IUpltTrt5vnOVRSjyhnbRZN33FEHuKp6G9IfbLuq1y+LTPuBRlQ68zI9azWDgTFk
6C2QLAUNj5mwzqHUYz1qT+DWNy0g8Qzry0xDwpjLFDS45eIb/sUkiaNZr03f55SbFVg5X+XanseN
XE4lmL5e5xvX9FzHqKXDwVpwSPQZhaaYXmPXyuCRosOA28RKse3iFsvu50bU/KitrVZ9F+12J6OY
zmJTs7N2xigSZ7zgGCfG1M2/PO6+ARAWmxqTgvKM9MRwCfjJnaEYgv+AmfGfpxHBSBUY8Re1/6Dl
JsYEEO19KMFpog6Oo65t+6NS7k8IhA+S+6LqZOY1izBTTS7SdbNVj3nEmz6psES1Kv2HXk4NHwm8
Szz2WEKurwPwNQLYkX20C2PtLR+WcgkSsiyj7hO/g9KucDuO0yBAlQ3AkzuR5UUJ4dxBLfLF/ur6
qYcJb0794gWrRVjRFX/ShgzKg9L55yQuvUouhKWwHWune1ZBawcX1raK+L55+potlSoJOM0l3Z7a
eqyT0YEKX1OX0xoKtpv7u7Yfii/UIWEBLSaP1DTOf9KOsVlwg0nA5g1i7281vDRxBbJ5+kg5YUHK
VGaz3bOC7ME0p0fLsaEfZPvP5+ZnijECxrDUxkluQsrteCI7h0b76M4MftuuIy1zcedguhxXsCSI
Zy7jnVMAPQtRPIyA9sRj3oGCVJosHab3f3Ctng7M37lynVoWyb+GseztId1glipPCOjABdiMIVSA
tll/4G9+t+qcmjOK2OVtr9zcxW3zEdZvWV6wLC/CvNmrA8qUjeMlAFatMySrmkYBRvde9PGKIIag
I4npyUOYWGFm8T4dE1lh8rQ2VfM13X3waY9HtSeTOKCdREKukEzjYTUlt3MeqzOj5SnlguCdRPkI
Ko53WJ2004QdcJ1eN+6IhjyvbiYoS9pxX6b3UOctg4RDSMlscwwaE6MeI97CvJqMlHrZ4+cE9pZs
qqy+GFZKsSuQFjJrbT5O0TBMmLgqypK4Vre4xHUqBo0zewh+v5952+oRL4mR7oObezOQ3i3/vH33
ZIcTbTP0Ph1eCoe0kZ3yYhc9CHXarlaDHqxE37OLbERqN4VbinjkD1rp6eKCZErgQ+zDAWUrUW8U
yv7MNWT4O5Um5ZxOH9o5+X4ByhkrRzMPU21d0hybe58XwFd0ZxcfP/n77IMMBs/k1sCCPRiqP1Qa
fyA55pBD5mGb+l68Nv8jPshg+PtPSxT1UpRyfHiq6H6hsziEmAbtJpPU2eF0iso41NfyhXD8O771
6nsrcdqJJTLQ/Fup6E8wPQKYJyFd7GtvJv3SioNO5rcEpOiZEnfG9n/XmWAsVzR0lWfoaXZSx0+/
TF9c08+lX8WsqfxJQL2UZftRpaHryISJdKgQD0YQDPgJNpLoljnBPK2q9ErkgbMYgV+t8dTt63fy
QF4cxCoVnvcIUYyPoEEkuYqx8S4TZTe52k8daMemecfZlBQ71sx/P24rjZ4wQQeTrhdTHPDaEHCh
TeR8b46DCPn1krIwZe/qhdvgx0VR9MQOlSQRMrSa0HE+2yzjoJBZdzvzGlVC5K51t54MEFib30hP
S0bZMkWOWgzHwFYZfqjQZeZFZc09VIHYGVvypAEpaa+32XutvufL0fl1KCgS46ydLKD4Ljdg75Wy
ijHfP7C4/T8viRQl8F50LsqcRDlbmeR1Q7Ppr8ORfCOyeIoF9sFdmjHIgOmCYh77kiJIhPvgXCyd
STSiX5fWdB8LP3nexGekEj7l+r9QmWS1YmS8e6SGI1n9Tvucs5ooZOvXiGCrYSY7q5gs608hzSHw
FcGVoSrh2wQqAAzn4/PHUuwANocCv3KwlZ/r6onchM0umiThXuvG6XhFxO4tok0E7Z4+AJ9DmjKk
dIDP5xC6dYXLGOl3Dbu3mRu2PK1C0i/8Tm4ndKejWkcOwNwshkFVoiQf6eh11upuewNfoWDkRsQI
VZB7XoK3npOyDLnQD7Sjq8+uZp7lRx0zTEhtBq9gNKdHJGPuBaZ272okfXN4YtotAtRFwM+phzIB
Loh6el/ukbny6vdXLMD227POTeD14C7qiU/nNFR7HdBvXZE2Pd+KbMD7ShkqMAqvlYSO57qTQVLz
tLErNFODpXSMJFb6u9xJUt11E+04tTcipdaVA5hzh3WoXBQIaUc/xdvaNrS+VtLevC60O8D4Jzma
B8WlRdBAmwg3W8QQdyWHg95fL/5yqLSkWDimGoMFjHflMo5X6uuGlQBsdxvHapS6fPmTU2yzChHE
4pRxyh3MPnzM4cVbjKCjUyFN+VzEpiS2xOU6TyFvJq97bY7WhHYmrsYWuceB11Aq0X5OIryDXNME
c/FzbvhnI7fox70WZ2ZcsrbNwbqBmZq/JCgdCGAGNQgqVyZ0Zuqr+9vmJN8nt9bQSQuqhKoQsQFm
7T2MbH5O07CgzGXBbzT4AlaDfPQQ7X12Kl1wQY0OWNcWf3WiQFolj3TDDWrLFEdIPhBPcpXrbB8z
DM4ZqPNNps9gW9oVSwdzcQ7RSe1xkl/FlBGg9leB5oLEgXRpQkwFxkaKeC47Qiw07zvNsLxV2CaR
YtQfoXhUqaZMptDY0a+tOVgU572P/GsrQ+1w4jvVvp/dIzT44rFnhLMXBRHSx/HLvZhVydL/dG4s
iX1kdWbueu3ekTv/BVFmwdvEV2RC8O0Zrnj1y/Cf4r8jiUP45N85bHOtPu2zEnStFJskP68X+7SJ
VwpoMJadJN/MoP3AAfKPulgHVPqqiIeTtj6eCSVWmOmJUnum2/QFNZ7vX0I2nxbcDrnvVekk31Oq
KN813vOVksRIQ4RBMR35U2/RQu6Ct7A9ZA9l5fIrGDTqqTb3Ol57UIh8bK8e4nFUHJ18CMX+A0bD
uyUeB4SzhgEMnxUqbv7efQ+fCiHZc14SqAPjMqqENRiMz/hZml8eQj2g33VDFne4wpNpUCyB/6kk
2eYlbsH8HNEtjruJuB7hzwrN/nNO8g1e38kVu9OiH8cTHEiB34Nh2bvAT4PJPHUmaqfpG8yFsacT
lnoMOzkp+oGSJ1xeDHujERdZ7POHv4HRneW+Z2W2TaIEaD1IQXLNQRGGXg8Bt+n97gf8eu3PHxI4
b5FynJHGV5JUmlZqDiZGZeK8P2IoHjF5j0Ube0JK15VuObyEUP5I1MbwbE98JWX7lL6PH24mgv3M
vAEHCtOtTQo8wQpLLpr/SmUPF7DnCPy1tBQlBL+r5tSRDKFAGA58ODEMs1kGcUoqEj+1ueSNUTk8
Pt/jij5TyHNM9p4ojOUrJ0Pac5+t1pb0VGHDX4yl1/6YzIUQkd+iTlAkK+cFZLj3LVXja8+DcTh4
EhsulOfhic5BWJxySyou0MImXsy3Lb1y8jjOaTzbgMZG4yHDkj8UuoNcG5cxFRGk0+rHItMnQKu+
YcRXJShJ8StvyGTaltjZXd0k4VGpXLfeCRtAuBwIZItjx2KA45VSmieg/miQBosa4SBzztmU+Mm0
oMTov/PrJ07DTecOakAKyOiJB7LrPsxUR4czcEd7GORVVUun6xg06JPLphZeT+waJN910J9i1Npt
XYOwkJhJvujjcpmEeQEs3vHvw22UcZ3jR+4xvSZIee+T8gFCXClT4xouCNcZSY/i3vz674/OjFon
cwhAHnRSZK836PlpV25g+gzo4aF0tpItD+v/FtpENgh0AY/SNhAmgXlkPRyYVlS6xa3DwUkVnfFD
t8r29nDiLO6QBGMWDVssQguhJEhCXrBkPSJZ2bxMKSskjLGs0on+Dl2yE1veP3TIyou6iSXu8yeG
V9OA6T7hXlqBI94gffAD16nFxYbl0WtTTBMRYuiZYV+OGdwp5LhjZBoOBVRQmvQuU++02WYNsPEF
cwT8Zqai73Ph7IP7nfymeStqtD3XzSHGZHD6U5Zl0IXA/EHun3hyKfUf+m5AFkftcGBwWYDwKs2/
1/9TWwnWy1xH3T7zWJpPXtxPEOO+3wxkQvnvO3Y6MWab30veTKr8qe8+WebWtHSrt3ReCDiRzhzC
gHJQnGD2p3Ym/0McqxUKUYFbXqtt9qWilug8UX9vd57PzCbCDI/CKmMIERvqVIIs0HX59U96oHKr
ekGdnGlodhowYjQ9nOBKNJGWJX+E1RjiWxJ6BJQOHzu0Ne6ZTk9KmmZQqaT0Ugmhnlw7433cLRMV
fRzpFnGABTfwKiv58+BCbooUmAJEzRMokB+W2nH7Rn4n/oy1lvqd/r018dd3Ms4OKN0vvqpNRqWg
kPz96J41vcUiBviBPFkNJKO81/puuXiK4d+6kmTpX7xtG81eHGxHNfWUts1W6lYfnAt7MDKAO0sY
9ILBsLKn45Wt4s2BYO7rePsnrXu0rDZJK18q9ugyFfMXCIWcxUuIA6zETlQAqp3zYLwYGAPOAAIL
MkXmtlJTmvO+r9rTcbDifySN5K/+3go9vHI2F+LMMeC8gS8ssQs7Tcn0Z5u3JBExq3YDCKLjT68q
kuWVba04O5hHDtneoKbm74SD5xNRm5QqCjMweS0cH+jrC86b7KVLMDW6wjn5WtmFuwTEu3MwhUg4
ZNrelOfdI/dsfLz56BgerhEZAznE7V3pGLDgpb55gzuTdfCuTQ5cYQC7h+mzidxUDMgD0gz8YNgs
qIJd2xlmEbtWcMTtl5swbEduhE0e36h8HOdwOdeLzv9m/HMAyOU8M+lTb9fomT7ovO1EGN1QhOA9
BcBDj2IKnzQS6hnA72yj3kA/zRpSzhndpz3MKspn7PPHOnohM5uocni4rw1luGJXeMjBAnAvRtTe
0XfFXEGrZzVo92Kwu6ep7ROibC2FHwXocORsuJx4gjWM+Ibl9pxJFilvFuPN1sn3+7QeViMbZV27
0M2IUgdcX3eKySbZabgw1ZcPasT6U6s8DofpXzAFx392jktG38p0/9JJHTssrWBBWCooSyPyr1NQ
DSw9eN/nsJcnAQwr0IcchXuV6HXApgQNFUs6Ea7311XrUENsvpVQoQQFCWYpIy1NBZUDeyEY63sP
kWsir1HxgMBSS8iU1bIr3Hh1qC94/C28FoqlYuRrbfoIca5jg5c2NGRmNvfMD2cZodTYrLUCjlOO
SViblPxYlrpl+VWuP5vYl3Rgu4nTsqFWFPNmZJ3hpeuNWLOJZ5yXgx2bMhqZLAg/B2rrzq9T6awf
G+Jq4IxWswT9ror6G+Ro45q/U5RCLCtxpPTxFM+uLtTcO+XCl7HMpXa1+YODPA7bIXayNsKtJ6jQ
L9cJqkfG071t+3soo4AR+j67d5IaUoBDJh396eQxILfsdF1DDa7opKpg1dslGB/3hsAKdCA1doCV
hyVavUpfQRCQGDQQ7rDu7FCp2LbtTgLEpomwsDH1aUMZ0Z1WsnNRUhJQhj8p88TTrTGUViFAyD33
UIMEQFW9fgT/hk7G5RN2D9Aw5mZfoPN4X2bCC2U8OksVhX+BmGxWMUFmZONSs6h//b6gMSMGYY67
TnVtg9AH2XSiOcODz0XlYHAz+4V74QLXPZfjOLjeaBMpG+Q1oM9ezSgwvU9n4W3VqfVfjAj1Ndjp
JeViWXv8IJ8ESgS4P2eSz8IuxkW/FmqvLPILJWaiylnfPxSn28pbBnd5jezQ2a1Rx98jN6fzKLSh
BRJzkEVdNkLMRD94hNJIIMJr8imZrn48HKIJbDcbq85MhR7LrG65x5i+yVAXDWutAu6KzgH4g1By
ZZpxmfBhxEfYZYPZbZAUiiuPWojtL8ccSRrH//hYFxJnFvbih5qr65e5KIlbfWCSEtEEiw5jq5o3
otM6dlUVEuh/Kxf/gy4h95dcOpS67KvK3CKjQpbK+Dlm+3/1l/OlwS2O0+dJGj1dOTsReN3Jws+W
K2QlA10W/oKt/PYf+qkFHe1GCJqZJFF+cj49N24ijQwiHgYlfEWayTFgPTEnhktzsYy5fAVHMLt6
7PGIBYKQc016qoX9Ly3C6F0oK1h+HGXrBA18F+EQn5tmPNplPpJgTdGg4gxlZgTcae5AEkb9mZI8
FXd6G4BmEvWeNyuf6e59oi+QC4uIZgbFImq1uSrzDr5tSF6hd7HGnSUQTDd5RYo1Cg6SK3bnuQz2
6Kq/9YemDVQbE5EVrJYx2hNvpOw++MOokpsB9D1VATptNWcFMJZY2p3SDsNwIgpQk56e4RsZK5BU
+2bmZucY/55H4l77XsYv/c/KB6cQXKFoazzjNO8eblBOAVG5DmY0iisD1/W9fiKOiJtGXl/zxtFb
PgEtsgJdhFhHUj6N2WJUbyDspq8mdCgszOBbZLm7Tiws+9hj8+vm6hdVmVb4q0sAWW4rFUXTWOTj
1n0X8O/O4Ua9vX3yhTXlpN5nWQ3vJoBZcmVpZZQzgHb6qOxdGZ/2oyH0SokWy6xW4kmuU9d7zJS7
zOebEJP+ZaW+u6UHLIi76k4sgmxVxt5CFFuIDcXSizt2ONXREfOpvJKY00XWtN/A/buU+g6ypGAb
RJJCs4FhFkE3f9o+ISPw/9mkkVM9W4ChY1lkZEh7cIPb+9lH0YnOXXrCdISVUcuw/LjPpIa5gJP+
DrXNTaivDLRtM9ngIIaf6wEVmIwDR0rQNuM/dcm0tujdx+6NL4zmdFiva57CuoSPnb8Y71v24Da1
8k1XKNE5L8KNFe9T0eyRgQfXNoo+gZxBgyeFDIEbqYZTYR95A2fYPs0AdOWswXzAdHXyJiXZjg4/
I0ZBKS1PnjkrSn1+aJKjaKPEmie2A5EThB6/u5Hvh1T6uYYnLticD+XoxpvEpCcBLwRrCmOk9btX
0InFEcK8ilN5yL9XPtESTT0+ZLSqVDMSAtW1YxfLTYSrzKm8bHq0makOaBF/i0Z8pgS5PZAlNAbk
OTCSvpAHvL/Y8oIiyneZu1JahfAK4nDSSjxkI/UkZAKVsKhtV+WZYgdPGVBv5FzcHBPIptQJthZj
+1DuikWEMqhdmAH7gluHR2EK9IiqVwJ+yjRYwfaL5YMeZlgdmausdZUBDEWC9pbLCtIkAPgh1wdP
pJA/WnpXf6iXKQK84Kum1T015nCYrnqzMSDKQnTNT3KfTGwoQnnjVvtuYOklKaz+gooevgkwzkwQ
J9BG+4bH0xqZMTGvPhz2gAkFbZdnjrvDLe8dSS3VTSOkBEwSk9cnR8ydTsrOPMvAadd1U02ZU+Xf
lW4SgSbepBI8fMu88TMs3egTwwBKHk0WF1kKhDp3jVuPGmvjnGSRHU7BnN/6DTm+ozBVLJNX1a4S
iIfQZ8pxvs3zm8Xn36CONGOc9NoYaYbtjL7LFDZ9KAYGaCMugiOLuUD3tnDs4bz0ssDLKoEb2b6L
HlR7Bkv7vHXCAyTxRzcJLqlV1neLGdDcl4EPv3TnB3WRBKQmuLvUDVmPq+kKsUx345PeLTWPRNW+
Wj3vftX7VsP/WUPceJ7/T3MrlEoHbUXBqcbNRpb5JKYot07oIJmdb6ZL7s6cxtGUd94NSS9SIBr7
IOeMBmoM/PGXdtcjQzLT9TQkjR464bvrQFgIHSjNxOvkAk8yCJ6Kb3iwz6SGlJyGOjWyOIzjDeXI
vMyDRvsEfHOLmLcgAUw6PFORy2bSBo9WY7ZizGd4MHsXal3i1jWsLacI3khNLtk91UugF4G8VnfM
iJF2D44t9WK2sH4PPUj5dewBvnvnCOw/tKizmPZoASLpRv2EOnBr4aHDAjq/xF46iD2y5m8ed4AV
ZfKbhQGz1WTF0EXpQFzmlFPvE25/jiB3yS9vqfeqyBe4uK3jajUoJFVe21rbg188DAv1oGR6FIuq
306W1wLAFJ5KRFm1DAyhTKd7vSAVIPFZadP73Jt/kPxDWChbKzQTSGv2KKaVdjKFvkQa5Q9aAGfL
q4OH5wyJCbYrUMRWVPc5B8S75GeKrZ0GkP1r2PG+bMsMvho86fz8KLFk4YiA5crvo4zmuvQkULQQ
A0/Lo8OUqWMXb6oCPa+Mb6ZJUhP5nHmzzuEAPLCR9UMwa1TTgMfL/bqrGQ2lF1felQqevthaqGTq
Ynsk1rE5rt2i2S40Nc7QAg4IGJ58At5T6cACjRqHKPd+9w33q06dXbtscApcxKxrYnQxeTRi6fNh
22mSN4Lw/V83ODbalRxcphHCMtWx4OqHU3tKgmbq1IsmEuVNsLdEFWN8toMPOqtEaSmjjwB16rv6
uByjM1MqWJmV+A4YwphZ++wc90JyHs2H1BC929ohw9wXPunvA4jbSxatXBp1ANHgNrWGJ8iVz446
Wdf71NitAykCE9UsXHQott+EGwWdhbG9nMdxCGodoh8BMyqeKa/e0fBwPz+vdcScM0Q/3RDRtxPv
g8ragCALEwojEzHpbGgtauQF6I72IyYVo7p0//Jy9uYGkmQkRT/+aQBWmh8lqmuSe8AkhZmldgxj
5vCbvhg+4WXx+ZncPeaYAxdkv/SM5xyes8mP31AEM2lbzCt9O7/pmyaYop6h9HwZ9We482gryoXp
F92y/wlgi1F1ZP9odZ0XMzNs5QzT9YTm8p+vFvLuCXl7GwYC7fnz2F1wdGITkWW8fS+DF6pOudCN
sK50Mbrxm1dlBhtVQyc5W7ntBMG0pjdz7vsitpq49jBr23SrhDDEXb+eyerrHhmiwmYgLuhjp6Em
4dbu+UIIxiIYLZEJyLwXScYX81NAHISlcXVsHD/CLqRp+08CIdLlYIrPW3SRVa7HUKh2O2RknvQ6
17N+SFcY7Nk8gOH3d/NmLmxJxYBpYKWkVCLBApB4WCsC2j9mQtFeuc9K3Yb2qubB36WPpxzkrfz1
lsYrgw/87qM1svoRkfgKwQzT4puLn7+2hlaBK4S46aWgl0xvyolhQwgmxVHzSD0fwhsxvl4B8S6Q
itaqZYJYAWC7pZwwQD+sGmiPMBnprz3P4RONGXmrI4C0gTqqJtIyXXAh98j0S9ulLQRjMhiRbqoO
2wABTEmHwzLust401ZdeOFzWH6kKhGvY5gSlDJ8nHr8HxwPOe1mwYllgoNUhG9fBYlCB9qRN2MMy
xyeRTPvP77zKfDGa96akJ69ufD5cXEx94Xh9lCkdSgC3i+XJFpdJyDlbvPTjKyM6APEm0/pNbrfE
VFSVXI4HxM4VCfGXIHeWMObbOm0O2MeU4G/Ps2lx0BbWfc5CHwtwcxWjdNoim8xcgWD0NMcLtSGA
orYd0rzVSx79A7lwgY0Pz9f7spPqSsmXI6qDLvfCuaOhfEagOsAy9AfSGVrmjKNy/oywdNaI+PBB
HZiQ7t46D9X3w3FTfvYuAPv1grwOLYpkzB/2n+VTLYd7wMTuqATStpMu32LzfENkHsd/o2NwK3nu
OS3zuv3IdkcJkEjafjv8fA4TTVhQdk97Y23rYiOzsJ4nCjM+h22ijcx9TS4bARycHqFo5PxiRStf
mu/2hcvEErOmluu/jAEl/5Ui9Ofcyg+spLtjqagSX1SJ3FlbijHdvW6Dy2a+vImDmoaUL1b/nHz+
GzThJSWOK1l78F/TfJyaqar3aimgSn3y6r81HNxmhfWBxZqlfAuGzWLAanWCIqd5XE32V5Ro22WM
WgWwot59iyq7oayz04rrWEhERCn7ehoonqSSK1hcYR1KnBaVvTUFrcfgfH6/yRsRyvC41VKDK+Ga
3yxRYVkqRRzYJaRFzHZc7IDc+5rhzPh/D99H4EOhNfgkZE3T4lMM8z5teiFDL+kbUZQDgtiJTWjC
z1I8kBRlxLjshUyaEA9GCLaBBgyKaWasyqJxtU3FfvWPRoXe1UTvuLcMtmwTGr6c+HfcAp8vj7L/
ka2L+PiJ1HbeE7Lu6UHCTMsrkfUXVEnLxK6WZ62Te6jkOmjYhnYTAVSOBQJIpSENLgQhpUqQfsVu
aVb28XOvnIl3uNF/ag0JNv7KhYIIsikXV1zdZU3G72yuHMsM+spHIGO/NZSNozq386hKcbbvgCyq
Q0wcdqb0ITqWLggAfYx14ECs93Wkva9plh6u8oL7f3r0NM/5wQvHDzc7Ia11NKDJ3tXKAkLQ4J/w
8AIPlSM8CVodOzYoqWJ9y2y3igIJI2seCIdFWtvOCPKDwkrYLW/qyZcr0Cp8xJQSNFjakiK3MeeF
K+igpkfwLOObng/aPoBET7O5uSFakohhcAtpmhkpIQIYJxfq4qq7K1NfuzKbQ0mUnhudgSBENOFb
g0NqAOR+PZqXFRsd6NUBKiXPKc8+YINFaJIwaOJ6z/oSwMRddo+x5zfmjzkqaln9801CcwyzsOa1
Q8ZOhDXuwDeRxSE3xJzShbcmqE45Rbd2hi6XmjTIu7bFhb9++Up4GHCJDjYOPIC9KSXkETwPKJZr
dIbO/VIjVQVe3h1fAhkyQIvXXdnk+tVkPABz5gtn/jCe5T3T4hoke9gt/mAhahSSP1n+25nbHbAa
vy+VSBdwBDrniGjPyEE3I4qH0LYY8pbsuqLm02vV1YF5BUm+qS9KmN9O3f0s6f1QOiFIC4ur7yYy
anZVi0RXUjrj4IRMdc67q++XQyXbaUgptRokTLSWPAMzxT0ppJWZliDrS7oNfaQqs00cMW9g8XJr
UZ8Uida82RTM6iVvmUTS09DACRnxw18uItgoEINcY+EbAZq7+cds2wClDKPEKkf84qe2tj97Ts06
LRqwL/UHoYlM5l0a7JmlRTX+7toyg00GsQG4WMTJiSidcYm8BqsLzbm8sSGvsf55UyYwuKolY8F4
auST0B6WCTyuG1dvucN0KmgBcECa7qj/4ObzeEW+NA//8V8iYapBGupLaduoj6KXhX2jq5P/p9lW
qS9HNGPT+ja3PgFPFmvsje7lY+42ZBAeu+qBfRGUJBlvPHZvCGKVUHNGaswPPpREI5YTirwGo2sS
G2v2XntUilwGDaqHJoTPvl/BWd36/Cvih6Bk9II5Iz3wr4d5cMwStw7Aux9e66Yq9nmzvfQwxLFa
65b8MEqSgVk+P2g8i8D7Lj6pg8iVVRLgXI77jvdPpze5ltzEZqkhUuIAvcbFqBC0ZwCTpJdTfWDu
T91rneqG6CGwR/fKZlInGhy145GvlduvEwKblUzF6b2xBe2BFjmJ268keJUCPogTQ1Jco/wEPZqr
CWORcOhR8Nvm9jLSw4GkhTqek2UyoHLlszlaZlqwNVE5mpP8lih0ZHDvujzHsj78FbPOXNtZ2WDu
zdyCECxeXOrkkpm3oP/EUMePxscpSbtUjw+aED/2OxpDyaiDzUMy3RK4JU6PfGb280oCUNFUm08Q
H1YvoQJVIkx4XbqccxshKAe/aWDYyK1bGqjc08OdltLN9Yn3MPNmvz4VlDGHeEDBGjofSRRmGnJ2
wmv1EILikV//XTipfRTrF6LZq5IfzvV5x3rMOEcrySJLZuVSTzyCjyjyM8vKjCALjNZuCL6s7EVU
iAKFK3vcdply7ujsFA7zGzZKc4VlBZ/v4Mircn/dolwjZJjIOIq5Y8tuxX2w+TcybUdpm+ol930G
44Hg8sNwrQ1tkXRZwQNUVLgQ8X/Dx5SjGqyZD/L9GXvlkee+/QUF7Jnbpz3sAzl8Z62wsaNxfGNP
T0X8SHw7JuWqSrIYkKok9PmJTkKfptQ4f7g4qu0GwF17ih1al5Y+STWghCEX8/qZv714bw1gFDPk
VjLbEa2IlnSoUzhbPZIU2bC7fhwvfOBSDdaRbZ1nj/Iv8tprCpqXWkwUlDlDxq5Z1Yvex5KCBuvc
hw9iXbgQRj7RjlzvvhBPkv+Gb+0smYeosa221BQjFRxw98xVMQmVY1Y3sCZx345WZviVUe3vI8Hg
EP4yt349+X/rVtS3HGQZemrbOz9xnLXjIzRtklvcVoe66SxpRPEP4ODZhMgk1g3RjsNtEFoKdAFj
4EFF0fUzinV+iC3GaAON+XcF3MqqQ3jyP0MPJAyISW9F5rI2y6FpxNZLLuE6BUt4CiP+JhLWAEHS
jl+ZDMfbrD7gegPZ7AhZOuvWWMohV5e5yM3S6Gwb4LVIuhd5zCCStIzgYYs6pdkaArL/KkQ8s/56
Q1sRofG0WDxbfM2xCpItDyHOwn6FkU+1FXWvp47/ZLQz087IR+nPX3wj1XCWAfJ+XDCIXdVZFzQ7
Oezh+e7fanSsWhpZJv8y37mL10JX2GrqUhYyG2RJf3oy05j7qwSNW0tmvUaaJ86IXljDXDMlTf6o
K5LZGFyEy/ZPU4wiGQ/1x2E4ZD4BKq9UhBO5wlrEkslGzl016npPvETIzEMlWkl2LrYWeTaFtuf0
EOpO6dfy3TSfmQ0J4LycxqcOs2MEiKtXiIWbB/ezhX/pxIWfMwK94EcpMLaiJotgUgAFZB+wxH5u
+BozVhMtRjl0vu51C3xNqEMFj2mHK8wBO1CEL3V3IeoImmBCTdCRUl0uQuOlviy53Po/VR8xmawV
DZEvaL6DaKKhcxcWrtCy6mCGrduCkPg8bSsivTixhCe7D+q3E2HlCBjVuTKUF/iWt3yvFrRsJQwi
as7EfUv2yztEEa92e+77pTluzRjmVn+aGBOATZpZDxyQLiuEzqZx7Mx1+ntKHE2Z0XWRQs3Caj3f
jnbeHT7spxQ3RK0APO45DUkvrpjubLDpm5zIT0Y8u3QJzC7pWuCWx49qheKFaWHGidmhwvVn+nJT
pQz2vFSBB3keTaZY1E0rwmSbrifErkB6mVfeF9HHgg6+mKwTK7m52Z9octrvjEwhrL4mJvLzZlgL
uDb+m2rWFJfxnoqpoo2SzKPjsi6OjyF9oPSUAwsvPSDyyAFcwXIo8RY23ZQmGf8bBltVSKHBKlm4
2qC81VDyLjvpYinp507EDUgKr5ZffNBhvutX05DG3aL1tJikN3dfYxZbWoOkkbeeD47oCLHtZhhL
gN81PFoX6ZIzhQt2DhfX5Xbk6ONM9oQgpx4VkRAbyOdeBaTrNToSv9Xk4jvCxviYx5XsomTSs9Ls
K5heDJ/0Tp1BnKWXUst8NAX81ZJtQb4EUkCMqDc3sUon2uKcRaH6+TIKscqQ/HWElRlK1dHyAkiz
Fx3pfBwbcuP+KMkP/6vyQvDQubBrSvnfaLOek8qUh91m5Fk8Jegj2Ju+G1fuQdlMW6jC9eZzkzqE
H7mAU9FRzndssmAuPBy/t4Y8AXZFIZ52gOToiI28i4QbgQswZSyLI5t8djWleAqRguHIhn/tSQG9
rMapxC+e7I8fX6SdKY8gdz+ltKC655VTj58lTpNwVd8sCIzA1kzR8rbmPJDf48UrWchi1O0v+sdC
qYWZ5s1QqYHlBZyvd04SSdrCrjzqFDx9xkdivGNXUhdXZ3P0gmQSnhrmOe9AYgSCeoks3C3QINZb
BE6JWmUp4w3/cVo8flrZ9lMJYdwKwrbEELlWwiDSL+rh/BofaYRtVXPueb/R2uotqaTApdvotQB5
tTox7wE3sCdj2BvJcGaafIud9ssrSBl+Z215YPH2DNgPGkpizySkjwtMAa4AO81bnPDPRJPat06H
XVHL46BDqij/cc/rlNcyWeq+kYza5+SCIDEkPwiJnadbgJkN0hyQoXBmnDFsBVKU7v72pbkyv/tN
m52RhV2wKTIYVH3sofQXTVY7Ld6HLMBkoWuc2QZfvHGm520JMjf40g+Gy/hFiIiShK11/J3usQq/
Qj1kQpuDQ2AxDj6EzLSGaXgOUX+pi/xq+FM92a/F2h7p70qxkg8I8yZbMxYKjFDEwz1Pr6vuNPp6
taB+hvGy1o1WcY7PcAWXX9Vkp3Ztaly71EPnmaFULf2I5InBvF+vPLNRBsLD3n/jyrhcy4YaCOae
9BojypjT9rMl7SBAGh0w6WDxfo0gGqIoP5xcbyTcAvhcQn7gR6Q4UuVj44S97a+uENWeEDuiNgoW
/rPt6KaZPtkXVNzj4iSYIvBROWnZYcTwWid7z567TNZW0XWyfFPgRvgVMHcLlrzGlw5Ppt3DScGX
AIly/19FXwslr2HbYEsD9+gdDj77g1xFJ3OdVgjiPSOPfs4ffhUfCnllFG9WkXvKu5iUJWAk2j3N
xTjxUFWLNKzG8ZG4lgeZsyrKbFgv63PQ6kGs1GuYeTGqVK77M8rRnSWHhh4lrVsXGZXeRDISJ8N+
rcKUugZPRYvBjRumpwhIsCBpLmjiHEZA2bNrPeVqr49jaPhLti7X0QTDgEvEjpumGV6cpiRz2nMQ
tGT68qq2D5FnKLslEc4IKoTIfBdjraPqNJAiMUr4ILNtyBx+vxRQZl+ObfE3BzssiPKNAXtNNehn
PPqBBWHyLm7mcuMn3AA4P0T69MgTBYDHgGPi3QN0NAo21LaUfw1uhrPeroTz6/mLseF448wZwEB0
iZwJZCXAlJsvpAt8mA4D83OwtSJTUfujkDukDykh61/NF+r/6DPUa2HGbeW07dJeWX35S0aQOusi
Ak57iLJ7l4nJKSFcIfj3GBP05KMeH0Qxbi8jcg2Eki0NPCqiwtklc3gf7djinu74rCpQPuV6dK/G
kvPCZfNJVduixx+vMAK+jFhZuXwB/WGZlS6+SzIbqSSvrT/R2DrAanxeIUFEYaNRQk5hDb5M5MQs
KDr8620bbsaBv7iENzfrgEaWpBKtSsfdDyJfNgCvg3h1bg8guQGOafzSifg2/WttPWLplWZBrXDz
/++yR2oW3xQ9pUGoNFSuFbnqpZGBPD53VICRe/DTGRRkCDsuU1Mbk4vZik5aVO7ceLtMpNbag0Mt
RI3rRM3TnX3IbKsNyELjX3vWS7XJ7GOWog1K0J18kb4uwh6E59s4a+sTTCaR/6E9hW8Q3EcWyEZF
M8OIHXWiVCwxeadIt9a85xkroCOE64PMpaf0Wb9j8Tw0njWTqAtrs+zE4VG5qM0iLeOvDSMOU7XC
YdqIs2/fn4PYyoGoOLl+AcniieIRN/EC8OBqx7PN6SmEHgW09ef0PA68PqL7aayzP/7eVRgLem40
TC9Ars4HTGQL4CQ8hYb0U+hJ/wymq8t7bMpIcrsXbD7P1WRgF8IhTMLRKtXXpb5eeRZJByIW8GqL
mvnxNOSyBrukUM5alaAX9asB5Gv9DiZiG4x273SfIbYWkQJJNMGQEVOM3+5JKA4L7emcN0nNgrev
nKKRoZvPI3SCMrhXeJhIfkfY90I+jUuZHhHVGzQVDQdRT7wOwaxCxqSk432t/DTRvfujbU5lOAuL
tVKUG5b986wIAuLH7Nc5bn29dGQ7pwfzYnFdInHoXjkKx47z4Z/EjiPQo3X3e015Y2i+Fs0Txbxy
1K6Zqbeldprv00duudDhVLS3Y9XBlEDqCkHJR7MwdmtPePm6DkFO8a+jZzedL2fXUzoycOqxk3lD
dqAFDzKsm1uyaHzW7+3aCoBhoJUHueVJdiL5w08j9+a+s2H9JhVwQnTi5wbHN4Xr++PyBgp34fRB
xAq/b+lhmH1oAwN6L7cAWQcFCxNcKOvzObHz2guSGVi9Vatparwa/yy5P0QJEblKwxP/LJY5YMpq
x3KZWKEboGmsi3O5V9D+tPioglTiODKeUISzBI0yP71yV7AhzXn+YxWxU0YjF4CcaBL4IUwrV+V6
4oSwCBFrncb+5xh5AcYB85RuIy131xyl7/eINdMdee06D6PoluFfMAOISvcJH9NjiSUZn5YqCUTV
0sZWVj0WdtKBsi+a+8hjWHXv2UNaGsdTeaVXPxUk39BWGcv1grzhb7OM1xSaR6KskJbvlaVbSzxp
Nr99t1CS27uLWsn2GWkGWhvw0Smen4n2CIe1Jp3PuyIe61Z38JJzZVTnv2iMRD1MwWopcI6L4sDe
A9RuAsXkRl/M5u3iGm3tD2r8+kLKmq4UJ81JUlGIrUp5q/3uEQ/3rnQ48aRADJlxxRVmuVDtmKb9
wHwGCKf4GfvQAPdMsAqp/Z1rKoW/ZbySu0l05OHYUOIXEAhRO3wy/8DlMRDhXQ4oDFQJ9jIEKmCM
b/jotuYWoJ+LnvQLtSwvU3XajOBagc7AVwWvzzMxlwetL4jKDMx/xUTSy6L37u1n04fbvwf0Gegn
kYlzH91mQ/eQEA1JUswxqUHPivAtnxJqtYn861fLy5WhdTCq+TnT3m2HVbVaTtwIous+UdVllyIq
1ci0/37wvluW38JTlAQKuyzL+siXELIORFcJvKSZgkFq2SBcYu26mek1pE5WfbOsdRjd80qSCF/r
1KqOoHBXp4jFx+2bvjj9hUbfVr/iB/b2PFYAyb/FH1oat27l0UnUehxSuXrPWlopEVejiNX7B5hg
wObphhsh8VDzH+gCETpky42BTWxNFEiPpmlTrmt1APrKpG1KqHEdZ1FGufuEHHBbsiPNkB/ukQ2k
ISwSDvEeDB6Sv/mDwIqOFlYYVyX25fzOWJVyZAo+XVmj8zBIaRlQmSYWw7gzWcwaOC+OJvQ9Xtoj
xICxJMBPL0/yMpgEnfbRLG87k1S9+YB4kCf+mXNSNmTkqJ9SG64JcD1PG+gTIzOeHlP4Hr0P4vDI
VFe1QO+KPAu9rXssT+q2fi5wqERW/2JUigXfUjbvyeJAEjtHuYWRx4kBeSN8mSM9ApxUrH1uQD+g
f4uF5gdsK+stBVbIolN/UoNs1vUDJo+biPXCpkYdmGlbG7PTSGrGdZMbE0g/lvSOEiOzz/j7s/sD
zKA/zUdQUTBctyBHY8ZsAwkBwVAe/V1J5YHLZcUexP50VDewslXEHGAYUF7DxxrnBdWNahlkeVm3
hp50v0eGitwfifKAnfRBNip82LMqtKT+0boW8w0J2nFNfJw06c3XFEzbF8WbtuW3T8ONUYZ+s2i+
GbWNDpyIf5IneXiHSNHEYgaBv28qwp+LglqXRHejPBIJn/CvKY088L8rMzCamLDm87LdxrRQMvb0
tL72ctMiV8UrAbzPkdE7kgEfrArXARtFEaCCoq6gUAPIy/f8BSw5hS53q04npe/XpVsMz0tZLeKi
fng6FGcIe63wKnBwlHKvH1yIulwVm0AGCGQjsjrRsJk+OCdOoaQPV10m8pl+cvzZywaUT+98wnRz
AK6jEUnyIqKLiqATOctrIwE/kPKyTox9FiW6jokxxsU2oYiNcgB5qTXihf3PaoTZcJlWVr8tUmB2
CEmVz0f2k+JL7+Cvi3nXHiVQK2VGB2MUpou/Jsnn53SSs2u2FPYU7v/J1rngjSqoOwemEKJ645Y7
WwMf4PihheHRH2kK80mcQ3zsC1n3gMGUoZDDbdXBEVz7/d7AbEUqGxrcJmG47orz4w9pUGeYa1Gm
uT7Rf4yOV8ihEmb1LAb7Yo+NQ7ZdTlQ5bEofUE5A8MTySjgjAYpuppe/lJXR6R/SAUbxmutMDpfB
pNOBiIiDNbEkHjnQgX4otxhjxL8ghGyOGw6dUnfRIvOnz9hdiYiqUCBbUaZ7DUmExBzwhLm4fW0R
8YqH0EL+mgB1rq1N32LiSV+AyHSnNlMsaFWn/ggS0BmNW5lq+OziM0kzPSUYyYGYGiGQ4DqKg7H0
skEsuGqULosMhWfJ6cYBD68NM+LH3xyfz9OxawTSYSMdOp5eLDMKLN6wN4ztAHM+EG3tpF36nljD
96rUhggSqkiAKp8bkx8Z+tw06GUDMqu8xlTUN8DBuY8DFk0aVc8Tn7M71YxyWrDS3jymAbrLesGR
/lrqrbuzRZdmHa2Z13RcErypJnf/C6Lgb4PbAyAWRGsF6i4cRuHORYRlQJd9DSgC1oF+neibQ1om
CYHcr+/CcKoCQLdmxKTWyzv/ujmYZxanRD4t/qszkPR8AVFNin4fJkTkRFwhvUJzzU4ihH2lcTFi
zSYgiKAX1c8sl5R7kh7dqZS2J0IaoMm73DCtSIZt/5H3FF0zCf+K70S/79oq0CfZLsdVBLyulKnj
D2YMmMek6U6RDdq1CNb9h0dS5A01ojsvH8sPSpPhwxIxA/qlXKBT6dmr1qONB6JJRPJ80n/VV1wZ
BavtWCLtlxn3DpibWF2lxlZD4AOHzn+zVSv0tPKFls3Z6ulF9L87ee8E7CmV2CELCFdItHzuEmjw
ZU7AWhrajhg7ECfr71Y/GV60fZC0o2wu5kWz3Q2XqFiQKlQw0lqibU0dN/NjVXgX/hy4PlD/HWD6
YSLYp4OgYRB5RN5qYSpXZB9soQZGWqdfDQpi68dp5AabMjMqGJkrpU+PeSEAedGmJXiolAATJgNQ
4QpCn4OTF7JYkzVXuEGXOe22XDndOfK7f1jmxcE+YvfzT5T5GL4KffhTuschX7of07BPzSuepeG2
yJLL/P6QEm+HkJnbp69Ykr87l8F2x3nJtlhP8THfOaTxxrJma4PAl5QlWUYW8VuclfG4xMM97B1Y
Kup1JqDrzqO1wO1I4akQ6/i+SDaILGmdKT9+nWzjEDhV/RSXjf+bl6kKVPq451jlqZ5l7V6ItvFt
oltHSmpBc8iNe7ePB0G/oMqqxk47LZHh9TC3/82lU+7eXrtPGKz6HNyH+Pyen7D9+HBka13qJWCQ
plUyuHaLIH2uh/td6uMnbCClHhbmWmHr2ajt9KFTh9JdVjAjvSDoLnDDxqnjL71ZOoubymJUepAH
NZjXT+y8JcLq/Og1Oovru2gQJWFK8gMDPM6j8Msp873uJN4r4Tx4xzgxRC1uXHy3uJAkXyJ8XMMF
7vz63Xt3jCYvfvsemDk5GbJLt4hrAd67bL1Mwhnv7KJvy0msB26R0IGq/vUBDtd7sbh/smTdJXeH
7mJ5TeINAXmQLJTW76xtlXw+I7A6YY/vzQzH6FzYJOKuMSuKMUzj1ci551lyu5ryjLypAKa5oACs
KCVzUhV2Zo5mjYqeHEyxbGinrP5xNtyH2uw3tqR7vXyE+eronuXZys3oz30p+ANzQ3nOonmyGZxK
dxTFJi5vo/E4jSEz85u3i0kh4xmeBgbN4ouEqEiRrxAu+osrQ2Qg36zoeMFdCN+UYjEfwWB89Jqh
42SuSJtKt1URJrT5ncypgLBK+vsg77i15+yD5Dl1NW7Nmc3gsHkk5u0aAjhZ3le6kZS9UX+BOwVT
UO6LgG0mOUstJoLXSsaW6e7AQMKZw+JjJr7gjJKUxmeojnV2oeM6ojHfFf5fsfeo3idvUlAq/J9T
De+OeLXoSZ5ZbVCOmjqqi1aSR/tQuGTSQlMCYmr3x1zP27VLN/WIbqOkbZcHpIZJ2O1tDJSTWWSJ
qqNWElLqruhcYEZ5zVl4MWr+SQa+3A8KDK//66eT2ti4uYdBeT9qYiG/1GtAwHSPJ3ek04K7ePRV
gBCzljFPjch91WeIueqZoUAJ6CAVZeKoxwbGFFe0a15WcfT3NpEDcHbFU8EzOsk3a81UaI2++Syh
iiSITYfcCIi2iokFIXiRlFlGd5QpmrDONyStS+VWv1D8UGrizuGdwuif1Gw1wb7k20iiq99gzA97
ocxTGwnASMEeILFx1uzJtWC2uA3IlCY2f5W0defqPc+u51LqLr0o3bRN+CslwqYqYBxrH3NyqjJL
ZlBS0d3iBbGVD4t1+2vqmww9gprk2DNOUpyqggX3YZ+r6Hkwo95ZoH34pkkqRUMjR6TqXu2cFMhS
UbfoSsrJZKUx9Bx/zc8eoLJzfpficewx9wm6hVLrGvH4Rq1WELr7pX7b5PRdhjgeI5aHHVs6xjeD
IKc4XwLSfdG59imR5ibOqnOrZKykprotVXjzebmdqaLTeuwvkBR5UhOlLwVJkpmPpIirvgafxvFL
14KJyNbuHo1bdtu2rot6ZTU29VYN/8FTvzK/yZMyYBqCaHI0+ZbfuqpshpFET0B4wT9p2h1NI6KU
RP+qylAJ6x9og7Hn5xj4FEOCsPGC7K8jPWejGMcshYrXWQpppBNn7Z3U+Aqzlb9AGljX6QrMa48i
0EPLv3PbhmzNZeeiKhMxvNtuDjZHRlK/mxu0NwmoYp3h7Gl0wof8AtDz/NlZS0ZEks3z/PB7qge9
PmItw42IYMCNjDtfqmDh8VewvkNlpJiK3KObHWOIsLfZ77vnOKSOzbWqh9El3FOT5xC9efP50AIb
wES8tiwRwv+LZj66/JKNjtT0bXV9gTGGQLJckoz+fEPvzPNVJz3zyuka4cjwU3KNV0UH5LnJPOtA
aQPVIXIf6mGCyEnlXyj7GsoVchDiL9rU+Wk07D6Hd5xAVhOSt5962MeIpzN4NfdcEIqe5dOztExO
jrNY2co+UYESG+eHTC1VulhBY/MjF9BPGxtTqzC843MhGbUMHQxzPZTwdzdxOxNy5MHEo/l9CNU3
r7OYmW7DxGJal+ps+h4xui3mNch4DMjsSbtkm9wC2QS/K0SoS7ke5JGqeHTbj217cAiIq+znDGm8
G4vO9pp9pYw7o9VnzLM7oHposQmw15U85H0X8RjJVJxJct7uKUXEI72qLOktzbeok/Slti0dNcrB
A39egBjTbPattEzNY6qA4G2QTdYxNz+dkwFPGxr4NOiGWEV2+6pr0UcED6Mqm23AUuVJqJb6qua2
3Lg8DXrPMbTmBK/lcDyAbrLQgeBPVJnIcB4Rzji+zacYfZXhUFHmOH3ZX8tMsfPMyqOb7BXcefQ2
Yu5A1Ld1RKcw4fyCDDpQUTzkgocOAUAa1NVgg7K8vR4kGjt38Uag8J+fS2rngMIghvCF2WVFHxMi
sAh8SV8g4/7JkkgyenHkkytpaelffmgoed8yR3fIeSiQnT9fwIL1JmPE80ZJOOS+utitYnstSEBm
DWj/b/xYAVjgsiVhfgrbNiQa9U3En559cFxtY7i8fv7cxc97mKQYvSTzG0w5k3iiWrASeKT0MpBB
g5CE4Cab8LxKpWAGNlCWZ1EjcjTBjv15F+M+XMLGVILGOeZFPghi1+vqB0HQezUsGaTfoeZtkKps
UghrFG0txGQbGJ3tFVwYQI3GUz/UgnJypFRg4FRvNL0a5+TOu0vre9jhx7WXl/M8LUmap6ioXO6m
aYOwdbWpG16XGoxGeh4R2LXSArD5VRzSvoLQxkqZsRYcfCxHALhhh8O39yaAzLlTwIvgu7hwY8r8
jkuVvNyhcojrdGSNIJ3hitCXRGIWsYQjPPR9z3tf3UZhFm9TSCxMIfmLrAUIPnkN/tsO9FSeJGpA
L0faUSe+m7Jwi/6KYn2B4IWM08XKAnrHJFXpCr6L8VvMVWcNwA7digbynF0p3PXecMrj/eFvfFtH
VCewtUt8UZYbFBCjJhL42yNVoqdPFGwA5HdqmCjxvF9/Fw4t5YeTKCcA10ByzHVwjkr6GcEVhj7x
dvpjjbMVwjmJrsdCaJ5vPyJHVlVwRrdab+X62rH7CsvisAMtavyL7Jr32BVt9wXVUkeqXJkZybZO
XlQxjH6pnxc9gAqJAdjGjTDW7AoZ59wrOTcWLl9vFtEg/R3EgUwdQY5f4lv10jVT2pkkKUHuCwh7
WVYaJXCkpOeJZCxWcPkE0Fn7oPF5d5x54PmRf8tiu3KbZol2Ck/vORY/zpqh8OUaOZrELbCEep4D
VDeGh6tI2UmLmA7t1qdiqfdbxoHrqdfzkz8z4DrbVDwwvp22xo/nBGvTksKO/V5gqWAc3MLxQOxX
n7cX6Wy77BDq6AXi0syhYvH/8DTozuA+8VI90UI7m9Gg4c9PsHs1VvE+Lqff+B/vplBYW+GMbetX
jdeJhdw4+EkW8csPH7SDPZGDPa2D80uZtzkg2xOR574ng1Ce3MDsd5HwpnmSbGqeKEaT+Ki2lnYF
+VlNNyJlN0YIW09po8EOkZ1J3ZSEPmlIXVoUIAiiwHZ8KzP/9z1sH3qQ+rWP5SF7UkLmLVSCQ7VR
Q6ip80G3uqLgWJsep2mSo2A3y0tgJECQWmybRlQwL539X4kY937dBPUCr2ApPnRx8QpT09KPsFXN
rsDeHop06WcYUYpdLCp10ny1RlkIuEUoLXtW5MIK7Ih5XhGAjz9C0u8vb+IFoHWMAElHHnI4XUiV
Dc8M3fQdS+m+JsV52fHFCdWMGFVEb+YJBTkwfTXIhXuQj+ZvyrAcg8X085qGLmU1Me63zxotdUiV
q2VT8ps8uXAMfg7bNOVDjsQ4GKGwEDj4Nqd/OyasF6mMxfUte4trXdEkhi9nluxtgKmFJIRsZnfF
lXQ1O9i7kzYVU0EbIIdppOB+BYcJ9zsb5LT2BAgHfAxHMmdWtoUWvaVsIdJMhbubXK8c/tvq3Y4O
EGNSjWnbA0XYbjP7yylXIYriBTCQush65RmM43vI3xc3+Zea7zppydqLPjIYDYZJvbF0iaJmGdv8
4M7l1/P25hU+ijrP3UIJbQ8r57JRPLPdToWZXRseJ4n0QTYvSlzK5LjlblM51k9za1kxPhSoJpz4
m8qjg4U5Pvhuzn92kimDyZNB6JptKZHAoVbutLiknKIH4WvAKOGtQpnh3SNu8IrsM8vvgIH3utmS
yBSLVvC/WNwzQZoGfv3TLOhfF+fiQ9VvXgueGQlnuRiKz+vv5XqXLwhMbkr6fCgE3LRyLD0hrAqU
lKn1wa20euTZCJ/Mcg2nsOhOnGsopX39sozVFOfCRDlgSGD1CWTB8/WqE7+JmqdG56hZH66EZTg7
Dp6Mtu2nfOCS7/aeD/BOAy/LW4i4MS6U6+6r6yl9AbO3WCDbqeVDLeTJ+PSBjXoVmGOcYbpTIqez
2cfqhb80kes54/fN0JHFPojliJ07ummXH1V/23V5YcIgi27l3Cm8o/YTJbDnSIlfoZgFCP82wbXV
+EVuzlJiA86GNZ3XLh0D3rdmWGhXpV8V16PC9fGpX+RzS5McDc2TT3R0UnGpHgWUytYOF6lzTS1i
AQsFSfUDvFd72NOi9X/4ZGq7ECU9OtXhASvwbF6A2LgeLItPoSafrfsPtmz9ndsp0xfClDowT0kb
BVjetglAspHYOnaj6KPC4xpQsP+j3SQCfTk2OHn3sK1wN9AfkaZ5KjXT3J+don7GDrtHjcQkUEs+
CM939tJ41TywZhHzUyXYopSIjnlHFsj2/CBlOgJMLwjaB0qby/z8MOBMWDFwwrtprY2Lz+Qbsuof
IWgH8p2AT53Xe9i5T1lvXGb4EKF0hIciiRg6Ayqt+SyUg0ApWYnwYFrufgbbiCGhtAp2BI80v1/3
6gR8Jm4VwfdHZOYsxFqIxCw0AYNqk+29aMD1SRFWWyaAL0pPCgmhZ7mUbNW7IEdU0iUK5xu3prmU
rWRhlC8GVenCM30cSJcvdtLJohdwRF5hJrngH/E2PDubhT9+6iKwcYv6MwEr2xibAr1XsiNBzfIQ
GoQhvcjYCCTVXXymLYz+7IdK57LGUufeDVifU+CKSjBtGOlEHsvz9Ii3eKgr+uZCqCk0VpW5jNsA
+mr/BKF7/RfBKxfbkogRwq9FJlqObMfU+VeuyFnngi+7nBP2Wu95JqbN/0r8djp/dpgYjexBqmDi
xTEgLNg1xp8/nNF6VhJFBe/u6tGFFfSYhcuH5ft4k3TsUXedWBSyM7Nm9nDez9kk3kjFdZRLBsAE
51hz68m0DdDjgpaMK4HG/p3UjB+zUjEYAJnn11f1Pg4C0t5vn05LGUrE8ctOrdtahdjZ4cMsWv64
dwSgVoDTWQcSOz+oWmKWJi5rf8GV8GZ0L9FKg6q/unYV6M0qQNH3LTrvzaT9bT65xc95O8nPio/8
tm3igM2AL2kVgKzCFBrM4X7zIHdhW93K+CraRKnryx6yyvIuhSvoFaT2X/x15h/D7ipt5ASJ9yUY
Jc38R3y9e4gs9P8cT31owxEOY5o9efPds7Bp0GQVuTkhOcaJdMjoLBMjm5B//p2AlyJH/aHqWlda
Ped42POoBspat8zI/npuMYzvxzNG9pKsxARVUV1GiiwKjKF3o61vt7Ac/8maz94SCPn0ua9MgPF3
G0MQKLl9mASSiH34kYr1e7Ly9QjvYf+FhVxcFPOf61+XHhypnoPG6sOQyMXWuT9FExnmBAF7atSt
I3nLetU5HMsReZNEJy0UO3htALvQuq1ovMxiiAmSSDp300abH4JevsX8Xl3950jvm0lsVFzT0FPr
I0ESg7hcMqvoBfTX9gW3udzuzlDFy3US6awGcIV3/8JJML09XXQ6E4izBs53oydD5P0WKO72pvfa
Z8GnocYsi8tlbQ5Hr9NJF3+FdMlq9RgZaijgxg/hqfEVgFae2Yspnh+npa2T7bPIsPgulWotBmkk
Wj6793drAP99aIy7aK4Cbaih+PN9hC9OZtkGTkntsEPiNJv0pZuNxSm5JbBwTf3UXhxKN8Rfg8vf
vosIfKGBgOKT8DSW2b3BWp+0gtx+Ub/VPP1xCJuNfbm9LS1cOjAsqtliEDlgIzztDXjhjXoH0rn3
3vrI7FeyHNVWjSJD58/x3bJL0G70A1tmFYct69LXiN+KCWcF8zSXLBZAHAt4nhK1HBTDe47zj8Vo
1sPZm5wYjJgohBiP3AEUoK7p/wdNjLBLDcj8HBUxd44cbZ2Fx+OnxmDmA/8hCC5on5vMzdqzV0/M
JX35TCSxxnlNOBPgyQbLhhEAexHNNGa0GS+ZXmaMmfpGiAre1ISrRFyIBdk4NN7Nu0+tPV32vvJw
4WMAOntmlh/Xkbt+kZXOGZ0tocjMZLquLbyrFKSEU1XDklfSAIJCIuGBkQWVnMmkEEempXNJTqSF
FKmm0IFPjC82UMce9aB/a1Ip1raC9J7sSGZyXt0QSSswBkVCly490SCOOxcH3LkpTAvZWl9YaA8D
hRWGGi8fDvh3ZGLZrRVqMe2QR6e76Ham3Aj2ptvxhyScT08MPmTK9UE9K63/SHobdU7Rn+I7w/1+
E9PVxfq5hUy7FLNn3+05KBcMNrKUbREZyNaERc0C1Qfe/gn1dmB2G5Mkym7+ZCB27Uvux2iT4Nce
DjLz+vacxjfi48f5JWS/pDx9khKhiP8RL5KPoqdGlyedUBP464pDiHwm+oFzMQeF/5Vq6SS8hN+A
tny6r/iwHMnBqat+1DfrX2Eocvai+rqyDNqdvJAo/j/hWm4INV5N8IfkEK8Rl67GSqtp94yFANoG
T1SQ/Qyw62fqqRsYv+kVokhuJ2JzzLQNtEViDxrU2fSzIrJtWzK5iddHuF5nBcBDNm1w4nGNXlqr
lXn+LzcdG4ExogifK7+8cVIr+cRCVTh20X1W8ROl465ZTVz5MqrH1zurArm6iq33meGyt/4ZHrT8
8ClsXAPOSu5MqUi/fG3kbfgbMLY4iiQJxurEl9qS/OUVxNAfdOQa/R5zKOFGzWbUctLlavFSa1o2
SwKTGiaUjD9+89sadOlNDa6+D5y07/sEnnr8MaEHRitrPZ6F+K4wMLX04c6X3fTJHxxXRl9f5ZhD
ORbr9kT3z78+DQHW6jYCVaZvxH+ClGrccxBCnMV7odIJROpO4xwtAZfbkgEUSyYD4fsb4YDfGiW+
A1TyNkg7dV/yKMyP0JhWYC1gW1eVleiDaLqelDRuosJeL92Ae9VjEwu5z6rYej9NcQTwD/3grXm1
DtZoxj8bSnLuKfufp4En5XQibw2eGkRxjdLVbEd91s7dBhHA8FN+8DVJi0+JfBon0yIyJFL63i/C
oedEuCoJBh2h3UnnslXpIn1HjUxOSjak9G8ZAmC9Fb5r9iuXUmQ+4SWbOsYia6xn0PMVCtHkN6Dy
iQY/ldw+wwRDg8OZz838vyjpBuonN4HpCfv+kjQHps4ZGFsKszj6VxWD0/+gFC8wKUer/NxGhIwb
jVWXWrlfcCW4JRxmdLIn7Z20zwyMEqpfwm6hMi6LLoiRapAvMrQLgCfrnJvXscHgunVe7rA/cYoo
gZO54XtdoJnMx2WI21zC6ObN1kK0tJA3oxdTmrLmjV3OncuDD83LjYkRpB0WdhTBxpmCLbbrEDqh
XqOG8UZxTcUCUC0vkgeJkTyxqGJfCJuy18hZYTHk8mjQwhf/HZgkgfVcGn/LaawrUx4aOlIzpThB
Tb0HTX2OED3JU45MxHjX7mW8EtCEDxNgc2f+sbNikbwHE6WfedGe8P9IGoJvRGfROAuixhvSc9g7
fYdSDkh5vjDQ7uy444AdcReGN9SQYdxR62sqT4eaRiEnUPlAXYJwUNgOrKooEQTlVd0MiSCtmlTr
EDFAImCoegIoYgwNjMHUQP6noK0P0K1HhN0LFfXiO3hqQBsD3ZrTmyIo4TIrJB/k7nSwOBFjUzhv
jjxGWy269Ro/pgrAA0MNXvv0cvOsI7IEEUMY6cgcZ3IVvv63wL3NPsYI1hIprXyJP+0UKizVSBHm
7vIPJRUIubJeY45A7+28LFJ7Q7EouMvJo8XEdt42zso0rza4ZbpndLLEL354bfRIgi8LDjHwyXaJ
f+3xwx3pq9NmCvFvTFthUSf4j2JWCB6fpwv/r/uFvA9I0VqTBpxU8HFc3d6tsrZzea/V4vctzICL
jt7rYWxdQms5X6VENMshtetkR2zpRzIbqa+pI/BM6firUvOTHtFJYwrRJxV3X9GkoAtsq2FENzTh
Rcot2Vd9K2fiagciUtCBlP/jq7Ibo/uksHFdHoOpUG1Un8k7uIXpt58d6caBy+9wW/PGGXkfc7/W
mV3n7w1oEAvMF2P0ChUGM13kA83YFw1J5SHpzVOh92Ja29LMp4OnNSBlEuMVap75daaGq4Pbr09s
KOv65oNfHJ5+Ufn520HeVeOo9TI+Qu7B6vSLs6/QI2iZAG7cB57G4ALMjYzAes7d9GzpxD/czqpG
9LO26f/B7TdSzDexMQh0o4HNEKkLIGOQCGV8qsliPmCX2MWbhCKdObLpcrgj7QLZr/9FklF4aD97
HqJmiJhoJKR56oENzrc4ky3KY2Tu5i0jYepdrU9jsBAoroER53ek+EXMhVJ+z80j7l2/gpjYI7dj
mhHlxmBRk7f4yeq6QKktDUbuq1yFU4he9moC8ClkhN8YWZZGPLBKC8ZbieZKa1+69EJiFBYv/fFR
Fv6upXJox4ybv2vuUd012JCoZdOPZEQSyZSYryD1stUAx9XYsk86R4ccYqv/KxD7tiQ1wPsAG50J
x6zE82416bgy9FT/4jTEJSDbUl4zb/jz3uPjBDTnZZ55AdJ9+OcTvdNKOdXXZLvREpMtxKn8rmsD
oCtAZ5Z8ZdWsO3aAy2+UpNXm0rq81lRP+F6DOVOGYeDJwqYT1EZmWcqnvpLhYbHsaweYyUmCqDVS
PFCtYjdg7/0I9krdMQJV4lRxFqq+bMcvPcj/HuwNtnTnSbHyK7YfF16xX9DKib5GBdqs8EHBF22J
9pmFTQ3oGtYCbYXRXqGVhfDOdpgN2kzYO5zVkcC2ldzMCgVBnT2ifY6XGcY8ldalYq4xPbNVZX9m
lYegWq53q/CjoYR2X0SpkKnFE02tN8mY/SWsAfvqEPUlyc6w/oWo6vnvdkyBrfZlIfU2IMfx0Ecz
bR94qoZ2TOK2PjDd9qslDo2jCrkBzpxHRtlu+ytPYPnmjZDw3zq+U2VSatkH/QD05vA2MZ1PQWKz
E3rvLrfrD7Tvc9BTQCaMsQDu3NJAd/rl4pdcZL01b08J9Ata2K3rgLE5eWzaz0SUdlMOR9conOS/
9avjWS+ERzhv6HZLrxbuCzQoQn4tGedDcDqpdOOQau5FWIPXXlWlJrD0OiaVgAwSKPBJsq26JZI9
HZZZ+YFnPUA6axrBO3LQe1Cqx3XyV0SsL7oKgnoEtpkTO7AGf8gZrpuzB0keL66gSzI12Qdoq1Cx
rlDExPeziYin2QSyWNzQTdMKxNWWREpL5iCeRmnuJglW4yuPz4uCygTYDP1sxPrxv6XEutk0lXeu
r2Sq8sv0vrd+z01sknZBKMeyFfTMDOxSWfvLFkMs0a37aeZT6T0Gnwom8UfhJ99c1+Akgclv3oQE
TeMtIl1teGQj7I+mWxhoG91KcnR/b/QExQ8oluudKhBpZZWNewCSudG/bfWZk6yxeDKeBvckKDQc
aBPcRa5p0vcYE2xy45rGlgRdmGK6M3jXB8DcHouWG3YLOtAyYe4ZtBdYmeaF70piu6Q9z0dR0C8a
v1Q3wKqG6HYmTU1u8wEIPtoEFCHezdxORmJmAvrjQdf0ec2hV8Mww1FhAXqlkbDae7vkTixn/jwu
jHkSP/GKVm1Lhtnx7jHFfV+DU9tm8yLglnYJqNlKeukRST7mzEvO+SmsHDUipLz+jbJxBN5HvMYS
gMW/zW07S5hSC58dUumm6JW6TYQgs8F7paFrmUrpfbHlma/6aE2/Qg0BLUPKRQm4LCle/a5ZoRjh
HIWim91d0BFPrgR57xQDniZZTPHSGmkcv12PQQTCqVUqMtmLJAIn0P4HV+LyvOsxmcGej9je5/PT
QZjwr2BF0zAnYMqf8ucooRV1Yc206HwHjg/+IIUHUEhaH1dWLwkrl6K4nbpteEiOsGwTpt9GDy6U
KZLr4g1ICp62qhRQYeYZcKov5rKIBU9vYqw+EPyHqDo41frGysCccSS5T7XAODw/icRPp319N4tv
atU0fnVyIDVP38AV4qx4AWX/OpZueGh2bNA5d6qvXarZxyMXy5nT7QPVQ0VR9GbS033+wwVBnqrv
sPvdpDwRztMy9faVPwTSINoA24+jrO1gC30aExb17AMigLHeBPE3Lti6PJlUPjp5jNqVt9FlVVzc
rg8Agtt640tJzvyJ0UD7vkYfgoA8u7qC5uNJxaJcrdEy14+uhKP07oGsWR2OFZnVQzTlYLakJTH7
Z6sM8CwaIsHhbzOPa3YnanBr0GXsPJzT+6zwbCmyQ6G+ULG9eVPqQqGQoM01UZzLLxaX55ijVo19
oSfsOgV1S9C8RoMtFHKqmPEZi+UWKCnGkLWMAy8dOLHqzci8SVfyJ21eXXhhD1TAKsfsJ6zteiev
5QiRQrNrXmdjNzh6Yq8OZX4jySyqxG0rB9gXEpYArktOIzigD91giDYu8cSuGpihtQ2wlW6t8y4m
E8njWe+ySZgLb7vOgSj8XbC4DbXSta/kgV3q7h3hFia4MNnZnH327XDpoaXo9PZhUqSWBXarxYTR
fRE7qMx1eV5QNND8oKxL6CTH1zD+8HfYCgeQMe50tfRSnFrCRCyj+PbjGf6t+B+i8RXNzlc/U/ea
Miwp2CLNqNr4q4PgtVBqLWcF4E+MdqpVxkeekead7VscemvyCkgnfH5bOjBfhef7Iio67TNrLiJK
iZnk49ZLda9e2mcgq7rTXDdO7p2mQ2hGUYLZogB72EFOJBUpBqZlIkR/ZZ6Mj7MRnofv6+4tBFKr
Go87cv8tKZ6ihkucr5b9whtqud6M4K2aDuTAaNJth0Mh54hVk1zsXWy2nZhJACp8Cu8UIg2yqT8Q
A8yCZJ1lyWViv+EeSMjrsWXzsuVWCYHfrjSv+RYp0GexUVB2AW+ULfUBxSYDUS7mdu+k/ifBTq9r
QuZPVYPva7kT45KC+4NZOx673boOaKTLNFfW4gxTnurcI9++5nPGdDQXaHQapXG6J1jZRjbM+pBq
j654izbZcT75w77n3J+HXcxk0J3XUIB0waiChE1Qk/kGlw0hUFKiPu+XR6pLxmpiKWp6x+igCFIp
yzGfTNeaM1oZinjvxQ/uFZTDR3sFPkFX6AWaERDfQAgTJsrKGCt5I5NFv8rSRzeytPv3juFuY7t/
dAOdyJhPf1DVOJNLwsoiuX9uHZ33Zc7ycNsN6c/eWQCLhmIbbsxardDW4RVhlzs+6xkc+N018Dbe
ot7KIiFVInqxLTdNMP7dkgP4kyH8sHjQCs9yRCGwbDRHuh0X/zDdjTjIrsvMy56gdotUmHaTpb5e
jrGShnLQBuNpRBEBHlnzenvQ5H5pYeS+9d9bMLCGu1j14F0UXf1jjE3PYDkgqDeeH0SjVg+2WwS7
i1yrRGvMWfu5jTGf1HuLGBG/uhYYEq+nt5iKzR4pB0mAKfJLB2k9OCn2kht1oz6RKFtG0HC2RRkH
SaTfqSuUhl8KirQ1ZyeCOTOiSmtrqEoZSMkzFr/icFPjGFDJ9k/CkxtQ/Whu03mIKzVIWn1kkbsc
vwjJ5YAgu+RQu51XxbZM8IzyUrRXPQjjBfbTtLy9M10O43kmaizLScmy7ipg25A8PqO+xT8tbG/V
QjEcvsPM/7RDXc3rFNk0jARbjBvhjNv7kzAdGRc9rDdS2nYoRgMJSKzgOd7Ktk5p5G0PgeNQzHmn
v4bCguVU9o86rs6mFzOfKYOI/sa0SV2Rij1qvyg1lnxkZidZMBlnElrwFEMMWn1kysL1rDPVPltJ
eFEik4QT120oXahcGIWyq/kD+W9/FehfQD47eARMZSPBOvxAA8y8gTTk0SvPIianf9gMLxn8BAcJ
LpnR71ZYF/VK2U1l2qUKjNuWsLa4muLECb/6DqWTDpIBZnzT+QHXz3lkLliqlS5NzSgDRjoh/UP3
J7ADHbIzdjg+ixZDVdrq3erP9xXWTIO7GNoVtJgLM9EfUGUKhDSxNmcoAN6SgxfjKmmGYW5qScri
AyESY5vnI21RrpAXYOBcx1RS07xQA3aq/MTOWOLuiutwBpFIz1MtK/rrDhqradx8l4elMMnFtK9q
UDtLHYmigts3zQnK3trF7bB4WgrH0FyZ2JIGlwFKe7GOAXUF3SfgmsjFMQTqC+VnsLD3scUryiq1
hIzvi7sTC2UCuGsxhAp1CC/HPFAvB9nDD3b+TI0v+19dFiAQtsBflYeFYEIMUymLaW/8bYxuyZCk
fp17Hl/kS8gSBSYn6YZDTvQBqnVX2YL35qLtjBNjzAhgw4rG1xcVA6nHvAWkLCsgpbcs5feRE5ry
IBQ1Q/kgWRXN/OLrXciqLtBYmkkoDOK6S3NoyTuPQEdOtTRK01o3uvsZ8U3FpFHilzQ4zIb/TiCM
WsDccFX6K+CYinY7Ra4tawQpBKlyGDqA+XhPvPgGwSV/le/umCa5FbZe+OMgSRAucIoa0tW+EkcP
vPDGqiz+6ZKWRMAcKSVBvq3nW1qOCdfTd+KOJJ3+ibUs7sXre/GNjZhqFEI1gBNosdkVKoE9wOtA
iHO67nuSlD4mhFNfTHKHREe7VQG5sgXj4Isefskxvxoa9ye3lnr2kUSuobIcYuBaF3/BAE0hOITp
iw4Ebbwq7wBgUPEOb8nzNmZ38ywAN1CdO4pGkiE+QtW4ythyC7gAU8XbhFUnb4SXkH7jieEnRNw2
R4rujG4+p+LPLLCUqlN2uh3utPIS4Gr0RVfUY/9pYvdBzxakLzI9Jq4+9RgUIm7Qb462R2RKzpJM
qYIYk4LsqPNsUKISKFrzCSS9WYozo89Ok9ja6iclWTPfCvK7PNlH0VH47CdqSvRfapN6GeA+ZRl1
ruRXu/RpyMdsUbSStz8WvmP+afdt4B43j6BkujRw1dLSNO85ncrokDxWW5LzVBZ24BQ3lbA9Jjv8
h4zetHNOHBUks2rNIVpElTA9SPx+acO3yFlp61zVOoD2nZ/ALMu2CtO/WoQ8VXd6zMZe+6Uaf49q
DzB5/NDJXJWoaJ/DCRHrqa4EEHQZw0eNs+ACCxbPswymvOPCB026fo61PaBvC3bnjcJhZ0WwY35I
ECy8Z+eAgarQ4e/dpRxluS1z5zD2dKo2dxaYhMFR+ZrpbJYFOhVldkys2IU+GTWfGa6uad99L6Z4
kfZwiPSTIru8PcSpqsRFqSO1SWpkhM6d8UjHl1xNNqoM3paYcetKjNfjZ2+H8o4PYb+I/jAzJGkU
UKePanyEgTrssaZcZeitLKyMqbwTPJqKvnHvABDebIDyDU4vbDp08OS1BjbMa8oQXgSub6U0wcuj
YZFyOYq5oOuOx58o+89bGdfvDiT+JAQIZOFHMv6098z5oCdorQQ5cRHnG5jp6IzE5uA+tM+YsVZt
jYuerfDmmv6O+x9ujo5Rs/rcvg4bNqX/lEUZPL00yV0wYxC/OPUlOGkAtJABN4Tc/WDo+Yh5hiDF
ofJIqs8QbNsELJHI80aaX0bDFVwJI0xUxC5PUUG3M2YnxUHML2rHPjdHeVuZYWllNuRlNhE3qVUQ
0hq9VdWyipKb3TdIHezYA5qahwfYsVYZYrVwAQQP/CYHXarHhRg0NjGlXH3k1HCxAddtJ97yMDmV
5OGfM8Yb8woRxq1n3OnsgEqBSehmE2YtyL/evMoYCS5z7Pb/o/2lnOvBicYZAW3jkoRL4N4JFIw1
B/Im64679dYnuuVC/KmRTQkue9R0oTrRVKGci7/AIuRYDvFeROJKo6oIxQ1RK0vzvzxEHWzc75vp
buOCxMiPKiVz6JmFF9DwZCINCEM0LVlzfgWu2JiS1+7CO2C87ML0gBH6abNqOm06uW5P83NLpT22
gzd5iMTs+eK0m8L9YatrQb1wZbryElFzkiHCLI81KktmZLlwnQ3s59ujSsObA9AJ5mIMwprdnskP
oNazZurz7c+pjM2et30Ktqak0H+eXND/TDoTupT+GtZJphqO6I7ug3NUT778Xp7wpUPiLXvWzgEv
UMEQ1kBRd0mwxskBD26Z6swSS3lsWIwCynKLSjRu6VQY/YpZhU1JWjjrmyZ+gygaYQxeW8cbO0jD
0BZUPuD79xvUu60wGdGS0ISdgyifNv0i73GbzgjIfF8Wge0FCk1X0/+bMNd31U/eZhMWcT0CO8TO
aTzpRAMvV+42QAsN19pA5bwUXrj2Oubk2WReTBT4E5qGXaVz/H6CFL3CoSCCPXwIDf+Jy/y6ptFM
0T1qujJAtjHPaMTWlSU/wCVM3XfhpxlNbLlUQTYYy9TNu53wmSe+pLu8HgS3NAdMiOApcGRQQZGd
4E7LMmGmHyvFtrkPPN02yWLu2cJ/Ls5ezQL7UQhP25iKHwm9/A3+NgHoHZYOtGojkypRuCn3UhJx
Z5fKxzFRmxNg7TgqLxGrvOZCrT1oO8GaSXp/O3Y4fx2GHzu9QYKNWGswABp71o4DkUcdQjNFZxBf
sjZOkCCipf3wUo61LmwZuonzBjdf9xA+mZC3H4Qrls0qG+JLmcbHJGJvqsRyjBiUBZ+t8ACmlunV
9EA3ha/a9IMax5JFTk3t5RXuIsQOIMKsCTXt5iqF9aqa5wPO0XflG/mSaI+M0KqOFZDWwxG6PcGh
kF/wWedxM+EY9k18KVAWn0Ww34FVTc/42iIWJxD53t2aU/IW9OZIYstWJqbQUoFoVfTcneW4Fsiy
W7x5LTOVAymVWWKf45AvmjNzh2/aVamv0xytcvmwkxIN5+clobEM4DENznF/xcjFMqqUszqIhDmc
91yIKCHMJU2/wX8UFjPE0JK8+eQkGA8y4cH17wQcabAkeEwcyvAHcHr2ktAB9N732WGqoJvourPH
FSPwHhZtlq53D9GbryPVEjGRZ8/9VKm7u7dokKEut1eNLfNyjeqKTkpTg4IbPrZGFjZc+NT33h4h
D9hbVpJfult0xiDMFvHwuFCenJvmV30N4RKAM1TuBEWfuRyxc0arJ2e2j3u9oOwc3onz0txkE8kk
jTSCFc4w3FRpZ2bAfFXk8NGDz8GokgkM6IGaxiVpGnSfgoC0jNN6Io4jypsW7IKeawBF6iklxkVL
6MqLewaQLOrWpsOroV4G6d4mTC7f8ChxGVQ57B0OJUHUfhc++UqKzCXIdQqSgglHPn/XuqyKP48Z
sQziQurF6qVb53RaEc46S80uCAh4VbOqz0q4VAgxHCdRNPNBsMbA/5O/y+UKkZEtdghTS017m5Ec
/OMG5x5j2JgmHb1LnmdYltgX2tmBukqstIZy/vAAMk24Ji5NiYom4aug8bDaDdYP6E8c4gKtHLgO
mYPdyjLruQl7qfaM2qmpdXNpJDG5xO/LJqS8trntdUpJDJXg/QrxQMMlHQveeZj6iCY9AIB4zIXc
wVDDQD9lnLCy2KHubqt8BfknOVcn3/+iiWCg7y2HG5FBLGoAc6zBXEB58/YI9o9UuUiGoPzbR+Tb
qGD/VcoZ6npXZ9xXYMwRsEY7CVv0EXnczi1aW7PhT9SwGQp1BwREdOn0Ut/l8EoO37hjFtpC6Cv0
yNAvxI+J1iR9PgjFfcb6e/v7/I1DrKtXbWosclXVgCdRcAgZufe5ypxFMLIkOZde0ETlFJZS/stJ
FgKoh9vWQf//SIiIujUGCCfdUa3L3CLdivkDAXSxq89jkjl8jDLpqxv0zJJdyBi2S/+UQE4z4hSU
i4F4Gz/dycruemmVXUXJcSwJbbbfoWq8tdXyw7hB9fVsbBoZOIz9ZYkP1GelsVDBuXglmpN/MuZp
B5j2XGKabtSGG2lbk0mgbke5UU7QkqTG1BEhqPTXaG7Sp7a747uXYxi4Nzyfh2+dCAT5nKFsdqE6
qZV+0Zsipf6g842qH6zEZsTn6s8mmKapoYWdZskd/XY6k4lW0J4Is6FH7gsP97cihVc7+Ug4eoSZ
NJLNVxWFqrzMMELXi9v0o9kxCvrekaWdoWtIvlEBgrASUStKQE/8lC7ElOTQFrTPF27cGMhYIDwl
eImZFCrR3wb0CcTB5oIR83j7pbSJF/JVZzcb37TDLEsm0ypuE7qY9/1CGfoq3PyTZ5xyQ9XSicnc
oVn8CXdsCckdwEIofEJBvvHAZ8rs5HmVdRa2uKQPlMjvzGutPyRjFy/8L4HLtjb0hSkx3mUMopHj
07s0ehnsxeplkBB7kMMQVJ88IDfbkC0yXjgQIn7xzp61fh4uPFi684XGAMSLYqdqmDNYlhssnikN
wRbQqBF3czEXIlQc8yAXQUFBjvEU+MVye/AEtAaepJCUmdQnMY7Zv03AIWme1OFDGnVteyfADRaJ
37Gqq6LIjgY+udYJ5RXkuOKMtoqkC35pHLOgn8ZMoglhVmA9lVnUDwgg9IsBrwKNtbUzWQ3aiDVf
4mwYhshoL7ewRGQapWYD8z2FGCWTe/FffedpTaYRgdts7YkVGLSbsAnsgIogYUGj5aLolLJePJ63
DUDPZQ0W5tlBEg6m0iY14xxt6hPLEewsATnygX2cQIQtR6VjX80GepirPjSDrseYQsJjvTb87Cmc
YmM4gLJsXAaXFT2BOWAn2XInKRYqs3miJ5V7lt1zZQig/wKhcEvUv4kt2+UPWbHdWpFTT1MA019X
4Nqc2TE4vNB2Xvw/L1Blf5U4k2mBD1erAW1CdkEGE4M8AYMre7Kn00pxAmOsE47L+L/A/kryAJkb
RJWDCnj+6SH1XNq6odrSX+tYM3HdqMcxit/RWB1rZQPgFoNaR/amKGyfWjw3w69T1U2zT9VQWnIM
v+H6Yc6/HhO3tmKRwg92L4NxoZmoAqaw6uw0mirGFKMx1vzF1AQ6bKrtILg73IpKSv2Sr4Lk1bMv
A/vlQSgbFdiniC03VmjTVpwzFBSlraxWK/Jy7vTHfdY1P/PgV7vlqCotKEJ+FmgeHG9BfGhZXXd2
+j7KCb0lHVs0FxRMvWJdoCBVMGF3p2qJWEYTZr2qqNHJul0dNz1DTsxYasbWnJRTSZMt/KDqK0R4
Uu1Pqz56lEoYL0DJBgV5+61r23I2bB9cvPTXmdPCGNrZYPShmgj7xF0ZkdNfhB9sDBHprm/vf7J1
WtBtNsyErrW7Abzq+mgotdjW5DPBN3PhW6Tb8NtlPzsMZVHACuxQwlrTHm5GAZyrq0ppXn6EEYvw
MbF6FnAFE8VBx4x8jUeS8eLge2mUGOxoOoHIF9Y9O7uJE18Va3mwapOCIW7beLu88SAKEUAHfQQQ
gTGs05Q83WC4EgAAaSpRjLgIeUZoCDd75uRUjadHdQJuFePooXi6mrAHYUf3fIM3JNrxbwZ8Dphw
xPirEnCLhHpRAgUb4FV1N8UsKa/shHgF8blwY3ifQOSq32quMG1adxlLIs+aQKrIAyDX233IV8hJ
jzX3C6i0eVPEas4WWmliy1hKeKHuPIDOs5eyei4ob7n9a8eszbsw30cG8IhFSCdb0s0mYwM13ZXN
pIEUu9zKfXB9RmAWzjQLQenOLrXG7cq0PK1Xs9UycpfxuHt4o/a+guu2Hr1oBhTYfKo+iN/s2bC+
vy+MSLUZ0cuH/VH++biR2F0OkAWV+vTHkerZ/E9kc3ufRafA91nklLm1rWi/qTFp05jac/AmUR6F
VdGMKX6haKl8+lv6PvmIPQTZXIR/BKm3KHAJctyZ2tucLREFo1UWmjdUvJ32NOS2f74e+J7wijRL
+lHh1lb7nYLlKGmjqHSOAT/ZeHPSQwCrYMmwgFsv0sL/dJDdbwh/PE9NBCVaqFWBQ0Y4bUoeBge9
5k7S0vPBRDSyqX6OeUYKdNLyYTGpHZBj6KmyZWqY4hzT757a8h3aH3s9ZLoLp8xF2nPcZzAaY3hW
WoqW4BVlT56gOvh4b610W6enqAn4MjDJ94BcL+zuALZbwuJzPNpWM16EQQbuooZ+7AtLg5Yyf87x
gyUnTKSGLNMqiqq2QemTKXJuyzwkClI+T6dLkEloVN+y/taLtUra445bYQ5IkhVcVuDtF1SiP8Uj
rFsOvihi1Zwjg3BtGSsFvl5OiwkRFNjgEvY4LpVKoPDSP6rkfgkFy2M5yoH+f/K8CJ1SGNdk9OJ8
RpS6w7wB8uxb3XQCHBnaVoBz36MTncmkD03DJyyHqy/uYtmjVMjgqJwNkn0XYkhvPwl58qVRZ/UN
lcwBc49JNNWZdV8f9JXGkdLub1Of33zFbYoPQCzPt8x2TmHUDnTAQ62MEg1eew1AH/VFnl+WK1Ym
r0VqVzWQ13OoT2UGQipJSJpSWbqDimmzkPcZYgUhRLWAWyPWmPQjDWqyh5mAc7010o83wgoLPn7N
YlsqzGimwKFvke7sor9qBmxvSUCQkqGbu92BWDugRKjof34Uozci7juo/O5CfGtJmbQEblq3PIz1
gFPbhfPXgzxSi2eFtlJ0i3//ThK46FupQj3XbW2rYubK4LKf+2XB33NNTHX9JLPJ1lMpgjF7rnsv
odpA+a+MmA43U0tzanAsL+XA4ubnZ1F8xPEFtSlLgJK7lh7HROH4LizdQwiEaYvpckniooihSKoe
7ZyPSBoNNyltjIP/uywzkwoEcZIeLdoOzK6Udvj72+CZWbYOK8a0NUE9CYR2PVjJIS6wOeoQ/B4L
XHWU8b2MGe9kPHFIBdkwiIgC+RAlNCJ6g+qcPdlNcvzwIjK2pKhPW7LKg4eFd2s2wHB0A+N4u+hd
TADXRU1Kitm4NVzvRhXp+Wly4OhZyNot2ySEIvXrY/8tu87rDAPLgwiHk4LYuPAkYcqSI23j+raE
bOfSBnanpJzRm//83ph8pvx5tlr9sZ+hP/L4OX8qACm91SOpiG0ur1PAb+RxTiy0PhR+RsAjqG0U
CK0XBtxdHbh+qwG8doTtrzM8N325JEqc4z2vmaiDEKaCIFloJ5B43LdtHvIHyGuRIXEzJxLZK/sN
ikTHUAf86nM7p1+2Y1hn8EobxYXZhWDfCEWkdSczCCx5Dc1gkeOJxPDR8hGZ2IQ0A1KQDTlmSdzG
Ie8HNbg4D1VOdFAwraRyGo/oit/lwNjOMuljM4Xqcrnai4h3Mhh76VTrLjQIGJqKoMUlMV5ByzLg
7ivx5bOQPBN0EwFrBi6qzxXM6ikUombe7GIlVDTYmHgClfZM96IlEtx7LYuKJFZwjlY6SQV09Olm
U5qO1rCPCuC2l5858BbZ/MdCj9LjHyfOKuMhYPLVjOLZrFDGD0Q0ADAC2bSBcno7hcBNsbCzkrCW
EzUSp5yM6ktIz42fWB3jYW9C1RCz+pjJZ2aLctFSXzUZFaWFRnD7usO0GGk1CUxSwJ3WBxKYL8xr
Cg72v7dQoGjCrCEwdYyIr0j1KeLF+EPvB+PfcSRUCQY+hrP0g8XyzwPoKdcM4Nesg9D5EURa9pQd
n1vQ1JZSdBr20vteGFqjUeaLlx9jmjafZO9pBlI6xj54bKzB4bW9ECBRPRRJhAN9cWg4lzneocrn
dUAhE9GfNjkPfMBE5VpOQ5Mm2WKIKIZeItCCvZbBgJ8nSaOFn7n85pfk+ULHyVLOSML+w044f7YQ
+bkHF9U2/fIFlMZcz/yTpGdJ0roUpU6q6z92Np3lSsxFcR26gyRT6+DHGOhj38Zo8JHgqFnF9lcV
R3Xm/z/hM0pV1N9AlE4r40GmO818SNBJhhi9Axn+swUYxuZNdzquG4keDpkiZqFMIQe5VNWHlxtB
6pCxfNrT5ZK9p6Z/KE587l3ej5X1W1xI+jGKNYwfVAV5zabk8xKQHVtvDyRmXVT/CjHg/ReISLd4
mJjdyd00uxAck7rQpqkyhAABmtStnjawSD/IaNXddwIOIN9w0Hk11PAwvHsethcabL9RxdRFQX86
lV5fZQ2b9S8xIads7+mVCuTkFSQvGCa87N2CF+ZkDYq5IxvEDMJ7ETqDtGl3WUsfh5WL8eIC15YT
fwq7k2ylVP0ewGjDVsnRk/L20n5Mm/4OpiBVmhDmieArS9EQ+Yi1qeDeJyy0UbtBPCRBp5lVgrbr
CzWl643Xb/ireigfuVcXA23JRqax3V4NtTJqE/qf+a1kaOB8BG9A2dxIRCjGu1SkN0/7WXmolC22
I2H+sxrxO0p8zCThTdC424ZkBvJWjTB2cheQ5YI3y9gJ1A8QqXFyKursKPk4aoWkaDc85esbRyHB
OHC1vzSOdx6Oe6d0B5Zm6bIaBtxmgA7+PyXywjVr3DrfkFOfD24iCkJMzR/UicnhGrgbgCgBtiHR
l80s1XP4URk2tsGOPJl4UxPCED1W1ujstAmNEDhp6+tSMG2CivsBi+oyRNiGnojtbg+kSLVo2g+b
F5uUes/xFm+qdJBpsMSOv4uJPA2yeKg6bv9UWfnL7LFgso8sPKmbJByhixpa3lIDObLiGQtSnybH
v/NwDcT3lXpLxt5gGmGUL1Dm46UfXLJQgdkohPqJcrvcN3R1o3Q2bDq2Jp5zPJ60RWt8lef1u6kk
kkNptUwRIio62MkkBQW6E9z/uipdqiCAiT4hBv/6a5wE6I3ADYyb2e83lwnkdKtUONcapWeAtRDt
hhRjd3lkNxxbXNTziBMADwkF29BS0bJrLED3oOBrlaB0ElT+EgFFbQcmtQWCwoerMTMoJGr2F8Pt
d92QA/GyZt9CsFc6u7nyJx2bhhvdO2ThVGrqi+My2Tqc9CPvUapZ5UCL/eG6RpLE7npCvsuOS+m0
f2Rdauq3r9wL9uz8KTljlT5Wc26z33jflLqDvmXkzy70mnRiB8Hxt6cJRSZUgN3NQ19P8e4DDkTz
9mZzFgtkjLlS+9l0JtmMvWs8Sw7s3ojvJnhfjxclGfpMq7OSCWMhzIJGglvg7Sk66NJl1UAfaO8M
zuayNfj6sKW/RYwAITgmnx1kHokZKjODCdxlQ7J0bDjRUdxT9pS7cQ8BxHDhC5gFDSPUSpkN1Lu2
H7KwVNF5GEfdy5RTF+2c3E9IhstR+K7YNe2bpvhPAzx+4Cb8gqEEK/dnAmgzkjjo3SQ90iV+F3Im
Sb8Ywy6OQoEf2BVfmMJDL7YT4o5MTQRWqqFUQ8KwMgyrtftZI5SVJLFt7QGxttMlAqed1C0fMBM8
wzGSf28fMCq8R/PIGoOEzoSg1Fgh735YBExlEdq4hKr/qPAgjDNTCKhvWCFLgAvgeNMulnNVYqO7
djz9AQrllRwhmSkJN2ruly/LPPfz07D1P0zpgI+43RrmHDUyjcf6PmO8jOVGg0lTSP/xf8o+ARrD
eioN8ZwM+egRn+rwwOEe7VUqW83Ir36b3+uKapYeWCXhRbLSi01C6fnsfXlZdNtxwTSqphlCULYL
vmmfCM6Ypx35+ybUJBX8dMrm4bMLJFAD9Q3kv2IzPEutel7xrozqqThEgmqsPfLLw6KQ+1u0zLsE
Og6/aTOjraSAyWn855Gz9+Vj3C1b8hoQuHYlIFYbCeEyT8yozEd/AfV53eNET/i0GC1fVzCShY5H
Wu0hCSL6tATtATLb16L9HhOJVLjzNuPY030TC7qfJSAKdRNaCdYsXThpIfM2p9QaXSECOZ8wcL5J
Gg/uuLPBglkZemUmdE+7qSPC9Q+M+BDK84DwFkvbWuD+NnxY06SPP8HACUkqgrIpEjNeeFzbgvw/
eAJwE57zdYbwjorwoaqeY12cyTAs1WLjlICnB4HlsNbRstgZefPBVseNttraxZN/Bw1cQCOvd90a
g49X6Llerg0kaprsKfs2mC+uM+md5pIznP7NpDYtv576WWSAAjZ6kHs+vSTKI2r+9dCMEy7hPwZU
2RjP83GVFVpy4/Ihn2eFbGr3V+VVYBlDPcGO4edQ5wWe+MdIU9GP0fHxCpUcjiSz1GANsgr/QPRG
aJjGiRvitxNyAW62n8ueaWf+bnoexoMDzoUNJrpa7ANKS475nVs/nX1FfRg2+dG6wxUsC+oWRu8S
ai3tu5oAsIAwQjoIG/qVGbLfmb/l3ojXK675H+mqFZubWKZtQ4kHHiRVs+5/Mw+e98mCupCN2YLY
+M+Cc1wl7UcL2yzvSHtztXMHlWNCthvI3nzW4T9/vzdKCAxHWNImWes8PKZPvp7vEVSIe9meQkFN
Ln5BdHpU94fsTt4X7Y8Rud4f44uU2orNm2IHep442Ot8HIeMxysGq/9PSfc9FI6SCDtM/IuV4PsF
kORHfMoeST5Y/oIEISFBD5yV7u90aDvlv003hy4aaNFPGlOHK1EA3wwkzRMcjRTdWWFliN9xeKLn
b6gLct4+370h2xQN1Rq878AQuQybohG8ndSp/zASy+CmxxJKwFz982grE4vCmY8MoS8bBtosXJ+k
474nCTCsG9WzMNySjPA7Pfd1K6TKgiDL/pDryAYOWT0zmtr7EsfcuEGi+AJx8Lkebasx6DCja+XB
1TDfUNBDbnIbh0pqG6N9otyg5bbu1pqkVxiDKmrs0P2BOruTYuTt/LtrQOvtOL1PbzUlOoNOqpj6
oFOGW7rMt5HfhgyeHMXj7n8XImUJM6pgTBxZCTtS002aZlwYCfAGZU52wd4unHmXtpxm4asPl/3c
iQaGOfkCaYbg/tFl0f8JXxU2CXUtfxNwrZPZK1cuOKerLnvRuXH60ou+0DRe144WEItTBkslmTA3
OMrl7k/2I2jSXtE4/hR9JlLJ23fHwQMHG/MaVvkycfq1m3bIe+xk09pC85vpymQgNXZDyhbKU8/W
4fF2RwE2YRLwew1HNb/6Ra+vZRJ3QCHKe/tOWuwrF9lKD7XenohY3dM14RJ+tmVpjP7Meh7FjDlm
s0jGeNEWOU/93PMCs9EbcdYiH6RFFZQerYiGbWNvDim8DtW27tk+zY43UwhwvLrZruSITD9EJJG3
OHHDPggN6vtL5OkSwCeYSLu2CUzLfpKeRGjT4HBLBeuvJUNlLDrjJvVyqCWXxLRIb0YWEF7GRjF2
bdEGjHGgY54Am26UbabcQLK+5boKYpdkmflf35JlvOQW1joMscPH+3fI21OyVLcZ64Em6/OW5XXX
kcf3JjxnKF3py4iMAICDcTcMgDjbAOP6FDYtCmR8201RsGgVP+9PC0MTulPT/MR7oWXSbAc9uDXq
fmFknR4fVHvuxiU199bscF4/cJn6tznPmTNUyxQNNZvoSl2vcWCk71WNA4rT4xYm7+M/JgMdbajE
z7pBAio4j+/mJHKH2u5beYEK6Cv0kO+iVT3j6Tzk6MO6nrK+FQPSDDCANNYcQZggl4eyEf7uwnQZ
mYKHGYhOmVwVrVl2lJdhSpMiUVvsalaLuRzWge2qcKZFNay3elkemUpO0yQeA2rTBRNBpLj3pC4B
/af/+Q2tmASuO9tj1qftMy6PkY2i3kRKRK/Vaceus1Tz+kTEfzu0I5otgrhVzsfxQ4k2EWrwyf//
qPf7480nxndQ7M1LcDAmqVV8nCSUtj6x/TwIE38Wmhw6mfYlih6IOnme1khR1Hea62xMFYxzwQUq
X6oyILJwqL72BqtJPyTAZNw1CSncK4xs7vENFZYb3o6jidvaePKTfDPtMDOFw9D8RcrXm8QpVtq5
0c+5qNpv46GpM3k5WtrtHJkXvZpI9VFYX8X5oX3Ehom+7dxv+UInrmnPmuzw07Sxbfc8U7R+VjAe
/yU9z5B0NZTLgmJBUtOp2vOfcr0+UZYOVnJbJI4xMiNk2HKtFrMHKnbs43PJ+m19u9GaE+xs6tEA
xga8BguoBjLAAY4rqSofQtsK2sfZkDhRRRhvSTEaEZmXxOEmz/XuRWo/tp54rqV0OUByO0exoaCm
WC0Ub4NZ4ddk2P7nYUHBeWRoiEBmZDS62XzfNXO2vme9M9jb2RhbR+LOW8t8Lxb46J4k9Ulv7etM
lM42Cx5b0zURXSPUb+LPA6aomS97AhM5OFE5QZf5d+YNd77F4dGQaeGWb6X8pN8RqqxQvcYIGqa8
ft3iEIDOaN5bkpoUVV37Ok/bsrjs3+9jM2yXRB4b69V7xAxb977trHZmVLd1Xy1Pfk+17HDCP2B0
MRda86Sxw/Br4GQwz9rammtlccKgl6wTWG5qu9H6hO1u1rJJ88c7WKnFZA4GFXYlgVTyBg4Y++Qh
l3Zs50Vv9mkKIQjlBr7AdEoG2n2yFb0t8jbqF3O06AfBzCHFocmaoQJcTXhkQNkWftfVkpiyIPSJ
Nx1p6y01uq8Mk/Bewvvuk8k/WUt4/w8HkejQjWZ4DpZpwllYK70xaEkOq7fovBGfWNggEVbpihdx
vJrbgo5bFhdUB1q64FY/pJS5I37LrFY6JaIFH31Brrv+IzlPOSvuZ6/gohjQNLMyvGbLXduXAnmV
B+N4bGNMNTxaoa5HO+qCJ8442axDnhSrnAjdUwaaug5xXJ3kXIrRYbuSFbaUUE8QX2YaPm7KMnys
t29jABrFMOV4tzS3znvwrWa1fjibqf7zKHRsQBx1PfbetnJUR2gsDStOqyGhKO92Yd5YcHPxg3Hk
l3UrVaWJp8B1CY75vzOLNAhpmLjs7zKdXarfp8XekuLQL74P2zm7oKouwIo6tQf+IC0+Cd58uFWR
YrWJsocStKC2qYHHRtUKtbf/qDX1mc3ct5g57nhY9Ll+LGcRoaesFpAdBKRliNBJNmwc/nfZziN3
epj3igiC3Bo6N0ltn9hUBcZTfsOuZfxb6TWCxtC7C9sEHZI0i2yGvyylwgwWC5f8Cb4lLBjgMuAX
Pa9fKRb/RlOyjNw3oelB4twPU50WhaT74YZEPn+5yXrTVzi7Ar/Y0fAhFsFR93SBvY2Zv164k8HC
fldWz71GzK42O6+/dhkLrPh3gtJrmVqcFKj2fU2CBGEk8DEkEY5Dj2hliJPKLKolNNP2usGmoOcj
qQyajnD3Q7mi/isiN/GbwXUIiTKlN+q6a40iR3iJOHrw30j84H8dsbXnVX4h8qlJgRHYtg0ZEfcQ
HxfPlE0qFCm100bg2+vO9KpsgHWiQ7MhY/cyB5iM2KZ1bxETT6MocvABUiOzsbJLjZH3Rxs4ajwf
5rdsO2I/5Zn9ExiUF64IbthO759rwF12iCCScID6bmJru5/K3+KjCRN4csLEF51dBleoC2f3h56+
3Dx84eVLPLw3cm24cHHS7thlzRMay2ABsJxYviQGp6vCB2KSpVP9T+UE7xcJAJjbzrL6u4G8Wxyz
RnEjVN3s/g9sKxDHgu5TT/9vfPNmNdLvFAWKbCDKyqs+g5H6nJQmBFKIv5TyN387Jlq6XAHEpdZI
N6r54+MuWVr4R04EFuM76ryILNCYQzVVeXMj9WTLgwY4wSzdDqEyuVlCQRRxiayA+iw6qvogX4Qh
tNn1JlxVSYfYWlSrFd7SRkpfdv/A6+liiwLFoZCsEN03ToolQM6VITVHGufvqE11iC9uE+ca0OzY
t1g234+p6P/suD3aFBSu1fVb4JSIprP93EU/SoL0jtW96JvM9KfNr1bZHtEHzXPx1CrvOQedP38u
TPSBytOwcMHjafU0/hRGr554/0msNT46xg9q5CfA41KEdkJdtPRFMcF+OMWI6g0OYoZc4tJEcgbi
KPD/9jeuyQ/2cCNDkGIUQGwXw6Q3em0tH5jGn/EofdnFty+aqWPXnkKUaloQCNdqdvKc31X08XeA
SN9xQOzVi6TvwbKUU6mHgHOUHnl66lvoSS4cZCxF3CzFVWZ6CGP9qFSAfufSuq5s7+9Yv4+jqu4g
9pFlppTcWI4si1z3IooGyWZLNCMQwqPmVl9RkYuU5DRkAxG+gr3icE+B/X0HIMuwJOJ2V29/uNp7
HfdkJeMF9OYA5Hw1GCsclgKTCkFDQd/KTg+G01w5vuIgosyDgpfgraM1Icb94aukBz6vMB93iwSA
fAgfk7qWnVCGoN1qooztwrqaT5CYNttO9Zw0iuBJydYXXfmqQ0fUxmbvbJWP6Tw5pjcw6eH4/KEw
FuSgM/w13hNN2CEOwJSto3/v67wairIXDmM7MzSkngHspqvkD07/okE7bqSn+t4jSMddpbJbe8u8
5SepUfaKK+5TbWLdJKpr2vR8SPPPl94ARRcGmT7JJDQpBkRIv0LGbP0QFCYmDdmyq9NRE1eNRFRL
HlHHS55MI92rwnQdCKA7iib+uKh11nrYNqtlxI3eUyFS3uF3PE7XVZ7HHm2ru5lz1u7VCmhP1jEl
F+a4Q84iTik8VErA91KuV11nx4LTL2/fPQlBwOGmSy2C/hGrMMrcIch21mgzmGxK9J5m4RAoYOId
Eax4Jhd0xihbO3RHI8a3lz7WHzfdO+SrsX8BNlDQb/rGSl1lHB3nZI07MgbKrPusmbvN09qHMYIt
sztFN4mr+P6A2J4RJLmBjGLmzP/xVyyoHk8DpvDQKSOgkLiumoX5rkuFQT11DPZHE3TnaPQbQ99g
UkRynyyeFRHFB7c/CtoMpIdUQCGpUBDOM82ov/Cz5U7eAL3MXAp9QoCjOfP7i1LD057RjdUo4PsE
/R5pVW67esKDEy76RcTZl5T3O48JkW0G+F/mtQtv9bN/biGhF760HMeIohguM1DVKtaN5BTvUFtp
AdrlX2AtUd9lnzNTTX5FbAySal18CqYK0lLPd33rK95iNRI4B0KCTRMUFZyNEJhD53id01cv/GP8
AlgbxIqTj9tq7xoaqnQ/onK7b4m3qv2pZ/V4QATutwDiEwHyd4NAZ5AI9aLC80TH1HoVEJ/VAM5T
bptfbXtPRsUHVEy1qJ8PO1s3WqIO5BS+jklri/att5gPqV03wLuX2XRuYmr0HCWAV3cczOssDR9M
n9TQZFjOkX+t+6nx+Sih/WLwXtnQGO7a2rONLUk5yG4+cXxojQfT+ui1/fAMtPiFzQ0zeOWtpuek
latDIjqL9DdwAVLsRD8MFx/gphYKMOhtDHAKoSMfB27TYGeSKf50wAwKr71QN1eJFBRgCcsJRTKj
8WkAXIC+gZep8Lrjl7DdhOZpqTrTUQje20KFeTRBvoThyvGkHdsM7dOT/+2zq8d8+ihswWDoKz1w
GpR4HdRqye8zSW6EeZ3abFXN5g8fjyOd3jVg4xNRuPPesaSVbD7QE5OtPy8qpL0EYg1pgNij9EmJ
cI7w042fMPgdKEFhiZDLYsEV3pxm1vDqvjYEGN/DPPrfeIspbu302KL5CIlLapNhw9HbHQPVXnSk
IBxc9pHeMWQW/VUjUYmwXGecAqo7PwRohl63BwlUIW0y1Dk9tTBKJ2KFDXjEgY40K4XAJuhrFgdr
nwiBKqHKZz1ImAdQQv/dawJo7xQs0KLBR711gVGZbrbGnzIOey3i1oQ1ICG4MUX7L5OfEEdO35XS
ESwqZo9Cc2d4C9uvm5RlQSzbPMkNubGIIGRwxprImBKA6OtI50bWxIerhBy+iLV+VIwDuVqx0Oc4
35Z5g1C3bm2TF2HwJLkV+MbO+kCZ9VQDuUAUiX3uZTzH1pfh80tAqpWwkZO6j+gUa+ttCxY3epAN
PH3iZexFWgD9ejwhQx9cwvC6f6pA+lDzsLvxkD4PX7p64PqgZkjrTHo5DXGvDLByum/uKl87HjDq
PSr0MpZ9ktI7QJqoWKBQDJUGUkbafyarG6tAp3H/qjWreiFMn+1eydugxV2ooo9lQ7VDjT127E6P
3RStqpvP3N7nWz8twYlGR9LPE1p58MkN6Y3UjMR51hlejfEmjn9S9/dQNlowSQ+9uRGNLBhaJ4BM
lD4D7KICyloReMV3bn0UJFWmzT3L9SbIFHRIuJKyB8ptLCHF1cI4hgFtWzrMTKCNTH8XBInIRMIk
B5vpGQHM/pHCDy7EAW9cknQQ+ELSQhUYB+4h98avHPZ/IUD73fkurFEYuYhGM7kCu+PJlst2UzF1
/irpcibhBzEbnEqqXaAxNuHoJZ/BjehJb23sDT5kLpFkOyUOHosyl5/xX5DDMEyh3uP5QAN93x5a
Q0lGrTrVogf+Uihpm13IsaXfSBiPJ+R50YMJmykYBsuTelkA2HHuU+wDehwrJ0iWxBtgZxG8B2af
Ym3J7l9tMx5i5BVvW38AddBwErLo2M0fvyeqZuTCoYiGIZZ7KCP0iGeKA6WEVtnA1/rBNHF958xU
/7qvnK/UPXqgJN5PtaM93DYEXG+IEDqdAqY3FgGIFy5GX9eg+2SjtkmcS3VK6r3BqSs0KmqIuYo3
1uv2bS7rHi16658ndlfawBFODpdLRF/FavhG9QVbY7bkEYp7QIW23JH6jp91BaXbeRonAo1R5Sc9
BDlys4yG41J/O8p1rJ3SDeEutaPHn2X1WehOzEfRobxBo0q2nM1oISAuhOjiMrttXGxFSzZd5FkE
cQPKc/fdVbJ9aN2S5/Xx4to2+wL0vhnMuD7F+4rwLQVNIx5t/w4APP+0LJ0rqcIwlxWtrLSpcHcb
I850tpi8QgiQaxXWZB5EpY/8ePL7zU/mP17hJ+28iS9BLMdIpKxUY31/Xu6LrlnFPDk/fCE+/Dcw
V/9ANyCQXqNwAUFYlytKv/z8HkPTf8bIJ8X93dfP67hgCXGYU2MIspO2/R9MxiQmo/EV7U+Uixyh
x0NO85lKIn9+Xjz5XZ8t2kKGZRzlM+kPSx1/a8S5BeH8wrt4U7wgNb/lu/9YW2cX6v4y2Tmjy0ny
JPhsXxdoYDuYsLtVsSmvSkTy59vPuZZl8z/YJ7s+DUoImYMRM6Aj8GUuWS4ZZqKGmTfUqJwfoLEd
hugEOSecyXC2cxekqLE222hJ2EsC7Ov6t0tX9LBj8T6qQDrBE5Xz7coTQKvV1CFOwk2hwgchPTvo
2geiWK0zB5T+CEmWVYm7o+CbAyWE2wJr/174a0Ry2z3y6N/IXCiofEZvnWFohlLbY3oBVWDFU2Ra
dvNEocKGNqFHIIVk0+ZVZ//gqXNFu2ywZs5OC1YxH15a7NQyizNfuv5sSrTWE03craGpADHl7Xru
wUeG1AyY/NHBIO8W0m52nGmc8Id4xbfSq8w6y6ZdEPNO5VlXCUUWP+Svw2FiP2Mtwhd/Gbebxmks
bomIc4k+sEeoJzw1vmh5mrt6iLlkPSKY568r/pxX9DoljnkZ9L3QbGMB6xZX0g+8c6i8diFs0MO8
OfMQnuwy7Rqb/xlXysMuUxH8CGtPLhVmWUU6c5pUPdBFKFRWyX8nAi1wLJRcAuHSkWAu8YoqdBsY
l6g6nC89ZqpfHEJzPSKNaLU4GsqiHiJpz4s+uBtMP3PhKsIS3EkaWPI/Wp0Pa4q43fgbOQ1TR+3f
xWhd1Wzo4q+Y/kvQKFKB2KHEF2ELXwXD4Ag1+Osn9B60/N31fNvBDdfvmR34BgYIhNtCfHm+lGK5
XpAS0xisD75rLw4tXGCwfZtYCz/Hv602D9T38oQA6vTj7cGt+zau/fFMvEYWRNvmejFuQOLV3Dug
JfyGWKFsng5FaxeZZ81QnMHNARVZDGFoxa+xDbtow2CZWSXXRFBBTDPaYx1O2BYBi2eoRoNqwQMu
vvEYGn1gfLt2/p+AzGS87M0J9HYun2wOyIe8oZ08Q4SeOTFkE+0jIqTJ9UBZnvmafxa/yEUa0OSh
z3eMM0o6LCAJl5VeRC3R8WvmkJUfE6zrmMzmMxKjYeo6SIzjeJKs1iTco7nLaP3QwgDsxhCUdKws
mx6zsfAHrN+T2HdMAiY4kBhwW1X/RSSZeD6Lq31bmyc905govijFKS7wH2DwJJCwv8MJTZoOjujD
JjSTUVV3ZQ7ntBv/x0aVWnqlw3SWUoEqn2w1aU1VAR4yyWBaiOxm20PrO+w7uNU3uhYNE3f51jVn
bQ8AOJJ0uX0xJG7S54FyB94OTWNfl86iNF5uR9Hkh2ClMEb1SYKQROumiCPpIlSJemV7M8r5/yLN
mNU55QtpSRAyBBBcjxben7jv5QI71DAyS3gzIm7aEVkhyyQUuEuAnvX0rut/zTGThpVyJhP+v1Sy
eSxWJ06t21bVoqSRuv0lLYtD1I+MwSB/2aNOnLkz+M1tE53lxAZ8//Az936vBoRWajG8cBQE87Id
k2Uz8HwsXB8lDEgnZTeXPMhHi+5T69SWZc1ZW6aMf/+fC7hF9iiZglLpokjsLnfBIfFo3C9bNT/y
OaMLp6gHbm2WO8FwNqPcTCT5VL6ns75sPRWuQYmAkeoWzH4SnZQ5wRtwGqajrlumUhbe3ccqG9ks
tGME3XDstYYRUCtBrS9OaaUHM7DdlxCbu7b3OqBmkWWZf+AcrSpp7FibalQ4dzwdsu73LI/YIpp7
yQ1FwoZ6CYqFva+x5GzIVohKlYYezuPwunPau74uOA+f8sFl33//oDjFia2MLHzw+4d2I+mdc4V8
BbRVKTAcFTpkd57p7yk4mht0yxka4BmXxKE21zoByMLELZaJMBbzTxXcWL+jCY5BU4AUj3bqzzJx
7iPLWs5EaxZwsmssdh1SqdidfPLsJpeJdVNtFuUbb96SijFbJbbzk9X6M+ynu3+isSbVLpS/XQrs
FKAl9d0+DxZAYanYKona4rMgDz0SFJBv2aujTvJnP/cT/Ztly1CxFgp0KpadAiqPXgbjxq6zVup4
+/jddYtUhD58lXEmNODXik8NV5HlhvTzDe157d1s6j7w+CfFV3Xn2BYVfrkSw0LNYydvgFUBziRP
u0DwryzcyTRo9VmksHcnPv8J36Hx7b+3ylsQwFvW1f/jKsxHjW7WxJdKv7oxkK3n+EBbIT0+iHO8
Ig5FdBGXuesU1TmSRsw2ZWm7cHlAc7ei9GW8bjX/0ksHre1SWSTlQN6vhnkf5BaRVw0ttgiqz61s
7K6fJAUSXiywtrDGy4XzZE5p86pauA3yQ3T8yAAtbMxDo0a29iGx/HqV0391vuNwohuwE1OuiV4n
5ai1T6/3oPIELRS5GVShNptq32KtJPYp7mRdsO/w7JBXbMZNBgj2k3ZIYzd78UMpPEeRPm7k1dlO
IMvFeTb6FLIdsUZetV4evMX4YVt7H2oXEARI0t+rRHLLBatUF3cUA5qXcot1vfpNHkUZXIQm2ftL
g2PhZ6J0wSqblx6I2GGujVmt5YzjBllIyH1jxWXZnNQ9D8a8SiYZasU5tBVcXSQ4VzWYVmYPaAYX
Cu65c2cSmeVKOxllKjqop6TmjIohJDlxJD2IbT2vik0fVn0AzB0EnJiQrcDDYxm58B+y9QqB+tLl
2Js3j7lonkJtcPm1UP76l+D8XdmHdhTbxszyoJKHM/QrF238yEUhaNQsfJDi3SQrrnlqZRPZttif
PpSfue8mRBgBqcoRpmHUD7JsYe6ue2O2OBxxo2irQkaC5CXm8UU9SMDWbfXKIOuWbYJmpQFjWKf2
6usBYHtwjduU7EjEpHSksGBqjJpYG2idwUYbSVcCy2Df+iU6wUHR7+wCqaMI1lQXkTNmOvaITbp/
tavG68RFTL79eRD9DB0QYkn6RIvaKBpM5mGTJiq18o/RXv3Db0yN24VPNreEYGkjB+IZX5f7Awna
o48X+lxlfjWN2hmrAO2RnKvy3NJGddGVM/FViolqaFD2iXdxakeAVa4xCmHhP0NRIEWNqp9vCuWU
n+cEErAtMOODz8qVGaGA2MZtiPREmqWd2hckLBeyLBHOkCOXOEtLfuTcOrCiyXUBmZvseZLbGHJq
dLWVQYfGI8m0YKCmUJfGFHQeeI+Rlc6HtrRg5EhIjlJundxhJSN4Gvj7l7CPdFI9McsPBRUzekJ3
efTd254JObVTQKGimu1Ez5x5FEwiEjEgJFu3UzmBhkoWhOkIDYm+bijohyqnYhh0IcEdQ4CzZfuw
0wqE+keWa8sNFVUSpA2HIstZoZAfxCIpKISWr0Gpg4oQuiZvP1CFqcJwhPoTsWYFMlPBNm7gvfOb
H/+3aM1/1cp7pUxR29sVirAsMcYOvfczuUayRKVVRx+NZh3Tf0hVvlSuCljWFrAgmFrc3h/Fe0Hq
722jnqByQguBE/cUAIQd/5DVQWN6zAdiH28nwa8+X4buu92h4yaHDMtIz7A5YhIME0i9PVeZLOi9
z1brGhhTNZOQWhl97yF1/5JX9j7VZfYz61MzsdNpwH5ThvEXaCrxKiwG0YlwI18wGXqoQ1l6GKYx
GpYRnNpRz1nq1Hrx3ZStfDtjrC89JmeCjC8Mnx8hjBoJ5kee0d3hHoBqQYu1sio/AtWXWKwwFJjf
B0FOmJwqsgsHAiKoBWO9PKEjb4Fibl2X9BmX9BPHRShJfkP3iwPXD8x4CJ3mb5n86/LZN/EaqB6A
uRYIPChW0jy5FuIjPotv0rmjfH5W229dkIJELJ2OO+3SY7M8O4qzp2AEmFSZ0N8Z7HU3V7fUXAiL
rWee18sS8ZFssd/jUfyEd+YBHupZDeROIPqbryhSeK6YLcTFigLw/IfAB6odqXT17TGOzu5ZiYpE
wfGXwxjzrn1S8/UaAH0FlTV+3ICX6rXGJnhljjn2ecLqpTK7unm38Ih8srtcUOhnGFRBscoDENrX
ekaunIrDx8Mf4qHrq/UQawRu74CCVbaLwMVRcQv7LN5zhj0vvDIr9xGLvBpTjm8M1UQqW9bQWCgt
p8i44I0AcsJ8/xfFZ+vyIQlOQ/074oaJyFFID64ZNA5HGoo2de/aCN2TsXCMLalVqC7sYhRKmOwT
XG9iY6nOuMBnLW9c2pPS+Bky4GZlw4VERBahBSTDIfH6sqoTF5b+LW/+71VNMVa8CawdOc8ot5np
AgLbaBGM2uTHM6wvdpG8nni2lWap60POZ9dzFlvJvv5t9FAJ7AbKVI5l+hKnQF7oD+OabeqYmUn4
MFzRAG64RUqojG6bUzi61btXgMfHVv9F3eck03/p2Pprzu1PqbdThYRmfieZNfAgQmYe6fk1JlVC
alIEmf6k++TmutOFhH2xnu4mV/7LtHUlM0X/kV8l+LpT4+jmBFHeYWJ3KZGxTdEy1hTbNj1Dlg/H
IeRp4JQZLh1yho9EqOBCcyoOkO5LtdEgQUy+Ufu23gK1Nm3dT31sZPHeFEAdvoEqgTtV/u+NSZhX
cUkKcMUTYRXdpjfq8kDkIWV+jv2MGqVpRc2RtqGoU2mh5EYXxpk2Emcc3f6+YF2TyJv/MvjBkjgy
RzF8Nli/9b8BkNp7Wrbykpa9p1cNQwd43o4vf904OC4caC/2DGBllHYLce8F4d3Zayr9oG+6RDaV
inBs4dxaSApuwly/hqItJ6KsGV2RbBiiqVUpClaxTXXZ3OY4OlP/KcI/dzL1lVLrrN/1hzrFj1za
I6d5eWHLTOacbq305LvIzFiGeLKAE41ycyTYvq+rGOq3MDhvCbHgTerZ/rld8DtHtKR05wkJWmGW
2Lr5430E6ptgS0yFKGQkLEhoJZISsqp+wJfv9f1gkdrPcRyOlYTZTrJDq98dGLMle5k1otZ4F2PJ
+LBLhr/Vmag2NdxYvyAA8GFruCqjaPyG9SXCBwVjOsdDvNjzx785t3C2uxTJ4uu2gz/a5BIlh1ap
mJrJQ9u/ZMsdFxC1z/HswLmaPN8gqUhTwgG2NRP6kJ3A6aBWZ94TVjc2JsYRMDN8GzkXc9nC085U
EULteaK2/jSrd6eyByIo9h5G5rRTo/s+YsDNijxrPveJ341oF/1R5axcLZg2CFcCj0lU81nnM0EF
qHRCA/tDKoeXwWmZ8UrOS0/rgzoLH/CEpYCopUyXL5wMnWvYPWjkHNJIjCqXHrHV6vJ4NwjH67bM
dr3S8pep/Hs28q8MZWkBRQFU3Yfmm47rAcx7HHs2wrWIOdeEaUqDKqySnsUSzI3ZZpSyVJSF0vc0
IiGWlcamU8gWkgFN4au/eYj2Qzj6irlci20r9mfJ+pipUZ+A8CVWBNiQL8cJJ2cbNMWXhW5CP6kX
lLiSzsx6zSOaVPkoX/HXdrgogz84QzrI8dR0aqRpz4HPKdRVlHL8/bM9uxpjaeCsq9P2DhbebAQz
V7Ry4SUWh6bKGdT5bYeTI3nVX6p4ZIn3hh6V8qeXBpk47AvuDl0CbdPaiy9tRff7QvbDCwdv84sm
jt3lM0hYWflJOfhAS6Eqckggoe9eYet4K7I6sq7TM+Co5UEYv658zDvKq7ddxfKTcjOsq5lD1iIh
ZFP0ocPgL1H6VRL/sRlaPr/D3rjHIGu608q5fg4V4HvI9BBl4sppfbCOnnTS6s6V1TIfBfnlHqjG
+CBrkR7n8kN+FDaLwa0nUGJF6ErN08uvO2O6aEwBfYRegoVVW5pigZi5b1wzzzipdNyEw0QTpzA/
lPX9iPseUms4KVAjKLVs1k58K2NKFKp7UifMvJKeSnaQKWVefoPu8uu9ULYKdzPjgPsLY/FKmbQY
JsgBzZY8GrbJsZkgwmxsKJoPNvL0AUmVm5nuottj16x1aazC8BzkpfhuZJBt/w2ES18TPdvGA1+P
I+2qmzNTWQJxvug8qg90EcYCjOUidXs9A6Qs0Tf6Hi5CWwsDrtmZP2MX5ZxDQP3De46YMTUGnKPP
8uPIKo2PYi9YDtVvbVa+e2In2ocXFzVi0C5YS0vz280kAHWAKRGSH2WhH6fwGvYBlbZES/rwi56V
We3u3yWbQG8NpFT0RuPf0r6SRDpQeyy+s/1xKCr1/w7wTAc0bDGb7yJi7xZyCKRwXM7Sl1vBH6kg
0M+/818HMCwmbXo/EAZ1N6hixLyaHvwm1W719W11uAH4noYB1llUNE11nwWR0Kp0Tgvgu4/Hwoa+
5dt3ZVDX6UMReieksr5IGz8UfjCgOSFD6nOh3LgXVVBlquF049Tvtn78dQGPHM20ShqK9sH/IH0q
pM4KxBz7fpozFLXuUNPwZMMCSkQFkk04yNzZkNvLnRFYpbsQwQQzMuIGxnpW6XSd2UaxzdA+w4FS
2EXQwAy5YwzmrRtoqdVTs7pqyGyOu+pWAh8sREcWlDNED0R0snGIJdsWv+7KsspIMNiJ8dWx3NKW
fjpMDkNbaJSOnO4cQUooJaaVEGPjOxv3fQbQ4KkoacG2QwJswZFqDYhsy/lH5T/Getlwhadbl0lc
EUkmeme2Q7Qrgr5Gfc2appEfU3A5B+jDW2t0BNZ4vetbep6op9Ft7Stj4kWNVK1EbLWSCrIbsawD
6L52eCa1eNOcaJqoXO0DT25WGlHZboCFR3WxcSi/lNiJGEevGBqeyoaQQomRmlrUaoRMRHo+awBo
TT2eqX4SPDfcvmBM0o7AimlP8xR7h3H+4YKikiIs6qDTYPwLFAP7cqLlhUPkeHF59Eo/KXhApj4S
7j2RblCwGd53RdTS/5FkENpabeyv3lzRgqIimy5fa5/mQoYMa/SArwbf8DifabNgCsCRV+wfzQw0
Vuh0MBoQUZdOJWA70uDBsHcirapHoRadChKdowTWAOcKbPthWQTDpQJNornRWMImphX9r0UZ2Cl7
E62Ef6Ihk3I0caBoX5Ldp0cNZQoZRpyYj+zKCu1ZGvahhCvZj0mmYLnlFIR1o26ahYB9JgA55t+O
21FOS2fzy80paMGnekDyEvt2DlrXqLwF/VNRTocfsyuB3DACQmt+ah2TQ2WqDhxoJiFJb15ukaAP
0L5HcfrUggOcjqId7jSpXZi9UzToxPlL6BhAFNT0t0+qZQq5vYRGKLFbBHxQFNS+mu27kesF9pv8
OIJ8SqwpcX69c2b9PMxyVtzziAc2Vy+wBvNS5jC4uDNJmpMQzvBRb2cfzwXWfBIL2U5J5O1I6dzI
0sweOZwQHYnRJytvwLKeenV94ECEGa4qboLjgrG+jgcJJ/Vsyzzzk3nLbPKTNUYMEUSkFquJbqC4
0l5pJU8q/utfgIShuv2OxefNk/VmI6C8hWcJeSfekt2IVJCY/A8Rm0othG3HGtbj6q/WZWM/QLtr
2VwYuH5wNBLLyjssVnrDlw7UY8Bb1pgvcc9dkuYr+Ght+gVzTpCzcHLlMEaNe1dm4ONoFQ+H19RD
ta1cf1CBYlLM9H3+zkw+2DVoxf3NJOfz5OFrkxZk7PqzC0awBKJtQQW2OMhNeSei3bKLvi22uADN
fpwMGLLsgYIMh+oKuuVAwzRY3vWcxJKTMzLrqnwl8u6H2X7+anHbDpH1S3wsRv033DsyGfeeQtas
dw/AIY7p6pwIIRAkBfAzFcXR7NJSjMxLO29bUqepOjjSD3gxBtXFIHvNeT2T9rhmA14ZLcFwaYOa
dQn5JiSHNXYNw9/qkd77cnR8W7nZY2oMRH5b7QxrqPnVc5xO9YODZdSMLbfmD3qwiXU3n0kFsNvz
LRIfFwlsvWFVXGTeHhb8ws303koMHZJ/LwZBV5tveQNsXBZJ4+8rc5vp0cbTQJpZaVwozne7/AXr
QfSEQrEU9dVnkkUP7xJAYqWdwxq9La20GX5xci3YhS0+zFhDJM/5GI0eQBW3lfN1b8ZDm1ZqNK/n
3ornkYvuub8pmAsP+L+ONRnwo3XT73eg8F4h5er7qKu5ZXLqWVlGY9YNyGZ12DJkO3N652pC1SQ2
g3j/eZDIEMVUy+VA/eNTiFz39IEFOstkMDOjJZGtmXutiRKh8+KODgQqon6Ojm+kRZJZkIupEaFI
i+fUg5nikvDoD66NBQa3DVMPMnEWuUi2MsdcngHinmoAhHfN0VZeAdkVfjKee4LidN0g6aPFEUGk
asKwFODZKY9Wm16mHxbNqFdXRFjugThOF/eTCEG+QV4ij24OVixmjdrMY1edFNYmai39kXhMlC/s
TPd3Ceiwl/qE8+yNSeVBPgHh/db2jIh8a/slijJv7vdbCHMh3oH5OQSpJ1u83GDfA9DeKedDOuWT
VgV6UXu9QCq8FC58Mi77ReYZfPTvnlAfI3snDAx1WWNJb3l59leceUOLP+cKzrw/wKhWY/QjkmE2
g5egvPGvgNxhzhjLmL3FQHJ2im0s6gW+FrlH5LkQ56yNzBuUqWd3MmkNkhaaPaQnDcjz3SUVNhvA
fJdsqrRONnwx0dTAhHNF3UjCDJQfn3hDsjrRqdaS8e0SsASL+qsW5/RLjxX3tc7ZVOBV6jqcHMbt
4aeGY84VFrlT7l6OclS98ljecg7rEUFuK/nc0QT/hA1ibo1etNow4HzcdwK4P9TJI2Rn3xLhbtGM
curPa3Rd04Ukw45dn/bBIqR/HeG0bpt/Dd7eHwLHWml4i8Dpkem0/WQ9RJlsbCQXFXFQoYTp/fm3
o4KbDRCwgsZ16mzjSedc9Y1pytgKQn6gQLdheJKttGRHfP2Rx9YPjS6+6lgZmgJ46rQU9izYp3i/
p++MclnbcRv8cCq9655cIG/h98+5Y4JjrzRZLX/IlJ6lCe/+HQzzVhM+OjlBM1E3bQw77vnK7Nh4
Xrtkl36DtawTC+ZpHejzoi51Cy9O+MfZHuRpd6yuVdXYtgx2LOI/rGse62IU9McU9HOCqn+05PtV
GqHD/kp7SnW5ix7P4lRRrQCYcQXVXCX9NYRaQ9MCTuYf3vs/bY9KN2aHyzlB7AtJD0TNMmV9BnEG
OY/oLwEsLsZByolj5KpCBMa3eqbz/o446afQA+46BNs2li7+ZDk0UvvdJbvspJu6fWlF3KvKgSCq
UH6SUIOiBv4nzDZ5H7CCntFKlE6jzJZyWr26TQ4tuLx46DhyP43E9fv8LdcnG9dI94LA6zBb8ixZ
wWX0B13TbxdutUWn93OPBRHSapE3is0Sp4fXcoRSlWx0BhdTDNyUW5OgPvRbP6h911ZRrf9mMTCj
aUy+l4LkzYLDGwQO2zgCWIG+yqqnrWWUgrGsbofKexNpQCkdcoX1l9AzI8xL146/apXtMjSf8kUA
Lf6Liuw7lmP5eFd6G2sAFbS68SihGjsCsD6v3DWB1NrO1njwkg9IaZy8M1iyJ9CoSuyJThqNajpB
QTpEaNJjDY5eH6gNEOMhtjwGPEI19C5VfN/24/yVN6uqddcEyOngKff3lxrTgSOtIjl60XsQb0Jn
KkIVytAwdYf8LBDngJl8vHDc63FpQsteLRm68WQPOrnqfxFngK7Jy3CEY03MbH+50xKPSvmoX8RS
6qervOLL/43mKHdrGpF7/26u0zgLQ+eOFS5VCZytjFbPRxv/xgNF709CXzRjmiD8uSH0PmiBJXtz
MajZO/nInPjuU5CBfX94X3Is9TlvWSnjNsob610tDuZnCq9b6pBKPgPOIbUDAJE/7NDIVuwSlizS
OHP69oYdGtckoxdRV2xERfBj1bv8Ppwn+BDIRXaJusMMLwgU115LDlmN6tRqJm7ysme6Vx+uLNrs
yiRh5zoubTjLDDELzIoCS50kQ9JwNJey2ugvbF6oQ0okWyvSUtid5nurRPqPFOeGfz+IEpAcFGZj
GmFo7bDiHd94eCOxngblpxsGRBYbxQtE5SWbmVM4NBP/S31lXnnq6SdRKC+ZxyRQH3u5peUpFTYZ
W41Y2iSaHq0ls8F4gH7e+gk+UK/298IZ2RyXW2VsBQqxpaLMYiD1Je7/V4+4PqID4uY9u29NbVAI
HDGse7FX+O4MGYfo7m/+nHFGK9AkJSj73FAuU80hUzzzmsyDsWF6SMt69BuWGIHOpZ2KoFzW2AVH
b4c1nxjNKsKJa7B0hmoTlP5o+eoyyhiROrYbLgvdUqME+hKUCCjjsu1/A4CwnPEpJip/24spkWgw
hoj2mL+K79slpdPlrx683Cn0+etXWidmXPBWm3hrifDZS6lI1qtDtgVvRlfffymGAhDxnaY0p5WR
4aJhU9qkzatiNTw9vHKkw7cc/dUlAz2vbRAIT6uDUbYH+x5TbHAMQAU6HHhIpK6pMiigm20lPODx
b5XvQ2hQdepu9KQBCB4huvHIEitvH0lIku7DZsmGMTpL+7k8Z6cU5qCnkb7HWk0lZKUkF73owOmM
AmVmNBQGhUNXbYyid+msrn7Kp4QvegKiNRYvtmkwPvD2xBgARchE3Z3vqDr9caMtOuGkIIV0LHmk
tPo+9aIVjB8Gp9mFUYON0I0q7jJ5K18ACpwLPnupBlSK9EgHIPQNPYcMFnxDulbCv0E1Ep7MNnj3
yeEXN8haIClYsUHorAegaxyaCCtMCAaUKCDbDiigCXC6+WInLaBuSDq79RPqMnjj2TL0CrDsnYkP
wvXpH0LS1zSHbuX22G2ZxtMgPItsXc16hfqcIoMyVktDkb2pKtU8O/P8WiZwfJwqsci0Ty7a4+L/
Bg/TVJ8+apDvDhZnIKipDVMnh3KGrAeUlUYOrBY/rin1qxKml33Cz+uIzbU2DJpM3fvmvfwAIIEN
gDj8L5qS72+nMOsaO7POpijTr2ngr3vncvze8dMof5LRMBnHFMaDLf+Zyoe63L6VKDod+qwhII7B
GQeVOPgpa0UvyQd6MXBW6TnjqFr8qzRh0PfqsOAHJvBMWN5cPmwxXR8UZ9zzDlKArJUu5EHjRVnG
Idm3iX8mUQ3Ugz6VnoqORfDx/ECx8aWTF9up2+fOee/YHps1ACLeZ/Lx0qKeOOiHqglKifahrMk2
xB/hkWquNuv2WloDvWViAFLsze3C8k5odeveyEaXNJ+8L2ojdGuWKMOFVRMJ433WtyI55F19cwKo
mlfMIvzLdrWgRq89Fpd6OeokhLSA0h0e7xKbE4bw3GwSXAj8kOa+keKud/sqMViy4PSYNRTX3MO5
hMRASWOIjhWay5QTFYv97duX+XPxgVGns3wO19jEEO/TH4nY2+H/P1COdvsA0Q7u6r+v8hD48WqM
sQIgyKC4P7Qo8RURsdHMKfrseQg9ie5RPYx1NRXDV0zWUViavrvN27JAUUSSMr/JRe01tCzOvdou
BYvJsPNkBtnPq6hzc+bT/PqfTIpPxnXZ60vRIqCJx07CuW3zKCuKXP7bX2uqVZSUCZyiySwdqTsw
VZjfikFwobghoP6qSU8VjCF177OO0khyO9k3ZIqivPOJN+aoa4JjgSn4emB/2zsgNiZYvrcz+uiE
ekFdVWwycr9Q3kx+6iaRuPZ8d36qhQ41a+N8I8jjXxz/D9UfSBx6t8iNUI2eIcGq63hrgrYiT/Ve
nPoyHLMK/pxUFDFUOa4ov4P1EItM/NHo06vIY+SNvDFozXNbM+8e0h2eFttAWwTIZDxYfSh781BM
IVEk6pAPAen5zMsnkezyXx1QvJCgqbTixO79wkA+jDZetYs57KE5od1xY98uZ1TSOU5yZa4Bj/KE
AqaK++sjkF6+jlh1dzmqJU3fT6ZdWC2rs8AHPDqJuPxTzen6jD5zqxpGTfqeGSXsExXQY0QS83Iz
arUXdMpfSavG6gevPiePwOgxJj2Uf/HPl5S3QZA2ZAVcSFqY7rvFQ8Eteb1GeLyBpUFoyv26BeF8
h6R8aA0qrVN3vN1nnJXNftVwqedWBHWVvIJCEhJo9iw2F7XdYJ5yRrdkQkB39N/1Ri0KdJYz1Y0e
z1x/SyOb6SblzH+mSxP82nPv7Hj7elw5LnmsNa68uniAIswSRpYl0c2/xG0oevz0Kp+UXolOBazo
Bc2MF1NOOEpVZh95n9WqxyNgAfYWly+MUak0W/25UcyCXOO3h3mWFVKO16u08UtpClElWm5dPCpV
pwO8MloGmGgWX9Nc3DKY/bBfo0bpsDeeXWSFtfMCiNPnHBT0pE+hrCbxfo/nMnCtzUWvGNehuzgV
3IZ+epK+ZPVkB8ockIlKethxT7Y+iASTgwsdNvoF4CNNkRGmyHFDs+LYOsjUAVjaYy7kdidRlfzE
bEirv72Z+Z1KU+BmJqGNszchio4t84KjwfkWJx/dNaQjc3744cRltjQEmOWZvaFMD5DV4zBpnoGX
qxMdHWqeeCtDXNFes9DN47PlDe3gBYBRZZ+xsvXX4EVXCJEFpO105+SeWAdevsP5a6XEFQo3M0L1
4pBoWfIGBhNu9xD/PJVFKdSVUjuGdPe/dbs/OhgTRPwx7RkqlcFuXjcTJBszxmWHbHwR5hKpv3KL
T6tx2laOetxToeV6nsm7OBLynpaK9DfMz6qaSxvgZ+AU+NKlJid9x5u0WrpTkNkG+jQUhNVaxPjb
WZSWOkaXaTzYqZdnc9wvaY8PlFqCDnh0G03Lbjrgov4dQ+saI+QShkMLes6OnbgxI2SZVTudtDkh
kve13Q0mm1tsoQiR5pvR2+tyJ/rb0cyMckeTuinapCw5gJoiyrbbx4IMGuTd8uB0cCQ12dJTuYbY
9li1hGEOzpquVlGSVrtpG5asP7G5msGnlQI4bYO3e/BhXyDZ6mOHzWG0af9LWs3ItHIhKRkz19to
eRBBCmvNyBEwKu52NFTP/kwqy8Rs3XbZDGh7PmIEZYt6L0+BXr5nwRZdw7YJP4BNFZqGoDkQRRp+
m0/iPIy4En7IHLCDImJPYrqdLSfTWp4U3Zw7TeNKGMvHsYrQtT4izdc088Y/umOgGMWV/SG5jTRb
4neRZve18cyCjsvipSiD/TIO1H/v9PeV9XQJXU+fkAhZhIt69bjvEJz6EEkHW/T1OyvfG4v8eSCA
vpy5D9HnVl8yuYFXa7re/6cRzIDK/+9n9Ma+jHyyRUsBtGNAo10TG23SXWdvd2Wwkmp8SkTZ/tM4
MOvCIvx3nx/WoEFYBCgNf/1Pf0OiwfxmoyMKiwLMGMZ7hKUaHdI+IsQv27uil0bQK9acjqGhxRKI
gOKiVOwSNGS7bCL2enXr93q0RKFmQzTcWEANfmuOVJ5Nu9fvBCRWHqsL41TVT00PK6rmCAfRgh4E
QTyf3gP937wKzhZdeHO2RQvVd1iNy7qND953nTEUfRh+Ys+Wuch9H7f47XhwratDSgN9stX61aWE
5JJ/jUU5X5GhjoiWA9Nc5SDNQ07BE1IaKHRp8zy+F8eii8GQNjX4b1OgZNfmMgHouQxUrOTWu6r1
iSF02l0O8gw1HNjTass0/qz7foJ8GXrUjlvrEw2FVwXBW4U2r6GkdJzNR24MRPtPERDruEfCgPpd
mGqBpFx+e4oHrvL+PVLuqHPM/9y8bttlEpeUbHBAkrF4EgRlTYo/wCR6hWc9UJL5lzcjD4n9imFz
BHndo5WmWIClLmUkJWMqPG0/qlbLj40gPdRTzcMaKk3A3X6W/ivOU+PLHt1s/W27WqIdpnln9FmF
f3/X2W0/LX/tm6Tbig6ZLs/a1V32hjKSpePnVyKsbrCeJVijTcgMhub5FSwI1DMXC9u9wzZMAhbp
qUEXuEmgQgEM0Ct1JKzTp5hIcSM+yh1q9zl3IVZuoTd/o+kUkti7DJgmZAuZI+tc4MYkUXbwcg2W
DhaGHCDBBeLhAA1kRWBrsO0oiS6MvjR75jVTVpT1OEb00fq8JmOFKBvYG3OK4Wma6/RhMrgMswDE
h9A3mJhlTLHKLozJfUFbRBbNspM63yeaqn9nQTHtZlF2odFojDH18sr7UWSp+Q1fbLd9V+8J2fc2
eCJcUqjpuCM2cgBGBFTGBdIHa9vpiqwO+uPZE3mVeDuPeq+81guLzC8lMIuVmmu/Q0DJ3pQ2DPt/
aQcZW5F8ns/tywlO4vA+VBhlx6g+FCzisQelnxKInHJM68rfXIInORwCqacUSDiQ3W5uF0MfP3n8
9+tHgpYIARfA9pLDVKxHJ1k6GPaU0r9c4pmzz9pa5Cd99Khb5zKq5qJUDWNQ5Y4c3kytWcALJaps
3TAkiGXlt2GVBVqllbUdQ1v2c3vu4JosbLE/1Le9hJiHkwsqbUkfZX0IQ+QM5L9Ev/mDcwPXf1KR
sQRDPOJZt9+MJNCvthMIMrr8d/GPXAGBhM8WAIuAYsvxxXqi7ikv+cuqn8JWbiQdtjmmbSSwTiBA
3Nodzrm02CEyFkwHoJAMPAS3PPrqgO6NUfvH/Ux1wgFISgsLEA1VJyn5iPIvMoF+NutxliFH6nzf
r+vzRf68hbBHbYHahFQpXdVclFX+J86i8MbTJ9tR54x0HRAhQF5Ebw7Un2VBuei4AOzaE0t/za0s
OxDj1dkW3kWdu3Dt1i5JEHECj925UCmQIxOCz6lLrbJdOz05bn5kN50eZ2KDKOp+AFaywe5jL4eJ
GgcMDFL+IL/xYb362QwC5OiOmZlJQAJCEqPqcO80yCJTC4f+PXzj+4zhDFoZItmw5H1oay9frcHL
8cPheOiUvGrozU4NY7mQa3xbxaqYUr6RRhXQr+Wjx8Wfygq1L/QKyhg02b6YeUeKv3WL9hrFiPTw
pMu7tDVSsVWSyQYUV94V/OXsNr6R4dcs1IyZCUrnsKaEocc9ku8UJ+M56v56XbF8Z9D5B9fXwIyu
TQ2xnvcpGafT6gvGlzy7vBybnKu/JsJHVrc4xvaIFxMW29tCLrsfK2jtSkFqeHvg9Qc8+ynmEDh2
H3JHYd9FJFqD4Xvj8hXTSsp9OGy1B5kvtDCpygW4jmWCAm8/gls5/OaZC+ypce/XxosIOv5cZrbO
GJjN/AXCDf04MiwAlts8ab27xivmJ3/Zr4TCGt4um6YGyUS0k1oqp5UuYRQWe25Ka0ykXW9EAkyG
4+pu5RN/bb5l2b/Ek3bmxkWCL+N+5+U+5mSg7ITrgdETV1ewG4O3BYTRm+xMj86Ho7E1ogQO1oWx
EWhj0RvTTVHO8yT+kaUI3NKiqa9PGppOdC55vzOEXHAyiKOvZJhZ953oeuPzzkWCdxJeAC7c9Bnd
TEwHb+tq4d9NR1ekejkq7OEAbR/SIBaaGQaNpm0gOi/qEd1fZ8q317VZer04aq8dQGYJ/wzST33J
Q0ZuqLurq1oys4le+Dqt9Cep/CyMIJIBg1AvF/gP68tqjFlGThN5dC/h2YHD6t/1sXLPEOkPgji7
GHPSLbyXrjf78C4i2Z7rOcSbGy646ly/JVuh81XCYW14x4Pneo66xrVWslY0i2gW74UuyjrDHNO3
xyX3Yuflo4xWeYfluXcu+cwuL1rAmJE49FRNdGHZrD9Iu4RA00SwH60lY4aeJ10xclu1oIOO1hj7
tWak5mHyM13RHb+KEVpADHTBDB+425JHFyAMsMy71eMH5gtZ6uBEJPgVnFeDAaeEx1iV/c6qdvTC
snY8o6Ful71Z7UqxUqrZzp7X1AXL1hvY+dDvBmWXcYwmez35RbXPdGMiLF1onwDePfa80bPDJCdO
3jm/iC4SfBn088TTk7mNZW7Ky9KK9Tmmpj8urE4xNIJelHlTyTPdl3EXimax9k81lE6Hombu5dci
XylaH3PXEnzCwnCQgk+5lJjWA6dnBMXDLSCE1iiCQBzzC4CJpm2NmaYSRbNx8Sv3cYS392R2V3Mx
IRuodHYguiPZ3KzPogK75XqHG04DVj/Ss2qCxozMvIGO84bF67+AYzGRbXj98+LoTGCa9ostSWle
VemS3ocals1M6xdKCuScXzaacZszKIQDH8kqVdoZ0Qe5lBRjViBx0By4rC6d6pb7kStmyjMSt2fP
Kw/qx8pQ42sPC53Uewf1kdb9a4qkOBUabKQvnzJvAAXxCLgvhwkz+mmzFFCsoXrMWTs1cWW83dK3
jEp/EvweRmBgaJqKh/us4VRFTmrB2sUDnoL2Z8Q7sgBJei47TgX4VghsYuB/A9H43xScy2l+a4LR
uo9fvMSGUtL1F1o35gtOOxxw3KydQF4fDnxPowPplO68F5R0VhKP3fDLWRhtAWxLzx0lIhHXC7ym
61AeeSrB9emEIwGqUJDtVXyWnvTzP7fRDbhg2rzNfkZAbEIwhNZpDcp5Q0wQzWczOlYAg6S9cCFd
RTTI3Vb49+KQfYHxJ+52v65hB3o7iL5iZ7HhMaOHSj1esgqbbMT42rcb8IL5dyGGwn4FvgeqocKW
jQMpV+1tebOSmmJORg+1f4j84FzVg/b6vL1FSAS0UnTToHXknCF6zxKNpCkATKz/r3DulyBVIZj1
yTgpKvkWuyDpBysrxiH5vXhhOcREFmhQZQkusVuya/0OU6keVV7X02mvXl1GnqjagsI9I5kz2eX4
2jiS60ZE4MyT3N/2g8Ou/Pihjdyvi4ia94kroZs0cagpHq9yWRs4s6ZAgzkTBQvgpSoobmcjb9sX
2+GuX+Yg8XqkB6jY2JNkxq4oKl2V71xGwpP+Mb5XoaNbUDMK0JpcbJFlTep7dRSdgUfowI2FHTmw
Mxo7lhuFdn9ffwy6K0B9e1RvJtGZSM+e5FXu1U7xHTHcjDKHvReicJLgrPzw1SJ8F24ozO78eI3N
5STkMYqqBu28xEyIHWtPu0itAE3hTehD4X5ZeDuha0Z/0exsgkWyV2W9FG7W5tWVHVq/rZ84kit4
qZJMdeYDxl3vZyH7p0rCw31Zc+APLHtmvUseCaRcPFdnYEbFKeXqQwek8sI5g1LDMUk4fztfkXHX
Jua0ccQHz/cPjWFsdovs5xjkmhJby1PCg/zyMrzHI0F12scu2k4hqyIj95uBsNBhayol4cBsPfsG
oIcXUYnTE4BywFYU4eKKUu9G7UVaH0jC5vUvjpow6QXcPXpkOsZEanVLznSbS8ObQBsiMqDEP2D1
0B+B0MkczCtphaoWqYNsxNuVBUtg9mOTnwZF2qsJOrc/o14BKRH/loVyylJ40LVGU+98a7tQ8SQ9
N+unh7n/9Z/XzaqrGkow46PJint7y1zk3uZFcq0ozebK6+njRwB8ZtrA/3+rUco97nAbuwS72dJ1
khzQ9brImdLVk1VR9isroiJs7T9pG6fb1r5QddaW2damvyDNbpDVNpIyTL7SOhmGmtqqFeqfJtqk
fjHgmw1v8SCkt4QXIMSI1dFFeNTbpNO0Nq9+TI4SWLT3Snxu/GQkczM/aFNaBJ/8nYy9NEycYxOZ
ppvpYbyhN3u9TSQWXjmnfmSKwHE1BBryZ25ANGIGT54zWsmlj7syWb61ua3ImYAvbBF1Lf2Ugrcb
UoCjABZJYP3BzGrLosaMWktN04K9PWaoTznbvQHK1kcwRZceOh/zh1T0EeVUTOkH57O4gSxPtv7S
DK3S7YZ3q/dULRncttR4iGKpurinr6OLBg68hNK/4zNgrT8Qu7AYknVY2+exPy1gTH8M84LS78er
SXkbH8ffqYHlrE9vMmn8z6qppctaqnwfJwUn5cNI/6mRkzzLfLzaMx8/lqYqGqWH7LwNshUWgkdl
cvUz6lpf2bAhrSTkzSJAoeie0wyVk2c6MvteAOAIqQKwgrCuRAQkyUS27WF+3FV6apTdQz0xLvDp
N58ALVFAyjpeE6wFBjpA8FfenCe7rzn4KBc3I7I5KOMzuCinSFynojL+3O0BkqZ8ZA8YWLxumQvs
w0gYU04/ZmTWS2rsRc2tv7qCJAgcw8Gpbpjohxjpq/gou7SO+VfKbyLvvyLB64uR6AUsxIlXRyrx
X8qdssiFBNcTZbdEctELEfGRzFwRTdiex2Tu0vArz1RiCCnvdouOtrpgUL+NX7/hco6EUdYDGExd
9TMFTqrMhXC0F0rBQSQ0B+9SHtBbRrJAewMrViIg+6/t7Gtb1Bj5qz5J5CQXuI+B9WHQ+wa5s7mS
nFUXifjmwH6GiCN/NzmsQqHFUKCFm0zF/P6SFzUdHBVMuw1ccPMIKi19Vm2L5yNK7zhyggYXIZCH
6uZ2saIO2cRDVyvEKt/VZn5miXBvq238Rbx03TTKwWRqZKnlUAN7LWT09h98hI/air3Tf3Yajtb7
IJRpWWiaZHvCqjSBbGMc9daf/3/5UKyrWnjTk2fmiXzOisQjOxRzzFMVgO9Gbbk06htCZ0g2K5C9
qagetvRrwpOA6ipZugF9kEHOuJrpUGnCT4cTwIhPP2N/Itmlwc3aHr75FXUCsGWyDKtE7YwBpc4B
hNV29oE/oFmDD0imZV4kgauTxKAegqBDKvsL78aigB4HWVC2tWbXan4FKH8yduQTj7u7Mb5ahryb
jSCU1mek/tsuYkNe1OLtGzVJuSj7j5nEWhy61YFcEFV+YnlJRUfuzPU+tAyc4VkWMVDaQ3M0FQaM
Xtql9WQirnIj+tooLpoEvEptPtYC/kpRD4rJjnmcmI9ehhaUFYhG2XvHySLC/ekBACZhRx8Bqt2v
5OiGR9Ci/PQ5Zcz3/l27kJ451Va2FvrukfvDDNfM0SElB12DlcrjU79Mhx9dXVVDh2LiicYePp7z
ReLQmFqcvKqcpssb8Vo+ByZbhoxTHxgFj+7lzqVNImQlmTqhPCxoRiCf0sAEANMd/hqZALS2mmIk
bTRqAhgNBFO0/LUR1PZ42tk3x4GoUuuK9R296pdlDzlZaMuvWunR+magNUH/bcWfrTjrao5geFyQ
XYqesvAWnhMy0FW3sOoWhYq+bG8qwLDh4w4CVSwzj0877xwYISw9WohCoGbOM7btUfEVkvXb/yQn
9494abVZR7Qr6uRAfXPzS3fzLgZgPiWc29rsXCF6i5tsptJZ3MsL605WTGoHdUBHmKDo8x9YfsD5
SbQwILAROTUhScRslNCoy6/6+Getv1tchlN2SOG42UBeHIfolxIgAGlNTzM5rSdb638bLpunlMil
wIkC9gH020Fh+ZloPuQYEZlUiCewQldkii6nk5nWtK2eKVQwcdIXBLkrhxr0eRRUOo21ckUovtLv
+IGJKOTRGWH4xUoncZF5T26kiB49QXZiwo2KbL7m4GWPn9/iCrAe/mS5VfQX9V8Y2bnDbWdxtKe0
gRGfwaRBzT9biZbpnaabn8g5uCT+FQUiighXkg1wno1yEnSUL3HDmzHCowPbeZ6XYR6I9jCWr05t
WnOCEHwERWP87lZ3XHblObeKj6xKvnGVoNYIBay8KSA+1oYnxtSR34wRdkQJ6AYflhtF+vsza11Q
FEhLNzxpZBzxhnOJTzUqJy60HpJLM1H6as8DYR9Di45qQrtaN7gzyUtSvWzCGQ/M7WXN4O7WFr6Y
TWqWi0B9oo3gvUVZJOY/DfJV8yzrGLn2GPuiFpsKA7phjlTw1PsRVqBtOGcmoQ8zj3mFX6khD+N8
62EJMPu0NzxJJDOKBf1UrHamGU0DFav5YmBjdnxOsiR9PgPn99apGJ3MaAcUGhF83cyBrXzv2RTQ
rf/PjVzAW+WQU0q5jJUGwwjP88rtlzj92Sa0SV9xxt89D4d4bh84PxjmpyXrwzDK+H26PnVr2aCo
w6B2ukKmT0rtqQRPok+uYEl9JHtIC+AE5LtG/xw+OgKXXJTPXK20gxLFCZBPjmugygNiK+ud7FG+
m73PeaAdOEqKcpCEIa7XADo+vsSBTUl2KZ4GaGMVxmjNWtWWqKRJJjKkNRqIWyS3u6/qTyOPM+Ox
6NccJl/oGwzAhLjV8F45G4Nq65eELqMRKUmF+cnmaOxv5FEUOEzcXQBvhFPsjhHGe2+dUCEUUm2n
yUiK3ynquJiFMo5KKJ4M/z6l/g+68klA1zImKQq6rEKcqUty7li+6CvEJsHMkgg62/TWTPrSeszZ
iQbnf7vJ9bom8ZiY/OQMslS6d96GU+E4O1GSlzyJdzZhub8DR4gYewJjbsCKR7sYGyjVJaKhVBl6
vOM6HcxTvTfEVP1MTtucyN5M0e7gEXGIFbvMv5W7A/CVUt6Qq7mU6nN+oZZP0YLJinDgNWgJ9IKt
oDW9y1crFmOZdwajJLLmnz2rzWfdFXTQgidx2jxF8a6SjnzJn5SJnoqp7T1KdYukxwYf4Q4iZ8b8
+j21OH2587Q0Z5pRbC8keJ9ud6kw3YrFyOu3yyluIiauJaoVYaTMXt0XtDELd67RSeQamgL4IgJs
U7KOW122YgionOXlBUCqE5PBMEZnjrjfYz93EWQfWf+cz3noDjRkvvtY3SVvTfhCGX9rCukjqZRu
e9PsJESSvYuRKLFjkgQOi1StMZBWj+4JvEBOWoekRaTupPdlHNxqI5XxBsEUurYEFx1c68GtR5iU
3eDf9A+6RlAdfgB79xBucsW/age43E9gbPxk4W8qqt4DAw2Bio7C/0u1KMM0YAyLfD9yiK42tZ+m
Yor4C3W/2qMCivbYe8CnyTOQnV7ziSFFjfYEQy7aV1wu3orhdy7/N79tnB+GWkwZzElfX+X3rejM
vE41KsO/xSzBgi2TLf0enYrQti80fFig3H84TakJDixhF9UK8mJVyYzZQ0H+wzPFU9tqX4ZpzF10
l+syoKvuvdAv18x+QoyGQ3Dh9DwrEZdiERrGhg1jATan5CiOwiTkXymtMnF2n2kShyO2rJAilQ9f
pgOxvtY4rNQOFRMLGJYEeFiejU1M17QDRHV2joX4UVX5Iqze/tqW+Rp5ewSdNywm2dmemsW5GF0T
CsXNVW3ynbj2kGHmUW5hXBsF+g+WRAggyBQFLwWNnhtDXjalIkf3LB1yRFGY1b1STBXqKUGGKFQm
uQqXec3jmpMbJK7vH8tHJO9ljB3K/FjP84JlykyF0ER6q7321zFisUtyeQmX4w0f+m8KWqQdGqlN
c0pvGEx1M+ig0nq5Y9TB6bGAExaH83vYz5YQvkUQdwe7VWXF5jLGtlLanYZJV3Ay9bf5LuM3q2jl
mLphJG5LvdKFJt0pQbExUJH1bQybfT+4nliu0I9NScf8N0fHmP/SXLFvYYIBiHcu8y/YJFJNohqY
RogubjFrHKVjMT40n65qlJ5xBbrXDi9q7arx6qwEG7hogAH7OsUBuo/YUEL3ZKTKT1QvxGXWKxl2
HMkesh4eSYMHRUm014OpgR/KtRacBcMZ4nlswGv1qvcelC/FGwera+T/q62zuU1L2IADRurbzTwC
SXIsW4XS2EWmtI7r4KwIBYne0cHd8XsJTPNDlbYrkMRfFvR6nJG38qJ7Va4clNPPAq0QiZHtZnlP
2UZpP0lzGWqUcG5HUuVJCKE8HgMdGYUG8di0WFn9WdvYAj4LKYZ5SdVTmXDrp4QdiQWB6DYF9tiE
wnDuR23Adp2PZF/S7Xv8eNknSq3RZW6nHiZXxjBItEjO67kPl9GBvLCRvJjyCGyvNh3ScjuKchGV
udcJfL7MW6EMZaluVqrsgb2VuyNpTdpJyyZXc9HFnpATwpBpJYFKv3nC2vNzdn0KzTAM8jbGDDpq
1/g2eUMEJmGDchMzn4VQD4L4yFPnyBeyCpRJbZH73OT4sfz7M8yM3EiLBbNZoS5dN4F5vo4XqUHE
Uvj4wi7Nc/UPw9I5F59BCYKeSEGFwMHxB/pbOtetxT3fr2jCFyf8d1bKUt3HafCFLD77qSIWem4P
6brGqyO0lbXEnRXySy6gCEqQoDq4c54j3pheyG6edlXy3HHBlFn9Anh8filtjCcmXshSzdzjekf6
kzPX+55qzyhggnnIQmeohngtY0D9M4+Hs82AT1DN++GsYqTOYE4a28n5SNvYxIcpP9vlMcUAj0zR
Xeu14ySUUwoBW3QwG/qb4wrrmmqieCuQBY6B+GtzkvhqcEOep7Ge7H2WGPyEFu6o7OLX/V/Es1Yj
0wIHIlukMw9GJrPC6ZJ8/HDUVr0q+YWWcRWXJ/nx792W7Q0YdxAnisdp27KXuOqZX8kWontL137I
TDfKlAgebtFK1xgckcDpgwozHLNpVe6h8lKpS/YUf+/mH5bsOz/A1RJm2HnVb2BTDoqf72v8AJxp
hAoYe/E+9bY5abvrrOT7MyHKyUIBKRxHz38GRpDDpckUgQ15Tw6UCY+fshjGO3mqoZnVubFvoqpu
EyIh6Nqhbo6mWYJ6K9ArE4G7L4nYBY6r+BDPiFEuchBPxIuAG4EFW+QLr4sQAyynJEwJu/HrCL+6
h871U4xjxv8ljwXKjeOTKJPY7pNMqqORfJ36Shw++CA76bE5kqtvCUeXdIUJd6OL7QRFZ0fOmj3n
Zyk7KY+B2chx2MqWzFx4pZXNaJm4dLDkISqpAhdXzS3tKm0kvmMyBbDz2o5qrX9IhZTxpC2DeBtT
au7+pZEMqnnth2ap2hpY16pyMQxbUU8ujPzx9qhPAt9AWlctB0osKT2KUe/QIx27UGRUPWkcHSWx
+o8g7AZ1V/FDx4evN5DeH85Wol8UZpxEVj+LoIarWW2j+VxMD3jI6GJVT/JIgFB3HrZdmPEQcgEX
VT/HE2fDXJpq1WuM6V8ZtKokBCeWHTEH3MaSMKsR0z0pyzXfuTeJ0i60JOHA3xK8BpUWNmMJfLZf
SbsDvCz93uoZSJ4/FM1AVpnuSUE3TGMLdyKM31E82F407e3oHew85UHnmJ1OtkJoSd4v7NlgYStq
pFrJb1lkGnE7KEQ9j8wGR/N90WpVjuqBjjKA+JGFraJy108p0UH6hqdzPzZWUMVCiuMqmu515lyI
Y3CCnPsH0gD2ZyqFrLkYN5a5CDGkbv1nLABtiyFmKmW11jpCvgRhbLXY/BEyHOl6CRT8noae4WEo
nab5XAeA60b7efuJkkGlQBEEv4FX0tQb+Y3CpQKpWCC8vWKHWCQvq/SfZ7O5P9HZzJ7sxy80SVrR
0bW/HgECpJj46u4TJnN7rU8Mp0DBc3psEK9JFyEy2b2+kQfga2DB15ypzLAlhnrn9fBbawcx4s+l
hvOYRVOSA8YwVODHra25OeoXrAJdqiXXCO4rv6QpdEod8z0gNS1iCCFeUJdltp2FNzFHANgilSfm
ilKWrL0noQUYNhY/9ViB4NjHZkIa8/celSheDNtmLHxEAAjg/wPq5id3oZa75c2iykZewC285SWC
uBbb7sThQg6y6fgkPlCtpmTe2CIFE4jo0V3PfT5fWW6lffskJqli+oiwEaihfZUsxfFo0evC/Z0r
K48t8DdbrpxtBRrIcSWOmnGccHBY8FYj+MwCcFLCgGs0rYfqDxxVAcJeACj4XPIxytar2AFayxMw
An3qeqlcoO3yhcPBIDuQ30y2y6vDbDSeWM7ZwqXYyhD4l52/XNN6h0vAKVjYV16dGLfCurc5u4bq
4yPnidXXxKd1R61aqba/ivgpBj1Azj+MNCt8YS1FKX03v5S01BjCsDqXr7NZDTXGDTWxyHg0gpsX
/2m5/CPD92XdVd1qKulufdyNRhcyljZ75Wn6NWDlkAV4KPT8ZnBF5tNfliG+dwPhkhEn47LxPpOO
Tp0RVSiEZp/1WMJtJd2vH6zNrmQ52lgBDRtVxHKMdmKIQ+37bw9EuPE7lRbQzPkJnFSCMQ6xGndp
sTmYrRUa4c5TMve2O/fjAXhQ1K11g3n4xkIRgDwe8LcApUls7HbkqCPEH2PKPDBK4524CClsVeqk
yLXythPuwzkkxH7T2ZbEwr6zpnZ2bXUlkxxzhM5nKepn8FbukHmlg0ngCWHZF76l3FUaO2VjCQdO
UmWXe5hc4Al6tN3Qi7gcnLXhBARU/PKUDSb5ien/ce50EV/oI1W3rQXHcUg7NychxNYli+H4w5Sp
jw4ZWFkIhjkNOg76JoXrrEYXMhVzs/K/0QD/4GP5OeDWAdVAjfdhYchXh3BpDIE5C+GGscG5iC7I
tzjLsE51vDspcyT9uzak06LzgeHYtyT633Dz6OEVStZhHKB/CWSH2E4GKFAdvmRkolL1jkrZaxGC
6kEVXhKtms6fSAG2xT55dQzHQoP56W2hpw8ooU4f205cCopUTzmyFAPoUa/Ys4I+EAu0WAAcYTsW
WA5v/0xfVDtR9Nenq2I7Z34/rMPiQE/FV+no9tUZ43ZGMvaACLwPhLY2xO4JjbKf1QNsQd5BoCic
P0+LrJ8iKIXgC9uFQ8yCz4s2dbU8c3VuYh2lmtkRfcCLWWLjAf0s3XlECp/lhi7/LmM2nkJXTGP8
UTXECH3NlFBl++Y1KMwEfgJJZa/cTUCGBTqew+C10w0OiRaJkwy4L5JYbF+LXHjfnGJBdQwHdUPW
COWDApS5ZUBzsRuLqV9HUL5C5/3eX2q9qADsJ+nRggxMWuI/tutUs18pKzsBZlD2Uphw2AJfaO71
UtTwmRgksBcDthEhH+7GOA8BMpPHDFUwRF4CxO8h0qQ9LM/ho/dLNTObblIydde8dUs7ZjJJy2Fn
M9lrrZR/ChsRcM+bMJUAOn/AsR72f1RoJ0WaDB6ZCFCamEF4QpsLAWpc6H/vjkpuIvyhN6SAkzS+
mGihneAFgfrm1kZQ12CbaWMrUJuxZo857ZbxZbMP7UCoZS0ntXjxzL03X5265VDICwN5ze3RyUEZ
uQ43uCSBRDbgbq6n3paf9c0ATP6qcT9H253rtRP/+yiuTIAR1sOhG43lBKj5t4mKAr5+XNg2NY8G
kMfg9/4dk/omoxUa3PieP+pF60vmO0zoRS+jytbsIANCJ8Jnnwh1PVhhf/onavpjkTcLvD7sgHq8
CvxKocLGr6IX3+gn1khZm621evbGcFaevgBotzdvyKLkFiA5Mxgkz+Kf4QxCpYMwF8jRzQzo2KAk
WGfv0o/qxDT51dko+dbXMPWlwjg41LIrJdzpSmq8VMUpVqdosKllUiWS27GCmTLtN2DvKyPVmNEx
Jh3D4KmWWqx9PZo4nEVBtxA+Gml5AJJgso0qBcXpESnWXvIiPwXQtqbxcWPyFF5uB1BcsiG3nVWg
/0Nl6/E8JmCsSBdIAD057HTdzL6j3kvNEmxYyhpsUQMd+/YxOzIO0vaAoECT6SDoL8T4dAhVx/3L
4+6ek+4VDeIP6OKZitYKQV1NVK5VWsd6xNcWYw1xdYZbnssYf2yG4NGus9pZzqbjyAU95TJaqfqh
atYPQAF2vOMciFOJXw1VZfRiuXEnIyTZKoVqa1C0cpjTzC0Ye97Fc7xpDlN06Zm7P9QaBJpv8HW1
CR0y16jmpQ7AC9wcc1jQIohtNanDFWZ5mSAJ7HJm+PiKCYUs5nlE1Z9Al630nqOEIigpziw8WBhd
CaBrnKu7O0kCa6UxNxdjy7FwPy/sM9DhgHB7ERh6yx3XL69FUoym5QNjhgqLeGlKZYvTmPB9lzpb
P7jSLAb4fJWd0BKWJB1YNSdUh/wRvboyzr60r7rJZpWIQTMpB/SNv689UYp0OUegWLdx2t9IqTi6
K7qiin1JIO1Uv+B3VFan0X1cf3xebMpUe9qjEfMoMu1DwKixV/RWEZ262DgsimbL2EaLUHnfPLLY
3//wnxcQS1AHB42LSIVYjdZfhMFWoOTykDD7JC6UBzTbET6n5yu45/C+R5LgQC6S7RwvI9r2U/Ve
oFjNnHgdUKqgaqk7I4gbUO3ktFy/yQ8Fb9KfWYknWlVGPskjZ9wZ0ARAmXwsnYviDnmemRVSpI3H
lv3W+HtjtWS2vPKBRpCLkQAnPoV6tYgcbsGYXrH0XYOb6tmPO6JrM55GUA+gfxOiqp+Xz68h+6vi
dauHYGSYAYg4bsvb8Tp04GtnqWB1DqVdF1C1XYFqTSsxdM6IIzwa6GxNrpd/Zm6GTK4z1woIZtsl
PjQp0IrypM9I2rmlYtkj9ceOA2V/42KW9IovLUzBBRtHLAh89JiGHPrTfunOhcoCmdO2SDZ0lqiP
2KVKnrrBW3ocDHhqk1VadvpMj/1ADjL1Eh/ARUBkeQbaf1/HXQzwb+3R0p8z1Tv5lB0TyDCEe42a
KDnBeHf0UIPov0DYX7yrcOWAc9sslHghp5MNzEvS0mUGDGFi062TKT8l3DAicY5sHFwI6ybnvr0c
ytl/f3KpAyS9jfyZX7pkFLvADcexCvziWBQltHdQ3pMcl5aLYTCab6ryCUyuu7MqYDX8RfuCpgXo
ERgzL234t/1P/i9XIaAE3S7yQn+pECcaQWNtXPjZKvTIE5E7i7rGUhTIJT0M0QRPVKjT5hznYGpZ
wftqWY7vVjRz9eZr1hl6ignd14KmwpPGCog06LOrtE07624tlR467U2Yh7mEvXa9ne7jOikOBE8o
fwZX9iNZLfSfW2On+lilm4MPz5RLftpG/mr8BZHcge0VEblpSiBbuBnQKErU2qlmIo1xSdmc+Ws6
+1Emeb6bdvr5s8Tq5iqTBnuIC0kQ9cJo+07jH+XK5QD/y2HuzRntnYEYrGoCpuIaAWIo8wgyX0ck
0/brTfnkJzX3NEd1Mm780DbOfCMt/m1ZzAcJe7WE7JEaRUw7xfV7JfFhSixbgJYcZYamRlYswqAO
xsZVcfd5EzmKMCmEJHOBz3s1swVZezfhrTUPMfJKK+biQCTRP4d21xUExS9jiNPjjKKZZU7x+axE
NfhBEpPr+CQAbSXlJhJyY+Tu1L7S174q/OQb3a2qPWzwQSRbywRsu7pdN2qAnpZcCMhVaX4GqW5q
DaPzLLlrBtxfPbDJ7C40vJYhucP+yQbQumtcesv+G+lruFvDA2BBy9bnWc0IkzI8E0XZDiFS72BH
HVs/dXpF0k8rU8Rm7SmJdP0uGYE4BVxiowpShMEtOeQFczHHwWovygh8Dui+ZHwsG8az/hkMEeAS
GTSRSSc4rsTgwk+mfYOhI1Nlk2Q1C0HyC4k4EF2ycUhhF/EpBbOcoHXRLeGUBMiLv8yVz1cLKXjj
fvu1BeRVL/oIAq1O70Hf/JGua1usa/qpXt290StezT+IPUQWf4Ln/T6y4s03ATn1lQMjGUdnGOUM
FosbeOc5nUByR2e/hEZ6K368tME23/uD0QgYayYKSKS/OS/2ftDR1Nd2nCwTQ4iFKSBz+vICKuTj
bA9QREO9Vvno+xBU8zfR4Qx1XRrCf5W2TbLGGzOL/XIaSVso1locV5eAsrxtU+OjIFCnF7hcP7jM
1C2Sy2q0yN1n1pFtQpO5NswwhdK9rUjbMjTcddc+MuseY5IwkMBv5iUyO5FqyS+7UuvPBCkM7hum
UaHWXjhYMAF6QSrj+b0UYgdEhAyTzOyLJG0PN9FtaGHRVwAQtX7H8ACvrJ/JO7nMdzRARCM8baqf
KjSz46co4ZJV576yGRpgCI5FNFzIKwRv1Hu+Vd9jPAw2/A9jZtodSc9RnlYNOT0eJ9WQnbbgsSnY
i0yt876z0PLWVLFFOV3QQXx+A0XdoPVQqY8SdhN0lVT49M4RVSd9qadsjTL/f5EGThjLYKOoZafz
XvywMC3z5F5NTJqCblaEXMuei39h68CQBIJmuiSjyh+v5jEZ7cdSLN49BZBylTQeRXtouvbabJwL
GL5ItlBcjoConOc2hvf9jukbxUoDE8zJAAC9getODgMRF7kBy0MYpyGHoF0Doj/yzG9pLXXRqzwN
imYDgcZ2YbA6Fscjoxbg49XU/2SQciHgu9kikSsREj/fCMEhNP6/dHYXjkff2ygalO/UM/+TKaPQ
m6gr8wfp/c9RzKXaqdHalNb/NvINV0CEhwEHIb80yIV2C6OjnWSP3IBYfdvlGEA0Nts9nFxxE4Ac
I8spoasTC7Hi8Qw5SD0EMpZ8qLnDk5WOwzsVUszQy99im99somJfQ8rZxUEyttZZUDft3sgwsjJv
9ClIs+8v/w7mkzWGPeNsN+/mfJojatiRyF2bS025kW49UgZxwy9sfxuYH1KJvompWUIggoQDHTYY
dtSQwusUy0TPdNpBfRaePNoRYE6yhu5KDsBUNDr0rqRkUkBg2qZo66GLzuQ9TIHKPE5e0wgxVski
mTOLFGy78sDgDtkav1onIqE8CLyCbh7mft73jZVJC5iRPaHqysSre26fAe8chrmh0S1L1lfmoEND
whBcorLwddiwnJdIMKo2jWBB+A62mYphnC22TORvZvHejs5yN2+iopT4E9fcISRraU4d20KCY1GD
d6nodJyYx+EzTnCs36K/wOQZ0z1O1zesIjyLcExonbVc9rmBjr7Jsu5uT8YuDN+xhuXskoli5tRe
L+EsjNHoYzJPcolqKsv0UoQ9FmsV8EHMzmB1wX1E9Ilc8EH2uBDZSqbQlR93oVCMNtPRf8y6711w
gqvbE6IkzAh8TP4JYXznlBblc8749KTKYSCnfw4iAKGKMKgmnqAdPo4CsUnhARJbz19wFg/tI5Jc
zsPwh4YuCVT8dciTUiUFBUyQiNCdLbB5EtIPqnV6vHZm3HRM0kPvIP64toqS69xe2GD7+FuSlWdO
IR7CcMGnglnsI9jnHGEuLtErkrC3KEF/II+idRR+YQ9U0hD7kBg1Umf9qnCkxuo/f7Z6KtBFuJBA
XXzYLPMCHhdubofuWZk55wULXBkt/NxQ+ToPSN8guLsL7bh1M5CFvSlvFuM5t3aM2ez0gwLqK+04
ylyIoBSBkdtSTe4FqxolKAXdJvKwpTlVdHqMqNBq8TUUXCBRLEg1NKHoosnkgzp2x/ygZMxyu/85
U4xa/5yZ+p4O6YaJ6HcrfCLeenP8Pl3zAMET33UDhIi9ELN8Xau59jknEAaB1F3q/0pElfNAtg1J
T3PUl1pxQrBmelr1LmtM3l/n9ipBFpgnUaUfIJE9Iiw5hGI54+F3K6Sl63ePTdoPEckogQkRxfD4
NaJyJeIUjfIjOjJlKEk0CeH8eQGNh+Wt4TiktF3RhjWwAVCDjFXLJnCC3yYvrRezDHUExykTc2Te
HxBLM1JC4zCuPzrg7RJFpeC2P3y5zmx+5d8s64mxu+CwO7yRY6qoGsbWmf8fN5EKiE0zCivZ7tuq
5amsLxnvIIlHpmTHcYLsp2TR53TXp14b9l2pdnCW/hsngbl1TOWjDCVMuqMbBEtZ1GFOYaSQndWh
FTY0ixWFookF+vr0hMgX5xAUKMQ4NAZgrKZEz4myU+SFAKhMv14eXhaKfibkX0135/U+wu416/6X
4rJKHsKnb4Y0iIuurk84jOsb0JIOR+gXd+CCAiM0iW6fXDhmAKt5k1AqQqQlhHr6ASdrYc1IGngs
Kk8n1gVE8cujNrSeWZXA9a4w94fUQ6oSaBSAu1wt+Ce/rp2G33x/MMIdCf0IVVkt29rFw5Loy3re
IRMnT6OyuU78uk4h3aCALK8ue2mNCCJggarmGIPhv7U9xo+Br5UMHBUEk8WOlQGZunoyn6Cz1rCo
8zB0IqI26mL5of8y+MB8o+uN48AKOQ1g6N6kdFS2fU7wVuW473j7SYKk8zchXgfMceqFYqT6RIuS
m8fmR54rhOY7z+7L0Pc2gqOM5HnFQuJjQno7/XxNsCe3eap5HVx64jwTHJrVmxAptA8u1M037iKr
XyGbg+DDUfpjiD1udvWxIVho0ZbJ/mDpnuVEzpKbrY9jI0+T8Aq8SW+06Omn3hMEQdAZo8KxMxHJ
IQKG3y0Me/JFJ8VBj4qn43oyfZuZX6HhSx9nmTPgKyVeU8UdDcKyQQ20Pg+Fi+45kTdt8OQ2ypDG
t0pDbsXavq8ybLuWsTStSNFSB9/Kp9r8gmzJNvOBLYu1xpjCFkuf2aNbEBiD4hfGphDFgpQ6N3DO
6FztV592/E0bBkjj3c1UWEFIYXjnMH7uqXwbaJTsKHFHK8IQRFU513YtF0J4dgF8bfvZx6XwzC8p
n5ZchtXRjzD2cPT/DQcWrf6uYOR2wt8EgwWX0GsjVYO8m8Iz5cw4I0RvP0xrk76bpEuUzzvoJWz9
x0guKJz4EHWwGuO7g/a1x538OqHJ2zxYyLYJVJrPQFFIrFVRGoFxbBT7pmr+wzD5ornzEc/u2sib
rc63Ow8JFzgK3dwNfHVGIverKDqoKTUKIWyuOw6z1n/mxG4ivta95ixGoBQ+mPG9grZAW5mIODdT
U7agLBBB0SyqBDsiR7vdSni3gppANemVp84aYKDcfwxaFn8TktLetOI2dmKVlwA7uBo0fYBxDfAV
lFyPNwJobA9rN1P2Q8NGks4TdrSFuO89UrpNY7YmHD2T2LqoDiKaNFC3CP2R7NcUCGUQLQamt5ut
mmRrx9roNXkh+re/zSJGEzgJ7Fsg/oEWbN30S1aACTMA2E9idWc44FKAU9nBdfQR7NN5VqaczLfz
PF1EsCiaGKRJLNlhP3n1EFwnqOyFJGO6C6XnUJG/OamTRV9YzNYJnJOtht3MHKo6DG2JPA+IYrnn
AaYQEZJonJtpt/QQAgdb4D9lcLbu1xwmGoZNMf1UCNJaCx2+Ax6blAw/d8aX3aXYrRvK26oSsfuE
58Yfp1+t1/sMiKjOokpvwnzUZZoZ6JukWvALlSoMln3S4oqxD1vjKMjNbiFSnfTQbEdrL7N/TxZW
w4sel7x+Xz8Y38Qj6HDMEwnzua9Zz+4d5dZx1hIq9uiSaunwtiEIgEoXs2oyTxKmOokyQ8zU4YhQ
3ybEfXsjWVeDJdV87OObMFkUTylrz40YkhL4HUYP2QSY7/Kgc5SVYP1eTt5FwxqVMRUgOQwvxbG/
nNOgL+bGUZl8yL+XYiimxvel3EU4crzLdavkgVJadeJbV+5Hafnxg0YBzrI/awKvsy4XzWiaPImc
7mzUnsMQnDf7tzHYoX8xbIqrB7KQpJ4oW45kv0jTYP/Bq0rh7qZoDaKE/Qsqw/lE+0tZ9XazNSXS
3RL8NULzkO64vMHFxGbRa5NYHsNDm2sN01gpdhgUQ3bVyHh81Q8ncBQe8cywWrRJbgc+a4yNfmMm
rjN6kvs7OxfQX7ZikNCzKhXTnNg4OQS8c+cdDCtzlHfuM0fFa/oMv8MGD1Cji/GfAnUvOzySSflB
Ydu146PhVMnOZQVJhqTpsDOk5GNrJklOLhbAL5XSSUclSLkk2rVJoqqdlnFIbQ/Ttz1ck4uvADsH
0PZqOCDiX27o+Xc7qV8eVT4IlNf1F4v0J6y+oa+DjR8/qH/O/PKv27Yi0W76D/0idX+S6um66McZ
t7BaB7iZOy9hv3KT7O7DdauyLWuyaE0Q4FM/YesFFDa5IWSDGLJtoTz3i4m9ooCR/VOXXFjQ3bB7
7Q9d6KyVT5ez95/xEpKdRi4OoUaa7SB74niW/OG/NzsT6uMvkqTJhfXKvQ4YJWwuhi9dpeEtRL0o
e4Jr/5VO2HZcwyIT03CT4UPeJhjPrUD2fQXjj6okVmCmdfwyTTF+d5TOTUDPy7dt+ICiq8fgwc7q
00ZvDv248M6EoK0w8vYhveD7NJG08SSM/MleCLOvlEtI1rPgScN2cw5Rn3aC9QB31E3RwsKN6l/B
KEcyna7o4ToA1IVi5syL37AGKuMa50BKR4ZtEb8xyM5FDoTSH7QxsvFvamSV9/+707boO5PG/g9i
dvX784a/dA7rUT3i5FhJqgIfqOcot0v0tDnopchuoZZoIcdVvzMjFTCmsle/2boxAUi0BkDG9UpZ
tjxvC75PC2rcE4oPrCgJrpF7F0dlDDFnZPpjGvpZenboMMICdEz5vD29TBsTbrPKWRIY4XzyGL42
7XOgs4NHuq7jF1uBKwT5iuFKuGwP1vafSboJhjbMqqtvBnVHhTxAKqI9AnbpnMcSbezNVE9RHvsS
J+G/UBUvnBne2bVz+jf24c2wSVbEiQFNb/ZLgrHnQ4yS1lobf5pYQnnfSGNZdWrdkddeDzcd50A6
jNw3eaFffbkY9WbENLUfV4i0GcQZdVIqvsP4y0x6EiLlktRXgbJ7Bx9SmqDZRnPC6nzK/FKnMYYL
gfiEDlsQIqJL69CO62fzfer0ZLpc8HD3zqf4VX+wWT9PKWrroSr34UWeihgbBiIo6spNmn7ej0iX
BV0/2V09vMXuKTL5eUGzQHuKkUZvMyiRwjCr2SCy4u9IlaSDABS8uPm7e97a2D+HNyblrYN52/Mw
GwJjEIHzO92wLWFAabZDxbtUQ6JQrwnIu5Nwha5v1Ji5ZW7SizEgr2nMwb0kkQku3o8f+LIlJsik
u1C5kjBpspi1FEE+b70EWulCxgbwNUw6vcvUrD0OhHgwNS0+RO8jFLG709rY0SzlssoetWAtgmk4
Q83QqCx2ZMOMDI6vl3wvUNTgMTLrRafiKndshfUE7Zk3zEYdRjudEwOcnkuh81akyrhel3JT7rln
nMRIyYe5bviS9YdwODpBU1lTEE5F8razDOTKPk2yQ6vmmoEUXt/NSbnAGF91+u1I35pheyRFbgKN
QGomHCrwDSMnrtqVnjUO5AUCz5r9Pc7INyVqtf1sw1UAMVZpdOkVdUpKyR8pW3mMJRGpRqsQRj4a
VU7Z36lVKx/ly0EUia4zs2tU3LHeToRndJMAuFoVahc7Q4mCBpLRir4IEJTogRYuq3G+4/ZiurYr
tinVJF2nrHln2IYD6SKBAbgWlUth/mg3Iht8Bwv1yjr2dPQGlTQ5LBPTh5Ya0LAOsdx3tyCr4p8H
mQIKNBUKg1cqzpOhqeS9AfZ2adwrWcoMp3IJ4wXP40kh+YF8MEX139wQxSiQmjoSnCHhA/Wa2lmT
w3j14/IhKn7tpADsCTlm5u0xEeUS1Pu951coNfUl0TB9OP0euRnCBxeAO9DVxTYvXPkHBCiOyzjM
RbxPzq7AYxtmFQ1ViZQbuRjVb0iMN7UYvMcyvqob71XUxWdXe5+Qowk03ciijOx0vimCiZ6Q35Fu
8D5N6XIQ4h4o14XCqjE6w6eTEwITonzifI/fxmyMm0+z2h2D42sgMtYKEU5LPiPpaH/LKHv3vI2D
X/wwe8+XwIhWF/eW1D2DM9PLHod42NY3iquIwQVEFpsFqeH5BzGynAGr9zIwo3JUwvubFXpK0cP8
m7fLL7FO55LrTlN31jVIjAsrQ4DCRlsVOHvTf+RT6vFVQ9BYRwM6hvu07c8FxmSGugy/v32kGWgY
MXHG5CwioMYYGavY7ZmoHTrH6Mem94gUygq94s7IU0ikr5npoK+vADDaXKnbT49ca01QMQGqbOpj
l7ulzCToFOqSwxjXxdgJSahr0f0+vbY1i/hlDy2FQ/7iVASy+dGKJ9rqXEVEs4msTMt8ntDxK9/B
7VHiD2e5FLnDoCyb95lesRbjTS/t1Dmm5Icn7YTGMbzzJJIdoa30itgkvc1zTp5AX+vb/4OUl59P
CYI3h6bKR2g5wP0t7fUUqH9KneXivXnw9su9w9JbhTTciEqiBUjLP34ddOAHJKITpQ8wNYD75eSr
QmJJDCzNxr4gSXOcpxl6NhyBeTKOu/ZombNunQuYUBTNMXUlJE4/XgnSeh/G9dE0C3XMUnJ8858b
P63sj2mdHUtBCHcNZ9TUTaNmtf/FWf5DLHVkA5t/9WvXTr8qO7NII4AK61zhq81lW8ohfytRcoBa
LnYRo1kCzNoIhjRRsrjLPN3Kc+om9K+4SBDGGljZzGyLy2f347WnTQvP2ToVtH/P81ArXNXOeSMx
q21pbh8Su2qUfo4WarDxOYZ2X/NImKLniQM6H07rt1NhCPtb0m62b6gEJeLOQnVg1oZE7GralAmU
8jn8XH/fuoWW8i5i5JygDrmY1E8eZi4q6lAwQmaRHyMWIvewF2gw8L/uYDZzvFfy+KipSb+uS3Qc
mcvzhTpTVdXWq+AM3+TyiHx+2NK4p8+h6lTgzfdW17A+VR/hFbpiV+/U49DQZ5q2JklQ3dDen3Ov
uU4fY/M9lixHBSscFvaS94WA6fxh5i7zAIep89rcLJNGrg142Jjw1LZWuSgujL05Quu7dZZZqXYd
Gs3bK0Imd6IvQ+mU9fhFrhFlg6mNFERJhsc/+x8fkUWBTFmsO2rm9zDsyZt1HPL9RoDHSFKxck44
r+RR3ywp47utup29jFyVNgk+Rz44ESKEc9Oyoq4PaBwHRJKQIZbfxSz5uIaRE/mKsM9PFK+8M6rv
GsO83WealyeZ7WOOqYCaUXeuEi8ddtxL4A370EvVDJeHHTJAbrmOO8FsxvJGehOs5UBSUiQtaKSh
Df2EkR8oayI29K0XcknnR7Tg3EYQcfd0MFAveALv44ixZ/9Ft0ZxJqtF0kpfsxFivcwawiDkEOF2
FmHM0NTl7g8EYitNK3LhICskF5IRmHdPZ8b5xXhNTwP/eFwtxt+vUkbz4izK0SLFmkY2FSKf+HRi
pY4QVr/RIE9ajIbpLdWFizFEbRUHd7WHerkuz+ZcqHIjVCS6wY+Nk4Wf014fBeMGSb/dLHzcaPAc
hg6U8dLZxrTz7UIRB5SdMQXoeeEqRhcpq8FkgQy2Z0B6DWsI33ZSMRg1OuL6sPHWgkC04xaWtNz1
DGDrWmpZIvPb0kzpobTCNu32AVKR2/U7T2tcscE9h+LST2emmGOFDd1bN+HPMIMPYSDWy8IVq8ex
eyUcBP/7dRHhwkwdGOY+Y1FMw41L46w1nr1PuR2jU+O9y9BKwzzcJSmz7tIyEH8J91CO8qPWcc5q
IF1auaP/5suy0JD6cA4Xlp7AcyNnPIouPcItJOLKLgpVijrQGjA3n1opTx032nOlRSqmypP1FRG5
oMd8jwb8ZyzHBPw5XlKVtTCUxPR0VgHYsnFYDQDFRsq8UyfwJb5Pam7DN3uNQrCZ2hAOzEtPoGB2
/e13NhorAzag7/WW5VJaY+FidilbyXW4xGmwqf3fKeXYElJg8A4DkNv5mtWIjJcibNQloySFPSJE
uZoOyI/hcNZj/bGLnQuwX/m+tZCsh55ZvyfZWxL1aCFR5aG2J1FNFkz8CgJoEdkWpvn8kx4Sl5q1
4pgOyl2+YfBok8eB5Ke9VvkwpUX9DVq1oNZ441aVGZBiPQMe4JjwlK8Fnl8IiY74QjNZ9qhuyZkj
iM7H5FHm2ys7OujQfzS+loN/eIMXdup4VFy6P5PMymQJn6Wp9AE8BtA1n1cb4v+ZoWwaw26n3rMC
vhBnrVuQ5Y2d895P0+yvmX0b/DJA2NMQuTzUChDEkYv7iRq53JAd/UyF9LPStPOVy1VZnOM0yzTx
USFdrXclQuzP9oajY49+QhQ4akBYbNEpOdt7yf/KUVIsH84AMa18vdionnvy3CpTapIKxqtXc15U
/U+2tZwCc1C6w6QRq+60koLAaRVhX7uif9RulGvcnRphm82375S0nVi6P4t24TaAsGXFW+U1EVta
vJ5T6w93UUCyPw2TnGTIA09nKKXrdIcdLqzUS8TnvfDoeS1wlsKly8pGdIy0jSyuRiFBCP8b+ImF
uWeBDsvUG+itN9k4jjjj7jI0af3wneo9mDo8qcYDSBMwMgS2NwDuuBwanrGumwvQXa3QswFAzEF1
U5DxkqgYNDDLsDM8x+kco5JNtg267kRlOPvniVd5K2Cm9+9FR9ogN8N0vfYQJkOLbyZafYF4N+Gx
gv4RGH8o6dqFkykXkoqai2M5cySCRcsmvbuy0BfFU23dCkK+uaR37gkQmEalMQQLAgbSMvfTOvlv
xbWIjuoCuKi13JYGXT8pnzCuN56JWB+oOxUEWqPP5PVSDQMIxdh1NRheQa3qL1BzSDVWGHR2/Cac
vVgZPwayTpePkExJOTyrL/G1xzfMCvWCsdISqOhuVVnAipppgL8WJNpeIz6wTbz7mhN/anLqh2cb
RjcQ6p+NvyUJ0XvrP/LEQ2rBjamK+hp09sbfeP2C0Df6eu6t7BKk3ugvYpOH8l7ERE/B9OfHJErR
Wtt8yp/l0Hnlcxslxp5RQmZzXIFKfLDBxG5K327usZhpQgiNJxFKUYeLjt+bfHjvGFJp+Mgl3Z8S
JcDu+nEoyloYBgLzfxTFajt4JQpJf7BCerC7RebGOOTiYcqaC3sAQksB5w9YSNfbePhFO/FmfjTV
53NOFZcsXK+juljKLvt8AiATLLTHYW4vsW/iYvL8LOEjzJWBdYaXitYlhcD5pq/V9XjLBNp95/8O
yvi288Q8t6M8qJezNEmqn4Tb0LhBrFPGSXTb0o3xDt7M3ZvRqrwu2CJ5pgOcrsdN3irxVqJ2Q8EU
6UXJsyq24O2P2+mGYMm0ang2gRR/vn96WiH4XxJRFGsjhMCbqtKy94vJj0gPLvk92By+EoxYGJ9L
d4u0oFgG1X3NKaRXnShPgX/UjvO/iDDtwCpVRyltFMOLVkH2/dMe+pBA8LObSAt57cmn8JUSKbE8
XF4tz849g61AT5PZjbQtoai6aLELx+vNLIEX9Ae1UP/U0p4Na4bghLmwxMlBrdR9GADUSRb6KRKf
sG+OTXxrLdL66P6ruOYURjYLht977o7bDWwU4naca4OIRq2L0i3qlqwbuO8t8zmWe9kjkAMZ9cjp
eOaIRSyQf/tpjrU+MszWIKlUz4Ll3i/MMKNgBqMPmyTrg/tAXX97PZCeWecATwb/wQ6bgStXjmca
m79h+oI9pFx5WvFswh43HOSgElJRQ4AnNku/rppwX9iMPK0jL8K3DdLlmE+fFR7h/CEjSH/5SKXH
5EtuIuUd0ofzPbF5jYYajbXZVj3T2v1qH/QYQ1n/2xQ/s9uLU9KYRPNtovqRejNFEn/Wat5gS3t7
aZuynsSQFQu4EjHn+qBf5gWH1ZXjP+zP7dkAJZFjrgacnczfvSVo3ojZZNy21pF4sWXGXxiKpUWu
XmFwnybpFN3Bd9q9yeT9em+m0Bbmsu5IU74/X3dzPrfIwDdt/a1f+OvYz7x8L3OdKNoEDiP23zQa
I9AcpKNovq4LZcibg0CP+Kz0kdv+3TGHJaIHP9mc3NZ/Ln0Xji6/aekMn5awgOo4qVnevpAeXaV9
2HczG7W6dOXhfgtSI0d+SkUS4mTWmMQTt/zxqhfKMrJNqpkzyutSauPPXBVwzaeKvTDxFA3SnOz2
pV6f7Qv2XgaIPwY0r27Qr2fjdKI1/VQxJLJLrG9n2+e9lSPF5YtgAg/F2RraF/6fC9iUPJcbJHRH
LtTp0DlgdbemIT8eH47p53oyMO8v8lRIxaoFjyeiE7zj2iFfPDQ8lkAXYYy2SZk8rc+Noo6Lty/Y
L0Ur3klSJYniopmB2VY5ibaJJcKYCmA1Zv4Ai9giAK1ye4uFERllpYJbPVfb502SgYGP7rp8YWsg
A+VehhNyzO1xtY+vyDgvNOX1LWl2N+MP7qgUmmhDXGqITF393MdkFIco87lf0QDORx7lYBPhJKuz
1XDEnUCQXhm0cG9HXbR/pCsKNGfkBHjYtvFWYV26XpFb7ael01UQ4VyE43mFS9SrwfJH7orZa6R6
s1TL8pLOuk4ou9SwcyJPy2Dc6qNF2thTwbl70RgH5ItD75NrKltyEvXjjv1Vn0XuvQpcG+IFSSCw
kGHz7KXx14L6hwBDF4QJ85hcgVFHegZvTmimdZ23rR0t9wNrUGZWhC4m+Cv3jxZPm/ahP3q3Otge
a1qib4YSTkZPPTwa438GwVkw36UYyWyVQoVg6V5GRIyleafR6yuZd+v2JEgRuYCBXE0wPcFYoEyz
CdWhhcB6dcq8Qi7ugiBGWrXTRuXJOGLg9/OuHuGTB9aTzcysCPgWofiTnJtP0/u7iZlO8he61UFx
dxgzJ2bcpHCdD+UkbhELx4SLnOSwW2ZO79RIVEpr8Jz8MQ7bA9PZjnHSaB8sRHfkiDDQx0K2fOue
IWvWsfublTuYne5UjjLsPmFWsDFfTKUwImD0UO2SosSXVCC7VsApjNqEI2e0E6/rSmWXfiODMZX5
BjK7MJoJ9BipsOj3vjLfYI2lSVOkCENSxOTclyYt/L9l+T/NZVBe62aZ9AOAIJMScmMP0Ks3GwyI
Ne0dIt7bE80nUi1MmTtCYhj25eaP2LTH+2P1HIbMhbvWe0zqU8v6fXigfVi0sHBBF+PYPjEaRY3I
Xra3En/8fKbZ1YVfV/M5xhIMDV92DAPuqGYb6ehEW0tZvR3OaniGt9RPsIMjkeJC2berveJICnGz
7Xf/svaEkp7yYPSsE2v2E7WdwVz4rsd7mI+nNu9G+K30QLQigvoSyMA7piVIAhgUpdTIth38MVxA
Pg0vuNXvP7Ty1+OJdR0iwGrEXkX4Dq4VkmhuMGA2IyyZgwVA9AMxCYf3F/7zT2rnvNiJY7oFXF42
wSpvje3nDBT2puLGEWB05hgKbsMt9/x6Y/dFukQoF9eEyeWSILGEPjIt17C2cKVGe+zUVOoc3SLh
5jmO/nuxnroLDt+oUcXlji5uX0asC8WIHpzKCbrJgyJU1aPTpNq+Jnsvg4ZgzaVcFueHOazEjkfu
RItcphv7Lr/ngLS/H09IHdkjOfJAZHL8IM/Yc3UpgYi2Nhb/+jys/oMCNzEMn1rTWn9Uc1tfHSUn
NTd+c7eynCIPR5+j79pywJKTX+gpAvbu7i06namdsH0bz1amn40iF16TFcpoonOztIqOwl3iMFEO
nUrnNYusVUc2OSdw9ZZnZLyvSF6j5CiPbmhkZtwhk14WI1VS+o1OUvcKQ64SZv8ZBFLfeLb8356u
EM1xtEYwsxC/VSIROj07Xp6YFqKQj9HyhLMlZe5KqegQeajEw8GC8SDCdrn9WuBtNBULlcppzf4M
ocJ3At580V+ZSkWB50Asvyw5unwpPh5PCmm4v+Ttjyu/uyJyIKQyUCV+boVuJFdsOXmaAAWFhu8f
DltwE2qN8gKR/DMVXtz6m8miHQsQXt13AASO+UZAKNE9MIbQO4LeMZ+XO7xD2vpvF1c9G3O8oZI7
Ed/tdkdNTr4y5cvd1qmoQUVfWl7jDite+1n18kkPuDJ9pdxomQO3GIxx15nJj999ZwzFusSNLBVW
P6PcwBPKplBHFEtR7l/sAnc2HcvPL1dPdc0odSBoQOqzU2JYrfJYHBY+eLWeNc55qn4PIVCXCFgg
zECi64a3llgFg+Y22+UKXJiBnRXTadxqc7o7ZZ6RAm7j0pGEh2YiFhhEnnNyBTgQdgRu544Gr9Rt
K8+OOgVflIhAQMppQUxepjpah3gMq4fhust8BDYv+7Ml+snO7jSdIjkVtQcmpFFbZwaxFPhIcG9p
GBnpLdJxtkjTAi8mGMfjaShY0CdxMQy6JpPEdBEL4TOnQ3KZW3cgaC4N0tkBU/lkFlbXwIDlaTbY
GjQGj3aWHeGY18d+9IP0DCIc6Tlnun/cuZCpr3x5kYpkb14UnIfszeMhKdv4o3j4ZoLW0vZZ2VHm
643GHNXCTg8hG6kRvx3rdMrE6kGuvOhXVd5r5BNahDugA/lbtgk/3kj4NYFdUgzKEEjdNq2RXo8s
bPPz52HbyesWo2nGy4m3LyxJqahPsqNifIt5iZkvyhWKJrsAN5TrGQEhS3U2dYDz8vH0bswMAsG1
inPEUYTRtDQvOYngWdthyb4fbzQ0k+malicPwndi3MBLD3HpP+uZwMzRUGcBD+n7FtIq1YDQWiRe
V/vJfj8BOJZEnxO/vtxWVkC+QuapO2Lan9DaJbaA0CR9rVgn2jE+DaG8zLrLjz3bXmvnNUuuSoGO
0ZF0Ffl8fR24BQ8F1xlJ6SczXftMfi63QTy/5coIeyb48/rw+PmFYFb//aOmkWaKaSOViF0kUOWJ
UGEX9zkjemSXVUne9QuLW6dfM3s8ahC9Tn36HXdmlYGROc4+bxpp2fng+ptLL4/1u1G46pRk/2O3
C2yzdS0AEVF2Ahh47jU3yMtVPYmJSvl53Gtllgy/TsQ5XpOM/XuDIOuqYwUFD1zBENZPZWbg0Byn
BZyNKvVyNR31VRDR8VeoJh3xldP9jE+rc7WzDpusiGL+yExJyjdAJW0LZ9YIM8yIDeUVUerDRJdT
RktzCivItj8AHiKDHB1OND/tTBWF3AuIsKCp0ZXzg9SG7LjKCyPdOEG233CyaEmYOvxmIDaZzbhU
DgJaZAkfEggtsJze+GAtqyU18RxcjHrrWehVRt6XCdbQWkiNG+2kN1j4zA8gyIr+LCU/WU3sNcqm
Ema+YPEyJ47nZOPCR6WHYq1RhiLCZYjeTWkA4GNlBq+frzwNV9K3CdBF6+XKv4P2+Y2+fmxiJQsz
D/G8B7M/5QbSyJCra+bMVlbC/1dxWSJnUXZ5DRIwcsAdk1EduG5rQD3dAsBVJuzF+FhcdgyMMeel
sW8hFDXm8ICWpt2tkdFJTvpJL0pjaHlWslJJrUsr3dt67SJIoC/mtbS3ReyrD5L067D1NlLPihDM
X85z/zmU6DbK93xJco75xa2OzVwpYt1OuZKrdqWHPL2Djn1ac01eJcbhzEJdF0AC3kevmBai06iM
xUJiGHAb8xlT16D8WQfis+E48vNLZnDn1op9MaSrxmFhmTcGw8js9QKj4heJz3AqEcDenoaKdpc1
OpDEHSO+LM02Tp8IDcKuofg+93qZ79RxYvI4dAvU1hmzd1JfhIc0qTAvbppyWmHLp010w28gK79B
4iVKGLvZhh4rZ25ER1lhZhhLIctAuqIhR8FQxGjMxr/pqEdXsOVi2AnsNiZMfunaEBr1cgXpzli3
AhMgSyUPZ3wz+Hqi9KebuSXZdmflZT0wFQVg6BfTT85tFerXtnlxMiKbuqL3145lqO95CxzWCXil
IsUZXxS/FGzuslxCWA0zlzXHS9A0A7RzFxX+4YLhSmSX12AoFk9ILdKK5cam/Fjv5gGqJfDKajkl
PzigiczQiod72/fN6WUNVL3LO7+T8ydAOfRPKGj/L6FrkwdvhXptjsaVgN0AgQxJFN8Yygq4HfAE
1ZkEqjWr/CePApaVG8s77w+SM1cOdVriHDACgnNFDZDEOBi0hZyVU/Ttnl4sdLZwdoAvECt+leiP
APAAV7DYY+t3PLdz6EgLlT6axbY0OjWRPnopfJlfoJH9TzXVJ5zH1Fa6aTrIDvVqBZJeXRJCwi9c
cIjxC1f0qiTB24n2cpoq4kJx9gz5toflG/DkfokUybYJb9IlXJ1+yDIBS1vsZFCSLGoxkz8TA05X
5/gucU+nBoB3Z6u5oo7HsCdvUgChyT2xuXcnVnWKQGFvKWDlOuMEDTqbDWc17YdrwS1rDnvFr3eU
ptfZqZhcbdluxm4msJFEnH4FiYu1zv1FwMag+s/J5R8/aMzumbOLCQf6oi2nvvrBoixf505Vuqwf
ANJ9HhRG+V2ge2RSiCwfzUANnZr4wY5ztYt0+vw11hqDqeN4IG6KfDS/9W5hGyqP+pIZPBuTs+kj
fPMmPAUVSwgX7jXZcqnOBuwSfSWouaR35cwNE6xDLwsNzSEjyGRQ3QkTfzBNlwY0QmakoMWKYg/+
kfzPa0hkYiKZE0rIl0rtHEGzG70e1NxeTMahdxcbtoYvRNM/uM1V07sXJDBM3H3dcxjq0qMyzhjn
9xrYsGp8hP3y5AMf643yNZFzOWxLu2QIRQWHwlk/FMNappu0GzVEN/nBn/sMIt+CYLemX4nqv8fg
yToJQMY9GIRNcjEMJjeAXaRanNgqPg1CNJ5vKC6JyOJjfr43P58v8BJMWW5w0doSkRk4s+hwjU2W
UAU6/xIB+m9kVC7/RIIsVAX2UQQL/vyGcCuV4DKfUiOlKLWEwW3SKX/pkikpBnONVdTYm64ujU+i
mVJrpiSnNBTruK8nh3Yqo05ESd7SiDB/3m0PUVXCcTB224Zh3NSpuqhZ0+mWCZNl/+pdQyOzMWxb
GWcJLv1B1V9C0MPpeEPhk8SfUv2Or7HkvfQKbASfdcC6tt7uhXt2pGfrppaawNqpsm7HNXxadK0F
UsrxjHmM0JwrzUfwL8cNKNW2UUtF/jtItJw/UFWpzorXN93yR/XFioVZf5zDKGhf7drOrYppUFp3
gughpWYDCqNm3iRjphuv4Nvcfb0GFN/CcNnSdq75SuQHfNrEwsNQwjUVL57V3ATtjEXWAboBX/Om
A9srWRt41jPi859Ubhdw0rfUr093j3UqGyHHsV72j3L5kwW/nR14aQWcB61fSLuW1lHA4oKL+SZK
01O/DLwAxpwGmeDipwYPNdbO1GDylOovnGVR6ts4GJmNU9k6RLxqTCqopU9Kq2C4/UonollZctZB
wrcWkQDpxkuQQfJx0GnEP5WK8iXhWNqkPIyJvODm0wVSzWVO8I9H37tRTfaUf7pUyxnSeqQkMGsY
65jF5QctJTk0VcJiJUossgEoHK3El5VrgIa/YL+HN4WWSo4lE6gDrAMv/+TTqck2G3uSj8UvEA9h
aRNygV3CqjvWBThWXcu03fFwu4R/Ik1oKTf6RpIL+4HvBK84D5xC/nHVPigMLgkKH6XqN1ZFHhjC
kAIj3VjwzDjpcVcfH184KFFELWOukVKmqndG0A3yPIuO41NaSxxoriEjacUp/Skpe0JSAaXZzOi7
5PBk8siTRJBaTMlN7vrhrxASrVwCKL/lIzWwSKB6v8fGIPU511wkj1pEMwJJeotemtoB5eHrRzgd
BLkIdJb5Y5e75+B2VIf0JZasItKlIiW1MBH91sam+okslcRyZMhZC6cLhv7zngr0t+HT6M1c6+el
vWOTBAQi74GhM8eeEsZ2aq+yXcPlPCmP/etrkNtbz1IyurBqVYvG/D9irWQfgyu17pZGpql22IaY
LIDbEQt4ZwBS4uWIwEl4MsIHzRrCtfTMWxuawbZGtmN7+caS8c78zTPsAg+1TQ1HP27uAhfzvDwy
OK9KxtmRlJWneaTTA6UfamQ6WlxHmRopHSvst35MBtd1M3VfcSvWBjRDmcH78yi6Peqhx3oscQMo
75qt+ppe9VQXXKfKveHbtwrifL7IPzMF/xL9Pynx5d1MOqpbi6QYY33Ogr8/VQZxGTmpEEBLvE2P
GVzpBAwCul+zz0c0YiOj2tO0sEdpZWftMe93umC60lU2mcpDfetlyEjbYZhspxZMmQmYvFGbBbDO
+OOGlHHD+BwTO73JwHWQBefdHCM35643n865YFLDQpwnt+773Mm/yQrlWcyUFXDQOBj08H4uyaAR
Fs8wqavJ7znBZ2N68mjtwn4mkZY/vWGAmBwtD5HIaoGKkzx5HFtX8t8WdcaNc4UVO5ICzLA5fIVj
oQ76Q5lUk/kzztCKlgWRZTOVpYr/qjPezsKneOhNc981m6bryGnOIit6NSpyygxCgCL3hdkorfVA
zqAU3V1EQb/IjqVaWmAY3FzAZBBdkfYvi+xFnOxJmiIfegwYBYZYZX87slDJv6FsWlpcaALR2j4X
cIjDfn4s7hDRo24LtC2ug6LBFdMSeiFP51UMBiARsIidonTKw5/BNFRIIEup0urQb2Xo2L24U0fO
yKPtmbhvu1aMu6ICQMVrNxddU0tZbpxiLDC/KP0Y6l4wCkwz1V4GjCMpUXfWuD1lJYp0DaF9Q8du
hfPkq8ZjEzLW0/xPdHMF/pMxKIVwQ4taxTpzzvk1z5BZCqaHS3hpEhHSGTamTY1DbwMrbYWcZpyO
3lCu23CVD4j9fpwCXAxNPTxgxY+k9RIYF13oSlrZWshoxDhP20AbINATyN5lzJNsV4qb55HfKRgH
KuIqNksY419vcUnmhzGFKcuG/SUWAXIB13Qi5BQ/lrs4BVylDCBxNWi5YhDkRWX44Mb9orx8+z+2
PgDg3MrJaxwq0mUclrNf1c3YtkiEE7XycQq02fUpKrZn+hqt5vQYrR4uuEkl6efkMRaRK9GUZP3v
aN9qd53226TOxs5wTBki3/7RSyyKUsxAjTtQ7b6ERVq2M0ubZoUjuBtjTxgMrnmgBHIrDHqiTbay
tDMxmLuXy4bZsoUQfsccrtSeJentXQRJRDrbjUxjYYXmIJIeGllkyMUxcidsze6n+Sbtnfm5aazO
fcLftY/o0bp9JhkRmmkYzLbIH1VSYfWl6XjAM5Ynk/dixNntL/xqpFnYAQySF+Q13ryFSDupwhM2
Oq4QpyepjXEeSfI4ZMJF1ImTCnZ8oqr9K8QdlXM5W2zB+210DvphThMSjOc79FioUcb3S8wYQUFp
/De8t/w2R8kn1UT9CdRkhTw4siLyU1X17E2pVn67abMYOe8dqtYyaHDmDjD4O7xuvmuRfwb6Ftq0
n7JCfHXC/eM6wyHxNvCV7j0A2CKGGGrh9ecczBI3zJ7+LSyEOXMe1vPGocfDk0xjGksHPzm22SEa
dpQC37FQI2Ac+rTMTlr1HAgxssGh1UGaw+NuM4J6RMs/w96XTjHSD22jajL1PGlZC9j32vNtJrUM
oLDxHO9D0WNV0egLThUVW/Uq2gUMgnk9RNJaRwb8tyABEZucDrVbAnrnyq2Ia8XViejkVdXIY9RB
84BDjXCJu34iFlvKBzEZ3Vhc5QKSNKCKCoq4WTYk2TEqgQ3S3NXVMznBQWUul1JBo9zavvD8FAnD
TxdhxSR+za3XTea6MoLGbb7Z2kslnhTgaMmsG0SRPVzjWoNwqPqGLAIXqzCPD9yftZz//q7D0HuT
hiZRHX+y12fW+7HPcSHzsu4vbIjIWriSMtS5U1i/MnSZ/Lpo7b97sipw23KQTJQyC1M8AOGSPUlg
ZOe0xR3ywvBwfco0HvAeByi75pws16NMXHZK05UwImoXAPZFQhAUDpjD2lGl5VUyon3Yz5DjldaH
ptnRwurTOdH3DZHcknHIgyK11H02ZeMwuybn9oaWU7ptolusMO3cKhf9VxaP8VC+EOfWSkdXEmWj
4ZsWy599ovUqUx+0pGJ3lJolKKRUwkPSoNA4xW+bq0xoqthzuIio0iSQ3nTDPBN25SvncxlM0o3J
BVU+8cFMrm3AvzJHB1xTohLxadxi8cS3SWLQ+HRRGhlOiQPPyqJ8AJqG/1MARMr4ic6DP5HRBxZv
T/0YUOkSmJe8u+6zuZXadA+gIpRSjLv+EVPmQ3WtUx6yr8q0B75IvHj1tyn7vAYDyuZfTlBmV2bg
pHGoeUaYS1mBtXOg42PBx6GQI2yFUwW8CzwEhkMHsCIW2dX9/36MLQsTOvXrqFnEOb1ibifvQGmd
s8ObKnOHgD+UI36L1cSY6W7kJntk6Z8QptpEADFa9dBR2CjOOW+/4PgUukUCNCpGQAabcNv3iOzT
EVd9cV6W9fC/mDw/IzMSLHWyVOVPOo8CLb9s3vtuNlnN9QfDk/IID/MzVjl4TZijQNe8vpPpDE96
1dJvTUoxIarKZ4v8h+zE84z43XMM2MG2wbj7KVo/Q9kJHhxF3EJvVn/ozJg5EnOtEqU3zMcGKPJh
HMEhSpThU//YBCmc2sbSN8rfiARv/RCRM8h7Nt5Rx3jHdDPrr2vpaLOp3dpeKgeIPPgT03zPftdP
XGlFC3+Q/xLRZPTbRRYwfJOHUS0bBQurj65h+yYjwtOSMEZCxnohyzIbG3h61668+lVdU1q0MJZR
eUbx6xADlCmnFPCOPTOeruQ2yB3KpnEEsA83UL6LAlrA4bVcWAwD8T7eSoDIvKRjLkDdOJ8WT0NH
nr646xzxherTHphRgTxGdftxKiHZpIv2DBWOkMiV3lo7JTQ9Z5y7e65K8bZ1j9/SXQIgq788aUhw
hS52gAolOc3trutUnc8Q2jXTaLfgTE8O/BJjM850n0fRJRs34sWUrqaclVNt2Pxm5Qt59RH4Hzsp
/9zGAAZOgkDWump1czQu49PJexgYOSvhGcLaTJfsouJxG1kPQJdy+Glv/mj3fhKKbo5zikUrc2bC
pmpAmKLmwGr4PD6iX6GbUEE6zfB4j2S8vD8bbp/3G5WmvMn5gs1hvamxVNwMSKoB6GqnwjYDXgA6
0VYaGPaHnPyE0nZH2dXTRj5pR1+vJNLGbTPMLOHglj+/HihMfH0/R60aWnWnMmPDDnND4RWK8UmE
VGKQHPrYz47vjNVGGwN1c0OQqXSXo+s9g+NmJOMFzvS0FFi65f37yomDZnQ41nCkrrLfx3KzTTMF
0HDIw9bb5bInZlKpegnTvCaUCYXi+F4A64Btffx/8gWZhA0uRv1wuv8CWF0LdM7F1o9OAa9MsRe9
TMKbfqrga1MABB3afqF8tQ4n1EpnX3GeJ4y7Vy/Jd57yigJjN/QT91Q+2LTrk09yf5keNoGdBkxw
ubTSrZ28dWKjAYhcbAU958r0q1rBrcDYVIuufQ5hx7uzD31npLb10tZZcPEbWP5olVgbHng3ZJNb
3RlwiuVpLWUMpy74JpzflC+0zqbASdaC88feIM9r3FWb6D9uH6vB9Podfi2MiTCdiEkfU9Fbcljl
iJWX3QGAdd93rJcemFqwdB1l3tOGCH1hWX6Z7r6Et33hk59TErgZ8fixcqA304TyqsJbI3vgKbFO
Zplmt6h4rr3yaUUSdci0XQNoeYq/qIdogZ+7QnCNLhABfq7RQENgVGWNw+c2ni2E2eLhMkDTUfvy
CTfFhEgZgX0B20oC+U4MYWdwQ3CjCERx1fEivu73F2uvVVaI6umYXqA/jkWq7qXe4rPtlKW/Msur
fW4cW54jss/5fKa+F5nH8obTm+vs+OrcD3ZT6u7tHiC5amRKWDUKojgX8R8DX8xnE8fZPxL+9ohm
jVwoXUqNo6IzSxMV+20c2rxBe7OPBk1s2ivljneUmsrgB/HxQIM2cvx/LR3ucsdZnbZ6dB0QpivJ
MAgretXLHL2zqiZFO0zaa2PpA4bCiszyRtx8vCqZYtUwJjYkUQaPsD/cMuVZ4eDntijzCKhnMDD7
KXZOgd1FeW65Dz7BHfG5RJBkwBqAnDRLhpXDseJLsEaq6wTau45wZPOsxCiWl28npld5zPfrL2Ie
kjxpd/3OL856A+q0Y6Cs0iv7Lomt3kC6ukGJ/NorA1EQT5JT7J4hLeg2bgBrLaESgDvXYBuIaQHY
hnY5LIOScsWs4TGTUZm6e4kpGpndKTwZVZ3jy+ZFu4QayOOUWV09b6yVgmXA+dp/tRRNWF/XK0pG
BTfQ9m+WcTvKQrZLdbHPv2jrJBHO7DA6Q+6D1+N+2rc5CGHrv+d6ZV7OtgFGgC8AiR4MjnIgpjVi
B6/sWTjhI4Ne6KeXaTLPl2gu/0/n0YRoKjwi5snOYxWtybyr9PcLouZXB0CTuc0kkQvN7+SNP/8o
ZBLawkHHFgNNVmfbSVD8Xbv0tjzN4FkvglqaTm3X4RtfLmk4tjmMH0A9K1KC0D2fOBdl9g3/NvXI
F+wGp1Q4Oiy9R5oi9vG7lMoFRY1v5w4OI0SPQihdjMvrqQDlfNkIPvDYjR3beMqZhQF/6Ea7WQIG
X6MQDoea0A4wBIvehrNqdusnQBotO3BljYifGedQrBw6x+kvAasW3KvumlyidDUQ21I+p2/FqXci
2EtDqN0zkfUrVFbzhw2SGXjTEDrNqyF+ldWN3x+y7N0jLYYOMz57BMbAFLt/b0PY1BXqeVlsaJcD
AaKBezOLUENToW44uOvU8rFPcJyN8VAgLNk0maUxOjptvu0LcKXX2TQ2UY5c7+A3tnGBVwFu1MCa
DPPCO6y+7fQruT+nhhBe3t0g9umpDJxZUMEPAhDcvIpK0EdE+hrW03fxpNBJC+XhBCeGTpPZV3OV
apvjo582YUkEi4aIZWxVu4nPNtjAAvUqyoDYNuZtaIzLUePleB3ZLA12ayFV9Ir/5+i1bsHSX7Fh
E5zdO4AFpVXe6m5uwPA4TjlvJffVQoAdk+jYfA+GTyFdtM5olCNdqMP14nlVhBa4YHNJOYJ2fsuo
wAZb+o5ZhuxyJeAhxSTHQ2bsElQlzPAR6T6xtWU1ffeDTCEhSAkcJK28yBoW4XuYshetpt4fNniK
ZMSNr46SX6i3eVHMTsDe4MoHpfxnQJK0DLGj9vifPjdQDmD8oOrLabLR6bEH1u6D4Ee3ebefOUOQ
AQyFPE4FJs7rOHHcgtIkPyvC7tl2FBQYTJbwuTWN3EF1432Rommr61Dk+vZRB9QE925q41t1AOOZ
epWQn1Kw2q5bp7S/hoO5RUqnLtSb3pGOltQ951A3BgHqxcFopk0s/yTnBao7DMssr9MpwMSt0R1Q
5pO3fECssZbPyFSdBb4K9bMBvqsqk7JwgK5BRGmgyGbK4THFJ1ZvWe/24DFw+p/VaTP5HZ1hXKLe
mD6QuULb1K0LozGTh7T2ysaz+QKMKa9nCbu1ueQ/ekvqfbn8s787cn3EQFGa342avpOd58SSg+nV
nGyTffbnabEriI69cSaBEUE3hRb7UpjmCJEoz/I2+xCfMUUSmQtGJ23j5sGX7xlijWuCe7/ntWMm
cEtpqWMKBVhM21lD80KJHtW7BamQKE3hzR0bxEVwyK5aQiZSjwjfaJuKcTbBh8sF1j6f4kkdzYo4
zhaMnUaHyZKRq7xLNmtEsDLgaSbrHXCgDOHwcSLcngaA7vq4BrruAs09t/y8wd34EU9oGuj7zARi
XZKkSfHYU/dvn0MLeKlwnobHmFfX+c6C3+ZU49GhwOGDs7xquZKKpKMcX8NUYYGik1DlE+vr8lKs
f/1kzB1gKKMnQ7UvPvMzuoH9JaasAPXozPBJqEqZh46pIjPcrUwj+/VrQFrBwzEMDfWdt7d8YCNt
Tp8wRJ3uUiUgjW6JKnAN3Ccy6E0pRWAzNUPILxSv5/dAa9I6f+4lMumaMu8FvEhxZEYohu6ZMSWs
8p7nUcJ467FmxZ0MOmMczXEBttTVEwwXTsHlXOgCU8lQhHQ7kayJBIK7Wj+XSTXaSCldGNfnF8qF
1QEolMmSj0uRRB979RrFd52s4I586Z2jH9tiCLs+DM0uKbooiD8pW0X8umMS1n+xJLm/k/KBJRfP
zeZD1yuXuZ0+y2Ow7nc6kfn/icQowKO210PSM/P46NXKdQO+CxMSaRKoonjcD+aHqyY2WMWcClpg
CxEsCcXUtAckAnw90aR8Kdn130CYW9t1I4N98KXTkd2L5Mt3SeYvUABYiCRnVM8tLzvQ30dGgiVM
zopXMhyATxvD1caf3MG3ULXwsu9e8eyesOJPXmJFaPqZa5UKgxSV4BUSy8jpcbG5/QxtKqFOMv58
aRvffSWENbA4cMFpyCSi3Dg0zFftS+wKyNEWq7uoU1Q4lA1/4ZlDpeQv2iRHJ3u50TlUQCnYJnJm
OvXtwZMmnVmm0hu6WwJH78aroDA37dcnye6VJfKHXJ3NbOCFXQgR7ZjPq49ZPB3c/Me2Z12E5y3v
cIlWHwjZXfbzkex6ycSh9DLwVH4PovtsJEroFIqd1kbdve0jHYx6ojng3ak86dZbMeBGLnD+frKB
IZNVCoBumaOsSRyjOiT+s+z3yWDNf/Ref5jFhDF52H3OSfUubm6NTRuFJ03vwcMG3F2AA0ecJVGX
MwyTMmvrNbbBNE+8gbK3H142ZMa6hX2sW8Cf+Nogyn/fQWAQeo1NgyO/QtJD3+8PwrLQaJgYMlqu
WnIPKF2B4EvDOX4xUARmP1c00NCN6wO7nvIIEbyed85KGUwItjdytwDY2oqozezWerOtjrtpK/5+
1Grg/kkzVBtjSFvC1/PQ+0znraX79NoS9OUA/IYX4wyaEOklkt6f2Usmh+N80/z83+ycYAwdtGFv
aA8AkXKt8odm49GfaUIelNiSuvQH8gEb0kXEnFTanz0gnUL/dRwxEslHd4lmGap5ezTuWewh12/Q
blZCWSnanqKKHdMOV7fC+bxPGm5VuR9YnPSNwJ4eupX+AM2CSpjXadSr3v5bfD21e2YR4RXa7Irn
+japhEk0fvJTAH+cYJTt/Hoyi73QypRUbvGFoxCW3mv/JbRsWH/gERYUgWfzT380tREcbXDIeNt9
TNUNP2j6SlzWtU8cRV83RJiwBZEjwIEdCJnGXJRl4BjrFfYUBZV3oeF1tyUGD3gd0j54WcCwSn5a
6j50G5KMXd9VeDm+1W5q64Gi5Zo26YrZ0w19TCHw0VWWwZBPLETUd6nfhUP214hodtJeQZy4PGsj
5hs+oQYfHDzGP3dRdt96XGrrH5DGvLoiV6f82ej2RODJXrMuUiwZ+cQJ/MgdkKq2ErJ3vb4wMavM
vjgtCcXJiE3mkM0Bmn0JvwbbqlOQAv6EGz+sDdxv86QEbrhmBxhonackBmPSGedO8rtM0POMThs3
nQLN6FiRI2Ik/6gtlekj9uYe3HPimCUiDuHabHDLz31LDbNqPFPYWf4LpKCRusQjLMazppA7tXh6
0n3waRgv1GyA3cUk8VFryglzgWiS8FEVqKJ7dj7OjQRW/TOkw4K7QZiN2huJ/C9p/Ask9o4mXg7u
VADeHlIRoi80veyEWDFqkddpcHpeshTJTl0mOgMgMIweVL0l0jirYYOIOFJD4ITIt5vzy9G/KtA4
EOE1HJMJnQta4yqmpJ4zbCDqOcLB0ex45dYjWKido9xu55EBIsLMfgtNltwDJCM9iOqqZEck59/a
i2S7TvdjjZIFy9fIuRqYGKbt+mO28Fn4NNHNU3ICFHFNxt527vQ4jrF9FrE86kvAG9/BAhJ7Ndo/
bQ5asOxig7jeMa/ZHCUmyHN0PFFS4oJ4AvQIwrh5KY/e4Vbl5IORZxrvPDwLxDn4HEWB+hA5bUUZ
ySSmg3kfFQGiKGfxVDoIFTCU454bK+vlJ6MPQ3jalFRzStI8u/V9tUanFRsrcr6tuJ5bnMuxKVcS
fBmMDxp7zLj62m9bil61Kxw0R0AoJSb3qD5nTh2/1+6AYQc/10LmdB+eCZg2XcmLfIpt6fUfCyPK
wN+KDLVn/coxZ95edVuWAS7g2EY38SnPLPUJmAwPtgqhgK69YJc3JCc+JHugxFARtsJ+COggflVK
FrM/clI4YaQ948C0r2bHXcxw1KZaAqbQ9zv9d8k0J9czDVK6OWlb6DTTargU4/Ia6+TCF21iyatZ
6hbOHJK0HwYUA543ZpwHxWVOjFEU43OW5jC7Ir7dOPYGIwTyQfezLZM7vdraXtSasWiOiiyXbUq4
CPrVTRQQum1KteMoFW73UDbJvKDSdVO3Ny3E7Z3aYlsIBQVVfafUAvFw6ls1lBOUp7Ym07rFFI2s
jzubvBCFNf9Wk9YfubJeAehnIfB0tAZtBw/tYoT3MJGfsOtG67pISn08s4Q/jpU1al70xo+G8xom
nhc7RrwxYc0CZLzY6lqIiiYNS0sa7pma0cokkhzWPpeuza60LivpR1Ak9PbWUWwn9TMue2saj193
bDKOfxCa8wVBRIEL3TN2SypI4fN0W8N9tB5bjq0aLGG9c4vOYXUfKCAIGu/pnfK2lVxcY4XunD5Q
3d77DDle4Dj+5uv9Ec2Ky/FXBbLof8KL6t/9OID4FQXOE1821VP2rwBMaJmO4UHGz2GcSSCtS8YY
j3eG5z5v6cW92BJxYki9xbTE8juz9suvthjR2Mdhx6EoUEUPBbLNEf/FvAlYCpBIxzGdR/InMZN4
wP4u3TGp1kri0TL4iDoh7ZFg8KMTW6puZS4pO2/VxrrVlAEEp6gxVWrhUqP++5VIL6L0H71tZU85
o27eVXehZWb6fFhlwK5lBti/50atFMakV9hOQdDnYG8G+Ik8HUCdda7058TaYeY6pvf/e8Wa+QMf
cAiMo9nJT+NECMfyPeMtLPnGhD9NGq+Z6osrnxJn7Ir/KT324wmIFTd0g8MFA5yO/QXmsq6ScCyK
CSH7xbxa53WSb/mvvf1zg3Bru1bJehqjb+kkC2DaBBwasLugNXbDfpTPbB75VBSBSAT7fbWT6dXs
HAW0kZ8EHAyLsB+Db2O/rJZj/OE10tqN5yEWIi4dM7Qt2J16RAt44WWPAUvKszxP8Lkeu19jmy8j
ArEChqMxdgX5ntGibV3oBTokQE/pJZ09f4o5ilEq5NniI63PIDWvmIrMg2cL4Wmg+pFOWa2vJYYb
qrlTMf6QJ32asruqKl/hvl5ZMAAQALcCCCYPlSlrUas133vra1uOw1e66By9yT4jfJT2QUgAgTiq
YQojFnlKyKIrP9E0Dga8SpMAJ2Fbj7Wyi5nafR7/14+X1BweuOhj2UJVXddQGlcngi1dNMlu4gWi
3QBOEvFr0+wR0gTMfj6sn6sGccHUCNWrEKAVElB/okIAn0axZbtvSmAHvxlaJlxQDu9beGcwaSX0
VqYippzl6I4iml+o4BUidupgDt3o0DDtOjdsFuJIIxMCV8MtehzZ60owLAsG92CFw3r+mwlFFq6S
/+VXUQEOBsxacY0/07CieytTZ4EVq7AkyMCyJRaZD0/6ILgBf50R1ZGhKFo8OWqj7xkn73RoVNQJ
GVCF/O9OxudNPZ05JYY5lAfgFlxEornIvSphNWvcBVmwLC3TflwLx1FBHLkf1l+RFZ12eFFmRQCk
7nplcsyEKbK38s8owXfTL3jLC3JgTfrvm1mD/bjSIdDZD2mXwsgiienq5SVC+JntsK2H5HyTTyib
1Y5K6zRAM/8wQaeVvfOzANrR4GtxWmFfCpubwR0DyJm3jaivOER1WzOz5Suy9Iuqfa9BbD8Vlbvg
u9oao8URp3tZBaFVvTRvVa0x0NS4uuI4CR1NKuoy+jrzxv+dw7D4SYwj35UlOqP9LaDr8Y0DpUGI
Y3jyOrT7OKikbU5hA6bXYPwnI9r2rsr644HYWmC02YHEj8XdCbYyA9Zh3kZ2PWYgDFs/KNmwtlCv
zWdr1xP01ykUyEQjlklEcXz6BLoVUt4lyLsVW3wovLM6DnKCF+PsU16HUmgJvu8z9PIAUN3DyK1+
wmYtY6GvtS2CY++qYZqh1Exu2WLC5FauGaUDT1/ydMhMhzFGMoU7t/v/d5+rHX3AhZ71Ocygjhmj
0ve9XdAac91ULrwMaKv1IDvnODUN+PCGaZC2TeqAJfdco5rc2YjWY/evvUfF8QiuUQss0s8Y9bZd
ynZ+Negtn6wKHcVAtrq3P0xAMnVtQTu14qlr7Mzjf82sfwAF3aw5EzNKsz3H45vSfwoJgA0wTRRz
Jve4af+G2qyIUIqytQMlYbQCsW+ZeC5latrERjG4S9S0vZhKJpv42RFuHH0INCNAO6kuC4xdRv1u
xNERxJqivrM8hYk+mVu3SV2foC4wZXGZV1vRkSWIYFQGUDwutuDdGcy5/mXChytCPokuBQCJUd0F
jZHhXNT6LFUM68By/bZlPfN6rSIdqpdAtszvxgR+4mmqavJGkgxFa/GmRxMXvYBV8TxamdENZdEl
Woc4bGf6yLfiux5Ssirb4pWzADEaxalImvXcd1+I8KNdpvYeTRCkxB1TOm6HsFvBGU0KaJBPHH/x
1B0ornTMESOHwBCcvYQ9UqxQxg9WOu5hJzO+ap7eAbhbWzsqOAdlsHS/px1mNLTDWrlxaHe1UQzO
CfeRlG5bxYeLPPLZat//SZYfpazbI7bJ8JI0yfh/FkQDJKcdZ5Oxcr7Xjh3iYDwiMd6X14c/H6cD
tYsExQJJwnqE3J55K1aCYOrblJDhH2XgCNrdfbFX8ywasWYDbCVa/498Pd5vDVGD4Wq0yhXGLbQi
2p3vSnApvo1gtJEttG2xIDMfNAkw8vVoGhlYt6XlUqIcb85t93ehMOe7nwleaTEmjtqzXQX06jbB
LEQliuuncZVhe0esJo0GxpYr3ogx0Ef+9d4jyfXh1u600pfY+pI7UZaWwfMG5tKL/tMCCx5JPEeH
Yhh9Vu7e7ADu1OVHVhJFrx6KCvpDaUMcbihazSj5WTZv2iSflOg9zelhJZZVsnWnbcPgdX2O1mil
o7RcznX2ykBNcdKUTUuLrjo83hLj1wURWRq84/w+pV0wPEm7za+M6dGXrye33Et/NKFMLT13A88Z
nUHqLPoig0PKh7NavYPVRqufBQaH7zMo1DZJGmtRvSXqxTtW0fst/Ig0O/y6niDZkzhWP/m3anOb
wkFDEjz7bHS7eXn2DcFpUy19x836HS92otNe+w73Jt0Fn8phCK0fE5NDjMS1/3q2fm8Qk68tKot4
hy5b0MdyQ8OSfatiYBb5s2LQEfTkYfWxSQvFP2k25PKa1fA5oakr/KWlV4cR+1HXwhGw8vOJ/Kv3
sKp7GRWtMtC20tIn+10JLnJBz5sxSs4rvXzUntik+iznZalI7uYtHBaBlbc6ArH8QScFrrzLl9Zt
FoLLYczjzBW7DaEaKZPtGDEcZGdFqXSLihOn3MVmcPYUqRatSuwqkH7tqk0zX9vYatJW+X9WS4lt
0gHNrgHCd3CPPPHRw21x3yi1LUDyNY0G7Lsj22acgqPgtLMp2hfyaq4D1pvUL+WBJS2f1aJwsHF5
muUeHvGAtiUFM6a40u3mT4XWBzriZ8HrqAybS93d5c0+Q5vHp2vK1WzkzXhWQQq9Q423Fvulk/Dr
RqxrvzqTln9Og2oj4wM2E5r4i1mU2ywAKhBoj1hRFAbrtdmpYHwuwo7C1JzWqWiq2lXadS1CphGr
waoOkx0d8GX1FRZclyWa6k7dNjvaarsqo/rR9T+94hX5AFgkPrZV43NYwBI0AdwJA/KLQmidb//D
VF4smarky+X/fXOxYzn6Tl0hn0+sezmSK62k/GxVEH+zDIYjAfsVd8O8iR7yFyHCdREMxU7XLopm
1p/5Q08+BukEQEEUjGutM8ASQPXhJDx3Oorm/hZL+JQ+IA3OjCLeOjj2Bqejex70qkcvg9uQ/a7H
DVOTfeWTbS9tTTkI+GuonkG/5TlMSxN5c1IUhvb0Lu96pNOuHm/q3xFW2KWLOORDYL+EJXt7j4AU
M0+ALVpjhDsrSRzdTf7tyy/OQCJM272Zxjvv0oNBeBx0HqqiryY4mDEPrlZqAmMkQeXLiqErWb1e
C2TRmquWjuAK09bPAQ1d8fyAojWSN5mmlWZHmOfq3zkoARjXXtCp8cC6yA9wOKp3X0PHLPuUbMO8
qCf5gGRMY3oJ6ePCsuFxrlDX2iB9CrYOdoTr2tZTtpFNA4TBkjrEz2L9B2clz5VP2eArbUoYXEty
EJ4O5qDBgeIaUEbYjdCs+xSNSOgH0E6KCU9MGsfIk0/Je5SduUQ/W7XLg1w/qJXHLk91koGZlQMr
QMGcY/yuzCx4xryBLu2MOH+blZOm7OdkZeH3cFqUf0OKo7NMw1wIqKl9FloZ/DIoh3+YKp1TSwv2
SMOrG95hgXHxOKs4W+Z17+OF9HgHvlfTHUHiE3iKbys5tvZCRc7tvQWyXx5JtQg0ZDySYTk4Jq7P
wJSyQrId/LwXdlDmyIavG4v3mt6gOT5kkPjAR/Fon4alC8FaG8+3p86WyjRueMhIq2niIgjS9TUc
lHCHHaQzdG7thrINl5wN4xSrS0zG5yImsnHz3LVQWeA+PS6qZy6Dz5KcXTP17VxPJkAECjr3fCQ+
iFR29+Bz9siv2RTor3u3yf53e47qeW+JP7xGE3Ny6RkGUtEd9D9N1yur7VFOof7P5mgqAyD2u8mg
ubFzrjsy15/fz7wxgcd8zbAG0YM+JsXiv2HifM9xTMNTfEa0DSJqOes+pU1uKvGdVz0KE/qPcOES
Q5CTE180iRuUMViunwMIefGx10UDUIQ/5/U0zwjpv3dE/MKDhJNmsVPt+qBsuEE+FnUoiDxNEGym
xRhc1y2R+wOzOUrPbGl939D3I2QVbjsre94Frw0KwRrq4t3VbvJnoEJ03jFqgiIwTA7GpWnTSBW/
ZkANvGazzjxrvfNkrYKPh69lBCjXJMQe+X7wUsQ8NFhmhMx/+tMaikS4Z3u02EFkzQCyPkQiXV2d
Pr29IqQG69XvGvxjZGIccJ54W5UL1EskiNBfLMIGtlabIk7hWShe/1o8XXJ+f6tXl5oTvOgWOwQn
3QOcybJyQYhktApS9tYzhBdn9SOJwgaaNQAtfyrFAlqsJCpmkZ5uCgSY8/gKCqwPaDHboE4aE2Vg
d9luSCTyuxUrWjoFBaPqz6TH6PnkVAoNryMJdVwQHvbwR+WyYasak7RIAWidg3gUkSWsiuqIfJfz
hDXe4mjD6Dun4t9MYgIes0D/N1j6VnGxxYO9TypmO/4TkHZJfvqTHCR8x3KjlJBE+gUClFJ6pOgX
LEE5BqbeRUB/PiykCYB4rTKerCkA+Y+qeN3BRee0eJDlgQiwrPaXdV66/nmBDIFx1eprCBDhd4yQ
QKhQcvEOK/YzfFMQLMcgNiGuVwNmMAIVGeLF7ZSZfZgfpn0Vee5UpZbLthNzRFKrvyFmwuLJzsjF
4WJs02p9FPy0xXUiXYJxZh7pJAv5268/Gwb37IY/FOlogg8mNAOmrP7b4FO4AHwaQoMDJHqmI2hQ
LQW43WJJ7XZ297QUnSYT8xX/hz5C7IJGQqnzmiX13yP7MjOfWUn3Qh/nlSg7AIA/2BaAULnR1KVg
iH5o8Ix9mes6mlIfZq4OQtf3K+e6sp1y7ivyk0ZEVQIUp0dYIfJWgw7FpJA11uk+0fKUP68CpIbB
jBk63FPG2oEvEuFUrr1uw5ishhmIhvk2Wo2PZ8lrNxDDxdSexE2nGUe2Z7fBQtWAiUbdmaPnC0Vg
In0ab5C5rksI723O2dzty+gTXvll4OPBQP/RyF1Mcj9CzUPejs1yX8qVBjRT4Xh0FbTFNWeb9Kx8
S726Bel8ro7a4lFqd4NuGpOqocVWP3mbi0iQa3YGL7g2A+Rk94pBboFvXnkBLrJOJcKJ/Y2+RjdB
QTsory4n0viFaETC+34I4Wk+jXhoskniOdUz5WFppZ6A4mc9WE7CJk6TDpAWJ46IX2M7gTALUAY1
ZJ5O0pyFWSD/If1yiGbnULZoRfyA3txc8iMnASeNES63XjZi20n3xbiIDNTnAnpQRtPhjUqbw/HS
gb2DqZKkx7vdSQf2vDGHCGSmJjjDXa4rGtHCbVpg+mx9ehAnYPTFYxnTDc0FEv2up5k5Ucmd7mpk
kTibqsrnu635xuo9bBs+Nf9livDQxwoUbZtdith+l+eWvIw/L0v9T989qM4jNYfWA9h66kzlttmf
M2n4L3D2guDqie+cwJ4cRGKQAPgKShJ/KvCM2wNOAmziALH3+aKTOk3+cWcT9zYPGjdHG+9cOvZ/
CUr0HKh83kwJxSjlJFLZP9u166syoqQ0B5ns0JTS+/MnIoK7KiplzOOTrTNiDGgtYwC3WE+YOIgq
LETNK3iunTVW00eebm3TB3CuiE9B7CiAkuECAjX1TAYJlOvDV2xhv3skrSmAgRi0JYk9FGVaOaLq
Xx1lIbChpSDlZde7lpQSZDe/G8IZ5LDwft0T9NrU2Y+0/jM5kPmJk8F7NzAqpJXp7j4i7qwFiyrP
7f0TnZr6+CeYu2woCG6amDlDgn9ceUhAbkJ/0FpAD9uSI38vH4qJBNcI929ErZwln/bOc8zUgezC
KbGZ9wXcqRuX9EMF4GbZeoAHOSEDK5uBpnJiMaTAzxOxMQ5SgJKJ9/a8QQttjI2L6pYcC8gpeDf6
1r4YLFU4i3UdjMALxMjPQqIVQn4Qbj+KanfAIrxT9Qxc50OflvmLd8OV1bMbWrZfxtnbnyxEkUU8
jahiMKvDOP8G2MONJokmjlPubKMnZx+eAFc0O2in7p09GyKcPYpIPThfo8BgwevhUPNN/xjRqiO6
+yJxTsg14rK3CSAzu2AXPDRc0bP+Yp18Yb4PL02D6AmSkdeQr5kTXEBArJT7hpAQFbEIWbaP+HAg
M/oqwtYOevll/2ETrPL9kiDu7ZZ5yhUFCdpNpJvfNAJM12qdPexSIlXlIVNGXVb9VZ/ZijdaL71H
ONeqli0OK5DYlYQPljLyG7MsAL5PNsug0pALDn+P9HXQFQGow9m778wbqHnfgKdgmUm31AQO1h+C
a/vsT98VTrvjWleDIICrxPGpoaCnI/IRhBPks8pMX6KAL1/UnVewE04g01nlbC+1yHXYZ+qlyEmx
TslrRee0HZh27UaTuuhbcp1CvrMpCI3431+GoECCmVV1ZVDQuTJTk3jRHmqTYrLLswvPE6RmEZB4
u16lSt2yJ0iHdmJCrNP8pgICY5nLbGCu6M/rsYFA7ycfBM+vvwK1A0JSCDHFCgt6O+GEJjN7ze8N
eF6O6UdqznjSmUcSXyJchmBomYjOybcVF+XLReRhwCnZtZo+at4gn4HPr5Sbcxlp9A0PY9lkA6+2
swzcVBaaa0EkaC9zHXREDO+mtv+YHnAZQyme8nWzUUtvGmbVO4LB9JN00VIvbLKdW6NqeqnxrNl3
oHq7hYf+sp0uP6ryLTyTHSkWbVKTjWltNsAOqM6ZNNklGKLDD8Jjyx2xj3Mm5UG1jbSCHEW6i5X4
wcvYAPsXg5gwWil6lgbayIeEW1Mt+0D7tOBtwmP0VHuQUm+iS1zpzPgqrJ7zmB73xAy8+xglDODJ
lrUKgGBETmN7CJ3QBoeYPpBisWy57nz6PdDJWl08I6q0wh1QOLB9J/iKIzGiaFE5DSQnYo6ZCdz1
Bk9LqTFb8xJN41d/rLuD2OyUsi6ytvuuXNkhjNLd8tX6eT/knLuzkLdRgnZtWLE4j5dxpaLFR3vg
YUhiwt40Ob8N91oKOz6srw75ZqlDUL1NGM2KEO6mnsTJyMc20ozGZ1ZO65DRqhi8IQRPU2pGd21Y
05B3ZERE9Y08t9zb3pu1KtK0H+DJxn6pdt1KOvCz4TYVrhNS9YXCHAgxNBwJbDEZhwnsQvyXQAGf
aUtmYNc0b5Y2I952f7r7cq84SabpNi2nspnRBvGPgCe4LmfxDfyYk+TxolRAzw0TgvS8CoD0ilpd
n0VxmeY1R3cj67l3XUenS7sEybvVE9GBocjLHMi1tnIvXRVr4cesjsYie9eILnHQ0hY7Akom3bY4
oNIpC3THh2X5SBIh5OI89eLUAhOQQBCCTRVKuaOeWz5vqo6defERBmSDqYcHyjMKDicndRmriVqP
zEKEn/KhBhqZrMlMoM17C3P5ETWkUO+jbAK9nwM/j8YvjVk8QAw7pTNLfJS4z7bT2McYJRlI+sa9
xnocWtNA1J/poZ0wSgf3W6CznY4ZhgC4uC2C0P1iIz6Ag6yxyoItOTD7/O20xVbUi3ao79w/l9he
vsiP1bkN1PvF6P4cf3WVNoTwkjLUuaU9IJwiTQ8wPE65q4iCx2Kh9aDSRisXmJQoZ7zfOh12ZG7h
FwPXhLUA2j5Gq/mhnG065zqZp0QKhy4EfewkWegrH2luep9FEocH2pMu8L45y+CLRVxH1ETUmRQV
6Jjv+UcIFrXSeq9VO8IujPi5AUhnL9hhy6ZFdNn9TZ+9ShMTb+raFC+1uDvFlyBjY6JCMApS1sMr
2U8ihCxrFDzIpD4Sd3BE5MZTSypcGZxrTYA0jSq2elqUZTkNKvzKBABt9+9heYAjmhoIeF8vZDKn
KMaiqnXMYGImgbrEjjBa7GJHcx51fb2a5uSn3bQlLPRyUSp5IjjU/oW/viInFaGaLYPcSnYu97xP
TFIuvgYEZhRkv4FDX3dBG7/VRFN7LoHqpwrGQU2S/TN1dCrS2j/8zwbuWTyMq4Y7JYly0hZ9X1Ze
iwUDYCbBM5jPjA4KlrUrUkVKpw4wd7ZDEKovSglI7+J5nA8oXYt/uVYN3Rr32mOapLxsID8d9AaK
mIsRwcSXHDLCpR1mIUrPVRT5dv8lobbUlHCpQYJSCA4kk90RWCp/CYlUx9n8fLYfPMgM+KoFN1ns
W6GBLKFEpNQOjeUjqHpm+WQGFsMjq8suwOpl6BqFqEZ4VvRT9tKkrh8Xi9rz/+/7jq8JXbOmMrAk
50OnpMpDXfcfdVAhiatoly+WidDbvSDjfYLbbwb2WhHnlWMuMdXwX8+BTvR5CdkGYWnStypwq8u5
HxPqKH+rz1f+7w7T3lnxfvsWtmEhUZ0vq5c2QQNDftFNxUrTYBUwB3ZbJNBBQiLLTrGSeOb642mI
WFhqlBsnpsOvD789iUUyz+/vV2RAoA/G2kH4Q+dxkmxiidAo8Zq+RdyXAL7Com04MTJO0JCN4B9e
ZNo5JNkPVzZiWd1HIV14loSLr9k9TEjcqPII9f/5AFdAbTc/kUAnbvQkpS+XZmfNZWbOH8XJaWEm
F9tO7gkKsfXEg5WgCOhqudjgi9n1YDNRfCnr/vYY50TcvStIfJ1tdSqFZUlYZd84F7ahBWIHmb/c
AGpuGySauRYL/vBZK6/QZOqRxKsW7Q8CFn9vMvkFJkf3MK2NlZirp1yPqik24GgQQI08xpXamQ/g
V+T5lAIZ89LWJiDlEIRgmhx5L9Dkoy2WcfyuHQ5zHnMkYsZRzR1kd4kAnnfJL5ZB0h4gv+jb4HY0
1bTeH0ufFLVmiAPxEn9KfpgIxZw5rQJOjrd+tue7L6gelLb1RnjglDAPiFYsbnDpGG2r499rEp1X
ftsNvn4SlyQIG4P4hXEAOxx9OXzuukH5nMfJbFOG+yRPl+hyxFZvwSJqWEpiFdbMvb1UXvbMUpmw
yn5YLCZ1457haloYaMtNUlrgUlNYjJf52ITa6ZpibNZxReZc15ucM29Ig3dLRqg+ENtViIWv4CBh
BXJgBAmpupc97c5L9qIRpvcT2KTG4P7gJFZrewy+NSruneFg9KOkYtvao4bCem6HzA4DQUcNbZPB
ST1iZonv9Thw6oFl2GdnzJktzmlS6PIn+KYnvnQt/9KiCHXRUnOpBWbe3SP3titbD2t+tjj/D+zH
DbyECtJioZDueOzTqv9smufefe8tO9xHLZY8Z0FawZ3zt9Um3lqOojaeQgZlj5MkDz1WMWbM1ask
3lCuGPaZ3DZqcnVj5dblR3U85QVv3pV9DG2MrDW5nK2oFMZ3SjRdlvZ+kNKKqiUKnpcAP8DRoFIL
RpscMNsm4vy+DyVcUAT9YbwuyqeVFp1vId+Yhc0aIWnTrml6UANvU17E2uuZRsNbCZHtgr5EqYwo
Gsx42860m1SR4xNKhs9SJn6Jacni/30ABi4SR6myJeV5sLypecJd74oisOAwImUh9fhhseo2Ucv+
C1Sn/QeJ4fcWmYaR2gZ9z8pcY3fLCT8imRM2ayZD8pVWzAdJU9/xUQx6uHyvfhvTzpIGFMVfPyX0
9dkDARgveJhlevNkF671OVwTE6COiwuQgc2hKQZCP8DObdmjfY9EWbKMbuBSW2PdoVZ5wBJGjw1c
j3PVt+3yRJN4j93vCEji6jDpZZ7p9AvYwsnTFYrOZct10NhjfZZ+pa5MmeJuvtZiGDn56A4np5BE
jA4mv0IdCuU3/PRk5jYnDqbGE8Ze6G1IPKcY6uJI1lNbUimN8uqDFJagbb/lXYZQBLQuIkYAy9vb
kIZXGlfOgsr5hJhNcHZOkWBDiQUvKtyiS5ts9VbcLYw/WCnbfdYx5ByG9snhipHhYoFR+XbES9+j
CF9PqcL5hLRjNw0LU9Y8GcrR1Jocob8t2n09kgairEQSo2Z1tmpFJVnVXqX/i8bMNGvSLgUqEe5N
NZ4PgNUq2z76+F4ySdtzFgepTT4y0ujFL+l2Vk1OjPJnGoNsRRtrGCabQ0kAmiKMYdQh7Wnhl0FF
3Jr7UxkKaN9+5Eja0DEheSkt8nectJG+V157v8W8NrfNTcFAfzDGtaSTVQuL1uytcoFLNkgdIHYr
ZfxIsWN+GAb5Zn5q+l5A2Bx65TJqAtTIZPxBlGpc/Wh6EwVaJPfMKAO993+4q5w6zwp+Sb0tsRep
firuyXgcd5HsOXyvvynt2omb8op3ObWBwcfkw1o47AMCxx/aLfNLPpF3hr+BLcmGeqHWlwjfBy91
E5nV4sp8ONcEHIJLBXTFOv13xRsLxyg88X/XfrAvg/0IfvXwUSRz6RHnYH3O1Y9fQGVk9Kj6mriL
M4H9Wpa1qtahBk9pi9SKD5eqv231SDaDDtmzLv9je0MAFY8iLCI7D+vLAmj6RlhMlMpCAUdB/rWg
lzCKPy4f7aPEL29K/Yn+XhPM65o77gxoJeVmExrxr+LmO4MB2sVaKJ7VP/3f8nVuJs6qGoCthQwj
6skheGGG0Y/QOL3SFYVUboIhPqOFeb9/a4ghzy76sGrDZlPz5E+iK4Qn04S0AbWA0VRCWnmXUM6s
amA0HIfNkzb8D78z2MTUqlJMFzJbv+D9xqN0qcnTcXssayHAYgc9eUa9e1RzlC6aof2A1ub7SyTv
A+AWlel9oXpFTAzZxqu8xE4eTAHMHESGgozHMNwp5S8+s9r+TDbj5Y+MhhevbiGTnwGwJcCKZKlf
KzXZD2AYcAb312EsXipytba2Y1H+QLQ6U5/TtD06oMSIfU08HvedzJbkRYSg7cjYc2c4weGSwYwC
fKAaQ5jIgCknuKTkSpoN6HAv2pwYNPmXhnGnwRqbMk/QjMCiHbCkESNal+PaMd6JM0QDMQnltNyj
O85RrcxOTsr0n2BW1WLINDkO+Gk9+1PgYIhdYwoEE9p8BhyrXryq8JRkSnE1Pb0xsJQMP30Q4Shz
D8vnF39oUKwIzDt/CjHX01vx8NeSrzsmbzCWcNtuAnV1jOOIwr3Rbyj8m6qYQysHf5fUFlN/PPQE
kzK8bnKudoh/IgdBuKWavDqo6rxofTJsCvCYOO/GXovIKxylt/9Tew3QCvO8zolL2FIy5zlmMVYs
GlE2zr5s19B+iUx6Cm6lS4tfErdFG7pEuHM9f2ihBiI2WXoIsaYQqHm/sTIAghOm7CDwiodTu9m3
Yd5jwLbgKi80WvNMqd3u4Qv4SdWGGbXwVtybf/gKXKV2/7SWQT/YG4lyXc0XtTyBu3iWw7jZ1IM8
7OhPCThX+r4bfmAdDZFqb/oXOz/wVDvMj2/HN+lMjR4WSQF8UZB0WmO+O7B8PRSSfzRfI0aetfcG
fPUrgegk6dqzN3yPoLjjiLjB7iohtTPkF45Lbjr4lLcUxDdLg6Yk+PJm6DEXifZp7Wl+zHo+jUGh
PQZvJvcdoWlhOD5x/QzP4pSeJp13bRD2PIEdmvywwc/vIZud7f3BUIphCF1FV/tj98WqCoLVPAu7
BHAnyoRlVIDvH3fRdfWQAY1NnskGH9HMrHcAkvqDDvE/YeIgrOCrfKv6JQHDdc8XKJTyasDfM5Gz
If2O6VtQqb53UxCJHuzsXbprK32r3FrYq27KftKYF+OCwfzrP2TNceHyNjFM8sNYRyDsFZUWum4/
jFa5662zosEVHnEbzRdeDmRr4kb49yLuJQ8Q/5b6m3B140zlTYnLajwK28kEmFk0tsv09S/vMSge
op2IWkI3kzMmOuRJ+bq1c+vsRmGxBQXbRySfWLwM42Kpn9oPdNrYnd9oqjYaaQw3wCizcAuXfoWM
vP6psXrHeGdyZz44pOnekwTUzolHlx32GNJHdCBcVpNYYa13nKqQqzsJ74L9gITbupALRtfajGg4
BbrbVNoy668pvSdvK7KIjcAfQ0g7fNuHKfbgK0wVvLKfkaRQ7ED3A4p6jprrgUotXGdpDHVylQXP
/yB0L5jWodXKkA7j/Oq1IH7glLm70DSg50C2e9W/iWfzkUSh7QhWJ+5h+NvoyLUE86B+hE5iPSIl
SMOH5zTbN5pi/NE2nwmWXXMBd5tSijk3kQtzJ52y60nKdEzsio5aMza/LJDoTqqbf+qIbtjogbWL
NrnkzHxvrmkzTR31OIOflA6/H4rZYzLQVBYe6oRDUY08YSXYZTkXWU6NdF9LU05q/nO8qx5BEbxR
QEBMYha3IC22iAYlBUv6ikX9eLXIqs8obl97pgBiaZ0KGyfzFole6tVdGvk/i3vf1n5bOc60mYu3
cJuEPs+A2ERdjehEz776qcIt84+sU9x8twcVQ8dGp50oH1DJTWpewmVjbRYGOX3z3JNrVeYpGH6y
6MfwMe+5C0CRLD1nTYtTweB7xpUSpJ0xGeS0MBx1xJWop+dRxgKwY4k0JvxEuWOaEyjq6ECz2p5I
ZOs3IVQfqZBtDAPeTY3H/Gs1F1DFwIbuY/EZpjJZtZcaNvyQuPJwghzmDYiT/EmiTrTGd1oVQFT/
3Ishu2ES+kUpOqw+nqscA9CVjPztfgb/IC5yWdto269rX6xsicwHzUP9fsHLbhunKngcVTaXUbMn
vNhPeOX4xx0E41R5+ZhHBGzDZXsrJVukHvTDovzJ5GusxhRlcCDNrrq/boSpEyeHdF5zmIzp3FwQ
wTRby4nJRMeyULLFVOZatcM3Ai7Eg3J51pbGk44sJaDWtHwTGhm30OJ3YOFzPPlOadn6S01Gvae1
vUpl4wpp02jJbGvlRgw0FP+SIOMAPd95v0QVLnhpXltujqLVoWwX1MX/bKIAZUqkMVqab4c8C9xx
feYb9gmk8TiXFWzcyKz54jkIQibxOlV2sWAEqmYksiqYYuPkPbei4GKSxNeJqx9XbeSpbBfriTiH
BsXtNqAHhAEwIpjeXoms6LIN7ypyngIrHEqAt3ObbPeK7NGPVMqSwHeZmPsW+puMPQDo17y4PT6v
FL08UCMA774hcLuBiaHrDpDKjbDTUivQZiKaOdVx6t2mOu/gUE8eqHucAJ+3lfBGQToI08O4SSef
UbaZYLNXjeKLdoAnpTw8MmuKOCwrMQcLGzvt989qbh892J0oI6pwhjVASNcXt9f4FrP/rQf3/1+Q
SeM6CiQ/SBLmRo4+5cBJ5qTP71vXy4MLDSCL162szkV1rRAmUBh0pl7ZDUn1xOIfLLLXYe5gDVop
5rtlc4eJMm6xfDr84wroZ1rHfiQqUlyFKstDTsbkk1ICyJ5bvEkVS8OdbbC7oCQ1/7TA8noENSO/
DAi/eKpFtSIQUIHsbRs9XhJf8vOPqkFeiOiU8S2I4Nl8O21IyJd0T108KbSY++U9fGRj9vwELBdc
T5EpX22XzLr/BFajYBkB9hs4593Dl16tUCom+smiPi/+omWHdzHjtP1gZ1K4LN6I2tCkq4dGTJ2/
Oi2S2H4A33b5daWBbO1rjJX4U9tjVQ5viBmpfekr6ZG2xlFVEydGYuh35GJDnIcFQ4/WVEBDgceh
RaiykfFZ0rrDrBOWO48E+QmWGtdtl6YtItU+yaz3LcRZYQeQ6qofqdNGTBHVcHnRKKdWIX8XCt9p
+uIlnFoNuaMJ13N3gCI+MTE+AM6r8jxw0N9HzEzp8sBCUNkdm8dmTLe3pNZURjjtDL2qaT5D/Ri2
GrylNSb3m4yLc96ezzgZetqvDqw3itXOjY453vzq4ZD1CpgRHutjvEc2k615jcIyraSpjSuBHY5/
dd7jc/W9x0H4mdEKd8M8DtjNsfQD5/SRiMf6TZ1oZkdfjjikOZFb1YpmXOXks24sJlv7FKDgz9kb
TmKYKmy0KnpK8FCE047r15cR9XAXOi8cslJib379lyu9lXQnVngj92M7dsbFAInLFzdoCKXOLNqJ
eEALHZd2GZRUpOQw4LCBkd1C94II27QbnFrMygTJUeBASrShCw3bsFQHeOZ4K5Szz7x/Hlf5ZteS
kDSPR7cf+IBszXW8Zc/GkDqr9eotGfY0bWVMeb2KeUBaZItF6rqzlWQu9Q/Ewzms3ZsMvm/VrE2m
nTQIvx/Et2ravFTfYhOPWl/UccdnRLbNL1b3r/aUoz5HSO/dLW8DdII+2YrFHQO3yjHEa64xvQ8f
YYvzNytLwKWaMysPW5BfliS4Mv4KXmvro26ZUyFi+arBGp/g12+Dujk8SGSESJkBYG3r+QM9iltf
WVfhun/eUx24MTxG7/aMCWoddwaaAhCK4TVOjsSbRdpORK8EVONzSCxgZar8EyaD7uP2+Gw9kjPk
Dy4Qw9JR1wB1bQ6lqM4Ao6BwRl3sSvVue55QHSL4v7+agyZwHdjs/qR6SQrmXHIvFb+IcGR8fTTg
BPs/Gpy7PIHD7WVJAOOjoQAMKCW+TKma+HyZfvzdwgmdSBPhcg2wv75udXVxIOmePs+0Hz19CeG5
/7y6g2OzPl7Wa+Tc4DeavybzG1i7rY4VxTpZ408OkwrJx8w7eeBwaiBQMHgrnlSX6QWf8y9i7fx/
zgqVTxhNs4SsBVy0E16ym6u06cOa4/nU6YowF1bY8a8ngd1xPA6LDkpT1FreIjEIzLjFqt5D3oiw
FLCXatdbyzLf0l2tg7b8oh4u7U8T7PKSU6vov9pXxr866QeFCWoG9vMFwcL35IVsFsK/CwzRBVVj
VXhWBlcWVeVVtIwjvpykfCK8iXtYO8tggbW7Fs8Fi52qnGy9qFQQZqN1llC2BNHr6B7jvK4GHM7z
X6CB9zNazydTmYwYOBs5P8cXvZbenMDiNXMSm4OxCBlN90W6lfLxupNBMhbbNfQCaazFu6U7gAJ2
xZf1VxXFwYLnDeMbi+8D3uFkb6VVdRVicoP/OymM569gboEz0e2hJKPx6vQdj9KFKbcabQ1MIAPy
9tMDTgRdWSOILniuTkJsYEsaXHbo26DJOZJGnFDJ+JrOztFUIWxScCgroAMWRz++ctFGM7VtG5gV
xcb9eD7rpYNbknzL9q/CAnzd84H+ArX0szpiBzWgUmWSC2oBlp3xQfFCQyFzJn2igri5SffRQyU6
YLpRX06IgWLW/iSE7tdQA69owopPuwbNUf42iXoxS7c94N0MEGowRED50NhE1sYQ+lMaqxe5hHUQ
i0zzcEL2X3W6p0HLAFJOOpD89uJ52RYkSjlhhgdbsYeQLDv/9iDglJLCEyH+Ob6zXhhikOemfabX
Gx75VEjN3gY2hp6bZkP0tcdMMoCNkWtXoa9nx8kPNFfGafhybjF1Xh36ZRwiUPhQk8hBBWbd+FH0
871P2VvKtmAnzyhOPVjI1D+IHQf5ubQMwLmJu2xLfErYPHAVMXR1FXy+5iZjNbnSn7Gydophs75K
zVH4RYjAm71IFAK8fuVKte1ST2/BL5bueX/OU5xKZ9KRaBhwlPpRfgBfhH9aD9p1P/x1VyiNTttR
Lf6ambJ+r+WUUJ+ujut+koEE84nentOuPzDH8iGBdAbI7l6er/ClSNRgpccTj5yas3cNwNhIx/gd
5Zbc1MJIGzLT/ozZm/HZ86Ewb5xPHDXzmdse08EsbAAYPd3WVufD9+s5CclPS+G5/zOFSnbEBVHi
SkBr5sSLrpjF9Q/Ym2uL2irjtHh2GC5NPElyTM7EbwS+iIDQmxrmoqrqldsLvZ7cqWdoSNMeBXJl
8+QsYmwtvpFEt7pSYdT7DRyzPHteiqC6+RG2o1xfIMWQXH3EULF25cV1GZwfR2MaPKYPx9th1Jkz
BpBp3ctX2JIHqcpIGekih8Oj7xAC0MkDDTGuUnnnrNY+Uj9gOjKLx+g/IHhRSbmkgV3HM2xck78V
R6U4UXFqmTsp44Yx1PRd5rHXe1jcGt7TIZ8li7nLJS3rg94d2siEqg54sOEJJ26zwXzm1/2I35wk
uFsHSvJAIXqs65FY1n4c2paKYZC7OIu7IZDYZhrvV+LBWkqpQJRiJXSvqDfYvtyN8dq3c+WrFP+A
r9IiKAbUCUe8B9e/WDjY1SXaBOr3TLRfcHG+jYARlSHwAYkGic8zDmv78EFmjrsh2QEbEnABtqBP
/CUePRXkAQvWoCxz1/46ro3Aau6L1GLn35+T2vAWSH9HjDo2uZ2czccVYkwZNaaR5+4B2A8113mL
8qBCiUeEcgcn50g7rgaorZ71naIUdlYSzSdpcu3sv4snVXMYeDnfaJaHEILqvOAFwfI0rO/9K6l2
mmxqEy12x8QF2avudzjPE7wRsUGF6PnS8wrZb8M4PbG+IvEnYbJEqrNbyJhzg4QWz4BajvSmV3D/
n0rlHzR9xjH2HrmWU1AE+lMlENBN+W+sAzpqfikNyMI57fSsLIsx17gsTvG3lPdmL/dLUFhTbk3s
yLLjzVQ7uzHoTID/a/gHM2mWao/Liyn8S9auVhRHYL6RXpr4+82veSpoPX913HDJyMCofTCMsCVV
LtAT+RUMAJTjWZi5RU/mMIs8H0Dsf4i4gU/23C6cf5ClyCJb9moM27FtH+b9gDCrzojNmsvMLVRd
MFeiIfXXAK5ebn93zbCcbrTe3l0qpBrc9N24YTyJ2GWAODI0I6mesTXTJkIA6BJxSwm8cyF6qAXM
vhSAOa+zHCVafNGGbZipnjTD+vVa9O9FMTt3/N1yvV77F9fwar+WeZ9sKTqYM7CWjLxtrjdViVUJ
J7ivh8dMqfvU9V97n5zbFQgPlbHYzqytVGgvmEGVz+d0hxFMfhlYo4TFVRO8HmlhPOp5c5r8Jzc9
iDwfR+lmoYYOs6Axos+UTSpLqK/j2gl6HlEE0imdK3LJWZu+EjLISRWwUrsPXnnOya7dBPIlH3CW
J9UfVRmz3oS90ilz+dXKRtGZImBObVjoAetPzpl1ZfGJ3t6L6peNff/bN8lc+0ojbDI8ccIAEI+H
mYBOlLIzcJ9gH9DuEXDBAnehMVIsL+qaPL4BQnGR0wXdjs9tGv5ifWwxIRCWzkaI7zRDN6OuvCHn
txXTcyC6Sytonmq4DW6sdvvmzNDV9XO08hWeyzVL1kP5TN2QNmnyVn4RUP0n5IKy50QDqKd+hVBO
fmwM9LhMs4HEac9ZLuxxGELwQPjNZCMMjPWtTm6I/YuIpQlNFMG3VrElw5RL0cEL/N99PGdlwYkN
anHjqYSbFUFOzs6BeBsUEFS+9hM8mHn6hLonfcd79/uLkaXNH1S33ADmQmG6WMn/+ihl3x7Hsdwx
gZ96568d3iRdBrg0Bxctr/mQdGQH4MjyEJfW8u7JaxETKLqoq9tSDRSvvjWdwYlZT+lAPQU1pgKU
Yaij+MLnR3bVNm/BNBF1t2+/V+grHGD6zs4T3oKHkE18s5uMXcZGavqXt+u8AtiTQ4VtGPsHrJao
pZ0AG7wAKAQWVjn70YnhFPl4t9ABbdD0iBZGOjb5U1V9WIUmyNqlfyuYxcMIR2uaetnNqrPVy9yf
+LDwvunefeGesjPQhVeZu4s4qDGSsYjh0dT16xn2mUKjyUKnE2ZN3dYxArTmiGWAn7CnzcP5XyCB
1Z5bzaMRb9Cu2+jg9XPMRZVdv1Vttp9M+qZ3859EyW/2GBc1yVnJUqtL+TuwEf/+Qt+N7OkyRtB4
6mCDprhRMCUlGPWbxOpR1VMbqhKx/hn6oz9fa2fNuEj7BY5iykOXSa2WjOrPznt6RVGNaSCvvOXS
RUfWWHWQTRKwgbMQUYdtWUx9qyiJhr51euPnP7GFCAV8Tet6AZCbsnBLeIL46JfQ7JSDPYfHVo71
EEDNLboKssi9pR+JIiFU7EEOfxz0h6SzoY43koR3wCy7/f6kNDW9j5szgXWTj7RgWQB9wy0yNaSk
DYOLnvLt8SLh2ktGLXHaUfmEWgVZKVbt1lVs0Xd7NwUhM6ICF1U2QnJ9aJsR/Ei9U2CUdEdellyP
Xjj32gDJZSN2RBrA2hp6qtEmsXn9Oe2lJAnamCWJ3pJRbeYl6xT7MECgzRE99BA+6G2XAQZHeMzY
32QYnEfRfRRIW/IRBW08OZ5DaGRLjyYOG+9jGy16VXkUdFixt+5NUNwCos19NbKfPCUZLOH0i1+v
HbFHkPUkZ1O1WWY5SwejRxBauOxRLw/+hQLELp29zBbp7IYdsXyutCgMvhA3jbD+KNHAQvbQ0MhO
a6uE0pUygW6yLuZU8KIBE0LTXrhdP6g3iQ8A7zL5io1XXgdIvpeEyK0KOx+Wm+ROYmKhn5tWbFwq
wTz2lpNChk8vtlqWgAddIipZXIwceLcIZSc817FWVJmXWVPlDgG/p5nmOv900JkId5d2EmwPfOQC
/+ajfvdzq03tU9m0Hf+pr3N7nrOEN361Bv8gRWLyMaMu4JKyDsrTvRQCQ8cMGctqhv4bls2Xx++7
ylIbLgXxlWtFRzx616/bYMdu50jvJeRdXtFVsEwR6et4rXooz91zeRfY5uNJgW2oR5u0D4SX/LKY
fflpLFNgFGyAr0Z/Dea06KTAiWweVkHp68XO0tzPJUitLZR0wLBvlQFgTayh5eMgrlLDTVJ8GqNN
12XPd09TIYzJLxjtA8l96JxH6avvhyQ1EUv8JSAGsxt3lELH/IJnfWqrZhc4Kq5dM/eNRStDyH7J
3V5asYbHY0O9VVgQ7dR9TxUceEeVZx4b+JPmh83dpkPoRv5vb+kbDPUSlcWwkyPTa6LthiBBx0la
foIVF5r295fpr5rH7lOcKnJBymcksD+jVVzMRKxq4hQl7nnnztIaQks7C+aH+9RvEvdQlmFIup19
fGQPgONJ/R2SSxDtTYbtREwSdajxtRK6AwY9HeQ1ykZX2APA0B0611sCLHzIsgD/oeRCUprJ18Sv
nfqyznbUft7LzdUiO5obkT70iYZZ5RpeE0Jpg4oWKRJupGNr1iGBH+A/RSv+3mJJRZktcfxyvRCt
vOY/OggO13/PnWij6W8xS40U3bWleJcrCCB3PbC8m2y2VbaXjW3xyfD0pdPqtu6Q6iEl9qyo7btC
BbFm6yJUu+SSALqSwWfSBwtP0q2DowMdVv9hlY02xYizcqZb3NL3m86gI70IzKT9/kfTpyoYFGQO
C4Ja3rkSHudMEWwMmQbAUst4pSYNfbgt3Tjvm6ziy8DBlOj00cDF5VuyYjyn2KuCjn+tyz7ZS6tX
drJKc1l82WtVOptt7uAYSHfxruqmk86iwHv/YWIHC27KTnUp0AHv0IZswDGSksE99mkioZ2y4YMh
3e07dYGwhtD/PB+XBBJ801TJnmFj0iwr1Y9ZCTQTJBuKCUxfNWdegSlZiiI5i2zpbdPcOvHKD1J8
5EQiG8D+yoP1mOc8ibvGd/Zsi5dfsU1FVohKYTjuplEVUaiiv13XZVYiM+c4WTId33dimIuYMKCG
pxmtqf+RD4EPc5dHttZGcg/B+iizVSiHKVPYwVAAVfHvXqAXqvkzLuFIQ1Zo549YMU1DBLoBdfeJ
2MMyYoQF68Zpgslrt9dQxEUNXOKguAVj2jLMITf3yryQAHDibAZXk+ZHcsbYtxW8dIR1sgP8mi7U
l05oIRXI0kVJS0GMw6yqtNq8jtaDNWIB6s1emBTQWK8nZRHIKfTLj0L5Vt077cmQu4eERUM5f60z
f5hX54jjCXKt3gmaBMVfrU9+miahblKz3CFDAhz7FDD3AZZRTrTLKj2Bn2gd++MDBO9qttGm2rzl
o+5lMN2wbKQzjM1GmJyLdGrBmnMHdCFMyaK0LWXkng7z1VMf/Vl5ZLe3FhC/jCr1WmL0zKPtb72L
ui0BsLiYAW6V1eTXuvxvBlzsVt47rj20gmmqJ2cVqLqGAYRM0NePm4vZ1QpiaNvM9jSt0VFyOdoL
rCDwk20FiYaU25oWz68cGv4YOBgG0D2tusJyFpHjduPZ2b0LRoAswJCLS6aSR+yiQ7TM8HHXXSpB
LIVQF2+jqSIG59nNflHtw3LEM6ng8qoYKbRyl+b/++vhQpSpHYtivVwwEhHrKn9kyR/FhJAn6kAq
qsW/A886K/yblam1CcFzdJ496IR2qNaSbRIH47fbUrseTRfnNSq/dlSNgbRuH1A8g4nqsinayf5T
LB+8h4iYVvcIq62HLHa1ib5wLiXgfiGlCgN6Od6msfIZUVNfSZjD+ucUFBBEfDbLLbKBbUNZqpN+
+xRkqSDds6QRHtIvWsx+BlHv+c1qgWaakBFZIwEfPYBiZgp2Pk7wdgOIAPtgd9Kg5uOInC8mhW4/
XAtXSGR7UgznLn6mU84kNiOsCVSsYsoxrdnqWpGSiiFaszDEBDXDgKxV2WkORK0Xd5/oe2bgos6c
8ZXFdYR/M7nWRsinyCU5/Nw6GNpCXG4hMN92RZi3ZuvHaglzw6ps8zyPV//U1b89PifQQzBgXIYH
7uc65o18vGhYC3UYgmaGmUV56vTv1U0nG39U1RVQUtcvoMaEo2Wsr/qZKKG8UVmPEiYEcsyrbqqe
Z+iwoCdC4c2nLZKIqVCstjZEcsXJLKVdr064XDOGnE/VpFeSCXgJun4QqIbajQZf1IsfvIAk+2PU
dQp3MwEgrFBTM0N1OOEU26tEXEzl+OMfGkVLq9dpbkoCB9TPqX0ENnfXkO+UdV9LuUf7YMuiATFA
iAsqn0P996mkbUuh96eFmE3FvBrFKs2yox3uNaOkrE9SBhDjiMdu9kHFWXpq5FGt3ZW6x5KxH1gs
4b52oV5O2v1pmaK9cc7sjk0Ls/cQwSC7R9qwRewypwfVw27BZx24paqAgptQu8/H2baMW+Ngb4Ms
BUE4rLpFGur034DaLOYhHJdN0sO7bPa2w5koHdVsuoWDOmiL9nJ0+/pwR/bxsvZKyDSlCcMaWfSX
9o3BbAw11DISvylC4/H0l0fTYF6TR/334wGSNIWkTtW0qwEdGCbIDSWahBqRKs6dShgb98+PvjnM
OEz+CzVyacQTGwb1XZayVJZKZgxZ5K2LFP7SFoOwuCOiobiME+wDjyMRtXFFjWolZOnuHIW2BQ8W
sm1uNiLDad5YjPAJ1IosWvgc+lrLU8LxW2SJnX67DuwjrpPq81XS4PJg0NoiLEtXxSU6SsMJKc2L
TA0W4kWf9lQ5ZES9fCA8AhWwDcIPSuPSwRjnnrfH5WganfZ1193+WG8V4DgOehsI/tTNBREqkLp/
iZjcbRwRV13wraD4yMGOtJDQB23I/FYGiJmmRG6KAnglywPHZNGowC9fLvjyXEOzCnPzwe7LxrvB
mgQx1z4kh6NkcugPvyRnmvzbX0WCA8+xqJ4MRZunTQno4kDl4Vj/kTxCGpClx4b1qyf35vNHFz+u
uYqdNbJBnbZY7jUJntA3iHCf755u1WKHIUGkkWWtCJp4z8q3UqeVWCt0ddR8VZbk79JP+lCLtOTW
gQVVz1pDEe6iozCipMztoj1gn6fCg8BjAT9KbJ9ALiYLLMrGNnmGbcpjHcBkdorzbjnEjKsE/NCH
B/tFMT8/4uCdKmTGWNcBWqgvRF4EHs0iE2wwxir9B/EXXwPtJ1erHkRauP5gSxFIw9aXXEkDvqo9
DJTz+rVp1BsuWRcIpfEQa/owDxguo8190rY0mD0vwoXfzLh53trhuO8FwLwYT9RvF9XfjhojGBcS
r3BXHkNhZtfM7vH0mRiZX7hp/cOt+OgH5Ijlq+0Q9ASL2GMyZRqHxQRVDkPyaj2AgnRaj8b48jCo
7hL+uY453rfLU2E/AHcK+dErKz9p7fCjM2cnfgp7oTK9yhsJ0SjnhpdMLdi4SsGn8tBxPjhHMYzg
+7WQRKvlw3RbDHRf9YiZXFWzGVyARvUuJvDhHtttSvec5f4tvVd2Kktcdw6FFRt6REzVr5ba+XT+
5K+WgTiNBTGw9anOdiWNCrrTIHmN8No939Fqm7HZjR3EFhBWZZLoGFu0tn8dPOasbOrhseftQHAf
P55X141PPcllwL5NlYeLzT79jXvTKlnvdM13P8rWGt6z+ZwPulALFGNE644rJvlMsTTK4+UaNQpS
dUKr5g3bLOMEpmnSxN9z5pEvE2+ql9deDKl/SJDuZnf5uYGJBcdrTHKDKRKE5OIxRL1DaGlBTbsC
fn0o1iCuNXTzlfzrSFOPEHZvf1MC7sAF5MXJ9zChR55ZYSKAm23zfQzmXiX4cmba+FSzqwE8LPLK
YO8gl9fsGXuA1RmSruuLYb7W4CL1N4sihOYngRMo+D37kLUhLnbJcSGxbRYjyBsvKQ4myGgHkY5t
DTMng4RmF/xSE5it2PvkGMUK+V7HihZqotEpaGgJFhwAY+B2zd4zqa/5nHbuRrRYwyV4lxwzIb4B
lAXGyKNwC0IXgp6205ToQX85nP5KrEeGYnb6bwPHrbdOtjQ3zPqoL7QiWS7yNV5KVb5eKN0AQerR
7U62YP97ObaJewbcK/Tsoj4ublIi3qiCdiqpwZCWFh96SRwnAHbXDalbuzp7hshjw7zsQke9qA9q
VwMOD44xxhSxLh627On0XvJ4Plav84XWHUr4Vu9A5lpaM5HkpdyLZBSmp//ktqhe2es4HCf6CtW4
lI9wZG7hpp6Ye46YmqQfuAc37sThnI5vDo8EJMa7Aih/P4b1Fb8QqfRLzdr5sr1DgxmFRrN42zdj
t8vqNtDGd8QAwSEfDZtrEwWQHmBYDTAOSlOcbDQod1ARaxnQjJN0ucBpswiCavB/4sr27EOAR6OW
EcU2mLoLuXHg9mYHvodGRDYvZS888by3hBrOIapAPOHKWWSmMQZUmloKK8PJ5Mq2yuk8aeOBJ92e
hc72lmecatSuvAqc0BpybjwarJvXv+2Ctc5LA+/xLbKVdftSwOQUxNJWdrcNw9+08igkkygoicL4
nRgg2rVl/ie9po1PO23Ny+8DLTw9X7I1XXvJE7gFCtWAQHAKMoOta1YsDcJyFbsI6tfgEHmpKuvz
LSy1hMUe8AOw+c0JuXSrnyaviE/ZFKx4XbWDIltQlU5yQ/TiOgeJLe1T+f/+7H4yqU0zTFppsL7r
iBBpmPooUGSlZLvVU87DlHtL304IfpLd0nFzln2XeCiVF9NkK0UjMQev4f/xVlJm5AYAIEifUcjM
hn1ObrtMeVAzpD7h5U+j+7bnkMjg98fkFdSkzR9vyxLt2rkHIyaTAkPnMucGzxYCnO2GeBuAc696
gSGwB9FD49Xi09VobMPNMt+xzVApy9VMWvs4h8+OALG3NtPB/sgA908BDk5L+zzFrpBQ9/TwoNsV
NNo7WZbJS7Nwnao8Rs/z1H/BCOyYtb/y+lkD9O1kbL9t4htUyG9NvdGbcSmhiwQllkvVbpJFPw1+
doG6lU+dxrGsnWdU4OmRrBV/DppMm60olD5fmVicGUfFXZlla/giuoH4tJhe9CQGc3n6Bm++II2m
XcTEZLaKARL6wXeCa67NFDauMWUA+Lux7j+CDW2vJE46JlojcMIlDYyOFNx5oPJFvRWGhoxQgwUX
sOKRIc0m5XP5oR8gq/sm6B+RqLSxFkSIHMa4OzO7OQRfsQCBxUU4sdDUpximbIY76T7zbpPqElfV
yVraiqdXOulMBJ5AlotyAHk5fTK2zDP82k4YN5wrF8LSGw4Gjqc0isFKsSP8HZ4PIg6NiHNUuDIu
JksEPmRVkaAAZt2823ZkiWVQdh0EaN4SsPPyuaThZYdWcM3Y2h/LhaIFuDVJ6GH0jBOjQP8YPj1T
cYLc221KaYkS1sP5sGioXTrYbQ18fSC2EdxGSdjXuHhYX4wpsamh49H/FNSvbfk+hMpH19ZO2hJU
QAfjMGB+8lP2UN9POXJ2kXNPRxS3aXAONgiiJe4KsBAiq9U/QZUKWcrx8j1vDo6WRxT1U5Z8V/qJ
h7yIFazdWMYBXwoTkLrqZf6D4AEg8hbNsZPPhYB9VHa6RXRmull407yB3/HQTbLgbXBctNezNWGw
a/UjYhVI2pWNcK8es8tqxOafUX8kr2erdNKUcQkFbclunMnQEgNbZguPc+nvDWLaNFSK1DhRWell
fsVoz2Bwp0ktSMhqi5Sk5JAOMJ7GXE5JlzDdiNhvvxz4BxBmjhqIC7e/p3iD5JlcTuImKfzzmKG8
o2Okte5ZJPQ2Nm0Z7ts6RK5v25s6oYaLtYPVZ/TP9DEy6rwQPsMTI4B6htZfiRyxkl96aen/aUua
ozZ8v2KRpBPqWfbcpCN2t5VuBvIcWZI2cxfcXlRQnHJYj/01U9ygX8r3mDThcNwl2fBeRtqa7xc2
v/VViJaNzRQLfTq2aogJcxGbU1P9aGmdO3rJw4oW6BDdVlJSH391C+wbDlBcVRrsDPecWXjpkEJb
Cu2eAscm8iCm9bgRSw1rQ7Q6H1y5tt9srkjtokda4hHxhT1/N89KgYZTqyXgO8zKMpYCLvfTTFF0
jQ/h7kgw8GUMI2uzVVWhZ4jQRfb82GaSfvqGeT2SOpme/bwEvMCzvUuBwb+4oPJ6A8cgF0VpAcE4
2ceNqj36kqmFwXhsjBhCz8b5uWh/ZAlmk2+lZP41SbdPTsyZPZQ8Fg7QVz8gc4vJveerULTIw1Gk
DwQgUFKbISyVC7GMcRMmZuWyhTCyAL4xb1CaNw46cKHVht5H43W7JBr3y95dnCP2dLx+Fj8xuofd
pJygBHhS0fAlqdYHJE1UkU48x2Imxe2BQPiqCheSK53+TN2fB91dTwlcwuzM5O3jrOS8bPr347pE
qL9i3cvOh6WeaiUnp3iJKJnz4cmOvRC2mtVvpGoo05yZltURzLmoaiEAI4ddwwwmMRoETQTRAQuv
HqcJ3FLpn3T4A8cxg9tqKKjQJqwU2YChIfVWojXI19ou9pjxzHMfTj8/ost68eyqX1bNikjGfHs1
ATmnSlgXQXqkZ+FVN5CMeTcOElKTNi0sd1khzkgIpj6hCShq7gLPwOfh7JLkX271yeVgqwNJG4Sg
HMaAoO85L7Ko3jAlHcoWo8cKGifsjIQLls1woxSozOexYUQ0KYYLTRJmdLRhsB+xSO6ZNtu2yKZ6
fjlHLdBmtT/g81A4dxl1RmZiT2uXaYOj7OmDI0AwZY+3bwg2ILnVYRF0mnVS5QnkolQ/EvEn8cKv
jan7+qwDImdKMrffwo1FsfMtg89N/fWg6YNhIYhjgyNN7XLmJ6YCZxiErsT23qDl2J5/7dAhN7dj
ESIxo2tM/b1mznIl8drLafzjNmdAh0QYbwZV4tvq4VrgJWLc3sp25Ep7tHEDIqhfBJdU13qWBjmp
1YXhUYU9BLerSrX4a3H7HCu2FzWWCT+20dPpf7YmSxXPp6rmI9kRqgyM96ZQ3AFTzIdd7BPP3lDb
IyYF20/KNQ4JHxHzaP8a0u7j6xIzAsIH3SQ/1hn81OfeIikb4Zx3oEXYEUr32OD7UJg3OB39Er54
hiaw3QL2nmDzfDAcGsonXRR/36lh8GMAwiJmds8fZZVQUzN3LxSBAfeiaGeYVLrjC9I5IGHCgYqZ
XR+rhNCTIp33s7gQpZSS7qStnvc7sVeSQST2oFyVHv42s6GZ5gb1D/Ci/XKID8e00GOo8Fpq8EOZ
He5y2kJg4rV+8+PvTfxgDnBCsDYOLmwcSURGb/SrivVd4qGVOsT+HR6BS11bZfo+hnXS5fkiidhH
ju9lLGeMTWqN80weXhO2psk5ogM741ovkMCrS75K6DxXpgb+5M93pE/IWopc1eFdBCXk5+NKD8AJ
d/7hedb09xmENPEdJKZH/pJvCXrv8Y/diTrftzoAG/ATMR0KcyV0NUYfP8B2e8dthhdaEnG9oLyx
GtRKG1cP04K4LYNT0oqrUmIBtf2Zm851oZUkj3Mz0SjoGnDplnypBD/oszZf/I2ahIf4UFpGqF98
1BvQXqf7VwtF4LaiUIRGF/FpkEvXRxoiCErYh5DwX1Pcg6pB9GT72zM6F0Z/jaFQY9Fg3eRh8Fsk
pResybe1XH/k54zNYcALqNunnFXp4iyY0scTa2UBxBWaqTL4UPZLP3/lUF7pwGeL+SKi8aPk+YnV
LBKTumaPObb77JHhloiIYJprLFkWKqx/eKq6VJutV4SD84BWgxUSO1lXno0UvD2R7HoM7KHDbq1+
osDTOkNkj4P/cbj7GDgEMq8lOJnDHlkjREZvYC1OWOJ8lvfFFMaM8w9vCeGQhIoJVMUSrS9v8FPI
eJzchcn2wS1HHgR9zthpdfOqWJQiWPJbs1cO3B7k3eAOrVP68yA52CmViElmFm8MqAJ2ktAitv27
uqnk/rK3EMuglgZf+U/ey9DWi505Epc3vs+hpmt2Ym4v9YmbpcLsmDqOutkiGVlFUmUVJyUVD1dc
vIwtPouLPkCDOLBxI4ZxQBMsRevdoBeYpHdAyOwMscqsuJxZFAGWsZcLaA6b759pUJyTY6beO1+2
Pu1OLyQnzPEEm+8FoJM862UNh2WlTgzK8F+bJK7620Y3Pesz15CcmTygR6f+hfEWmMkRPO2HJG6+
GJef/jC9gxTbqDcmRoWKIOPF7/X30AuhqZExPjhylx1Xw33hb3s7Oi2MBjxKFEd1uDBu7UfnQeBt
sOcTkif/r3yrNZxZQK1IzvBmuSo+Uzth9vPVheg9dF32JuweP9ykpi1rrFKS3RMytSGezeu95O3P
DuYVW6XwG5RtdC3DPxPVjYGKW09p9Ak3kIXviGS9bpDdAECMYWX2Ul8+OGHD0QISVgCWWl2Wh7VP
ISRPlAbbzl25Kx0pyU8Kj3H6F+RSeNnFa7YJbmEb3YLQZNdH/w0jj6DJUAkD3CYonTWpeqA/BHbi
k127pt3LAClB0fYgUsipsCo5B8zLoyiH6D32fOKD6XaDVUh20SGKbRAqXHG2MaPRxzHmASXEFeE9
moKa5WZAZnfJTjP2IdtM34SX4pAG5XAUw6lpfuJ1UkmtBkVreUr0AWm1rqD0gN6lumVqcghyWi4X
EvVYYqhOuJF4mpu3JL1esXA45eHXn4SERGmdi7S9CNROXkeim1nRnt6o37oppu6pNl8vDTUygMyA
4qFJP5v4ue0JYGbzp2vBHQ8X5FGrBC7L318PBGI85c8KZGH/0Y2gTyXFdKJZYvz5k9omC63LlIVW
9RmEJjJFH+BzQjGi8iiOe4yAncGW2GUeOyZoyaALDaH0jnlr9h0GTS88hXuLZ7d6RTgchmyIhsJh
InHtwdFep16Kk7TnVFyz9OmgS3880BOeqktWIww3DBZYxh5XlGxaDhjWcLC5U8wULn/PXBau84F7
t7Lj41b1Skivhhg6JFCiwX5pPDy6p2LsU0L0EoumFOZWc6Pv98jF0bB8FPn0zkFVYDwKgcybLLkK
TP7xmLGmapFKdd6N/Xwh0q46fsQOsEyWJNs5A3PulbAA/asBtfw28PY5R6w7CuZEkFzkAQPuJ4lR
1lzYuzNP8qAVajMndE6HmP8Yi7rFWEUO249V6LNSQsNRd0tBYNrW6jMDI+ZQ8ryeabvLMI3hFDl7
COV/Bd1pe53F0zUZldXQ0NhDzufCPS4Cc7GruhG7qBt3R0Zyj0nTlPSL/cJLmslabHCN2fn97x7A
N0OKaCvcsLTy+5839/7uNRtIKibBgh5fVzXOLJR+coEABhsxY6ZUkURnpCzRRpZAe4MnvcKGPEFP
mHo9aGQBAezHqatw0HP5pDZK+pAOxr+HvRmvmf4I+rg6riANVMYNVUXPmGJRcWlaUUHSpEpRqCG9
/vuh/xHsCDpI67q2CD6ZG4JU8h8WUJrmK5cmErNX6YMfB+Ob1xPmY0imPeQjp5OFrFGbrnKI9E/V
6iU9EHC6KsOqgeVBZQ4QRwUNM+OMIbrHIiUwNwN65ZyrLfiprLCHdNH55bDjGMFoRTN2Gh8fuxgW
tyM1iia2mibaC9o4S/RtOxtbmg1r3VwcLTY76+xSYeAMpDJ/bgneEnzMTyk83n4HLDnjV3Uu/ZL0
zr43NMr2VOmTGAyYFG1XxmhPlGKV+AdjkGRGHFrULfxuOHFBpP8Rgo34mtwMgp40dPBkYVlmbVsy
L2y2Dxn+WU5N6ok36JsEo6ucX1t78TC2jR11xzkJhWwRUpj0k1ZyCmSUX7RiJovY3NMjg3NsmW9y
ovoEaPnxi2+Lo0ppVjtvnhU983Nk0fUb9HZseYCEDjrrWr58i7sfF6vtd4fCy/xMXCchyJ6EMAqM
dz7+4j6bcf+lPW0nQV8ZjKx1WpQ/CmuHHG8jUiq20cL+csAJzr2+p9TFMe4M0sWm7zgthGajm9PU
9p3mRPzeEoTvDPZSl3ssC9sa2q2jZ1DXB+gkh/po77RZb6QJaMNR+p5RoypEMC3zXahRDHezBP9U
QVb6IfWGqF5LcKyLsnp9ieBUmWI8eUpyOW04l5EJ/Mk0Gw8P4aH669RZlf0KB//dMbiASn8p5i+C
eQY0G7p6tyAX0XkC5vrwgSyEHX9PWEQ7QW9b9+zCrjJ9CdSIjcrZ57mv2AfFu74iyCwSs5OMFRmg
iVM3GWL1f4HmeHvE9YCvVbIppJgsOZvMBHKPlbAm3WU2CpJYCX7Ub3dAJPbU5/bwbcJ3LVeOM2R1
9sUTVt3cqRRdUVuhoQ6xUgLkL/wV3HLR4xezcDw9xBHu7eLbhh2J5yQjIQkZgGP8ct8HDuYJ6Vqd
tLJnabFfii6eBVjH9dgWzH/jEAHeTbWS2UXQ4pG1sirIovM7yZvQnq3bMWhjqKWhsgr6dzwGvoOA
Bl6kclbh9fCVX0euLZcMqMv7K0P+VqtRov88clXD9PPSIRYbqvwMopqK2IFT0scEv/o6FgF+6u1/
nOI5zcRC6uAO7Ia84tIVgJdeDrD5SO5XADlIzrezSRe4X78TRAPoMpVSV5FYqaCOqtzOAc66h1eC
YVQOJsXE2Se/z1FFiV0ppB3Qq84SXJ+c5M5D9Vkulpjq9pvuSE29Cns6Zpwm/SaYI0v1Ra7w11iC
KyivCrFb01LuDPZthq9ybw7pbPUUc2zjN30HpqM7Dc8xBhE6kgFrU0C2To68vdtqhflY88x4dlh4
O3SSzzQJSvcs+AdAlFO72/ETu25EpAaysdxURcy9JOpIKiPc3UoP3QcWuWoOBYhJbA+wiEkEOUo2
w3dxqqubTRprZO9MeuQQKivhG6d9W/3vsENh7LFJO2lc7UuyLu2G9kMbn6g2ZMagl6+EXLPWg3+u
6KEmwlbjz4+J3S9YFMfjMkzRQElaC09Oqjb8RNEzWe34wTcOQHnIkMX2Le4n/rPsad2SyQCcgEI3
l6Et9EsKRRT/5NZvoOWEfiE1ajxWI9rp6t+CN6/ea/Xgbrf263BKpLlwdKV3nJJgO3JxMiNYn7r8
FMjYqHDemTPhluTh9/Pgh6k5GhCDpkhngkzZgX9rbPsnZq6HBabc4m38GBy0NPfQip1VviS+hFBo
EyfW+BCDRostnA2a1sALsPbN7Ns3fRkrm+4zkW1k1VcMth9wFRzWKxogK3JhPxwaKOydU4f3BBBs
CByjUZUK49MDtU4i4YcAav6BqT7TtfXvYZxbBoH3ApbXYKnRDTugfvzSj0F9nsVzYn2uLzUuB/sz
8AGqOfyQ4+Pd6VCwKKc0loatRBhoQZtCS+sLeZRNv0vCiqwWrvbu5PDrHa8GkMOURUumSmFHI5Ya
TnwvMEB6QdKjeaJm7JLd3EGl/nCmLvW6bpJn6Q560WGq36EWhh+7CnTRkNjtZX+nmPZeCk70v0CY
XO5938hdKecT8qvPLuC/dtLK4yql77ZUFdRRGfGiFoyKJ/H+vD9EndCr+Id9eRci/8a8p70/D+a/
2yu7fxdoETtz8eerlVoSup/Nsn8kr7NMUfkSMYDhptRAPCOfYKRwvd8ij1mufU1PYFvnFdO7Z1U1
bWkkHv6wqE1i5fQPHApD6/4pfGLRFQSNO4aDTfUFyv2YKUewzpoi23eGjlEsdgRNJ6iAJK0wWy8F
h6WNeqrHS/mrkxnyyp121h75dSZ53Y4jMvNv2kXafQ1YuUXkdaIFwBGPXyfBfkOsAXtufhyu3xJ6
9qS5zj1Sk1L7Tc3A899WdRvtjco+pVeEpGF4JxwhG4RjUrBxoNjC2jzaUeaGr4rDwJ1XfgMRKYpc
w+JeQ+amz9TDOwCYgoKsw577Yx0nXZU23tJcrqL1CYBWb1LSmSklzI4XAvM+/9e0UZmFgLagpew4
fSetJe3ROPpsgBqRyaSgFJ6qTliezsEqnNhXEM2OEKNvQelZZeUXz5dpaygh9xvannZz8HCW0DOV
IWgtjS9xLh+QNRZQNUTaFoSVB1U7c6Uvy9p9DfhzXv5Veo0CrFcFFeDOQsfPTVh3xknEeVGhqmnh
iRNpA0F1evNh9A4Q53+t9w57vWUsnCIR/z+6EC987IDhEGQOTWqJDeuw3epRfuK9n5BNp0TGGFzG
TRJpxVbk89kK/VQnekqblS66jPjGXaHlIRTBj2/ZZ36iRXuM7oUjJ/L/kvSqR/hl0ma52ui8R74Q
xSjQTiPMXEOcLVuuCkaTCiviNB/SuYt+EgEyCRmCmjSrcn5P31TWfClypY4iet6Qt4yKJGFrA6wN
GoSlDlThwk5zPiou86UyJmyN0A+Df8R/r2NElgrG7HAWX1b0JKG6wdNrNu/KI8M2bGdvX+kiOhqB
RA3220Kr9++v+DDH7koP07FgZ0kotvoRgAJbDzUJL/h82LeEo3wzGu58G3330bIEWq+rS1zHK6gA
0elytFjVt7FsHjOYkGccpIkn2IeBe9Sx3RHJm0yp+3Q30RbRgsb1vmhM13eCAnhSTExKry17eerN
wE+udWThZ/Iy6peBOY64Xu7cttV/EsC3oz6cOj3cmw4NKoP16Ln/TavdOios/4OtRFO38YBFJwZ7
9QiaPnfajYAtPNyiD10V9VlyQAJyK9JUK1GUYG7KLLDg9xhN5EUjyXugCUm6IR+99AXfBsVqqmRQ
BiA/H2gJMeW1/h14N5mmNNuchLdYhlhvpgqCz99Y8YGvGgsUDF5RzJ0r6Ld1Lmhz+TsO6pVVyRpf
WjxRgYtID6DGScnkwDk8ZjTzJPO1Pk4IJMy6FcoqDxN9TgupjiKldIaAi7XW602ULowG6H9PufSe
Af138hTOjor8mvq3GhCBGZ9Nk4mDcVDLaAzZg+kCDOfmrd2uwwQQ2K6geQ1a4zUtF+vdcDdhBJzJ
HAD2vdMQ8dtQAlqwK/QpMYJhoPpExhzXkpVJt9w2JV23iJyeDJSa/LS4s+F+Wu3XaOvCruI5rHHC
B9V/D1c9/eyitqIFZhb7tTTxyEZ6LexDUdH6NqFq1eanjkNvxexgDHMHqPcI0n+xMA/tCCuFFKGQ
R/d5Qyopjl+3bXdIR21kuBmDVyIymNB4+2T4MMnC4h8UpHYfRMdFRfsgPVaSn2P16RSFYgUpfxuT
GFZ+JD7qtLPC0MqGc1Cqrw85RhHw9jDDET5R7HgtZxdEfu9w+pr9YcarExt0JB+ZeomEQIAbCur0
M/wHPv7HDTLH2o4jHR6KjOKwktzD1QRJIHzMudGhdKCrSOfURYkDF2Wwxba71fBlLuS7mFnJNWJb
J4ghI/P89rDPpJkz3AoDjpo6RAfXPWzn+Fd6DT86VBHwoWmxXS7bh+lYyvX1IYgkGM4bN6Yrt3qQ
0WRmGdW5WyaPne/2zAIBgBqm2zKvJerqyVR3yA4JESbQgupDZI3TBSUP+pprWmbX7sRddeBnfDk+
5s/xZebTWOQKy22356JeY17KOzgZa3MwbtrX/cwfptLM6qLdnv3X0l1mJEDjilzf3OGaKAPiuIvA
bNQmbbc/gIpc5rgk6VYQCLTNLPH3EG7ENZL+sukzSmI20cjiBynGvccM8VqiUdBb9rYXIuEHKjmA
jzTFKFy6jqMXByn54NGVBbzXCAQX/JSKuaGeEtHjMIew3s3tcUre272iRYNE6n+y1QQBwcwVnMPu
H8gdbj8KVCYNewot5r2Y+JYX4KzKlcJZ8Z7iQFFIlpwaDB/DQWnxS1EwO1kZ/v4STl67SYD+Iemv
VNW37ZbgAoyW6M6JAGbLXJraSqCme8F3tMieeY2SxMuJGtVxGC99krqeWeQD5tOKTabw9JJM6Guv
zWRaR4+0u0W3Kv9/X+DSq6Pol8QzrDP0oStu+UKMwqd5LOkpeqYvIpubKRTc2I6f+skgHZAVjpDA
Uh7Z5JfOndnWq+RTmoJSGxSW5MX9qRYj3aAcOw6har/sjVK3jPh0X8PaX+OTkiAyS73bMA3DHcFV
Z/yu9xyEepE+HLIttdisJdA8xTHjB26v7rPpE/l2d1nXKjBP0I9zfDj2ORLnPekd/3OIEJN9Eg+N
8745t0RicEypr6d6sHnJYQlyfAspY1JHNssEig0XJV0zdfFLCAXTaDJdYGVRapWsemvP3ItUdYwz
4eRC3Ig8nnRmh+9INdN3HqojWLJGGblOODwlDIBxAVVOLok3ljtQkFSgSXsXYKScb5unR9WLO1lj
dmKEfQp+JQ5YDhwdAjeVSwuU1XrlQ0Yi/L3n799L8f3EBoqK7xvkJOyHeKzuRGME0DNBnkBlZ+NQ
3IE268thArw3A1C6mWT4l8YwsJohAXl9kJmEsoBH+nwwIrmDkRWXxXZlf722oYkiUyzqOKDxWbun
ZsPDp75wVKTj5xD/s91Y0VIBSNCyKHO/piymGLmCH3IT3uQb1Q2o7v2n9rG7DAWRH8tcixZgzyLA
0y9PgLD2CWn2VEJLDTWY96ZA7gLZskc7Yi75xMPP2tEptR+RHp/WBLbJIhT/I7/hS8Qy0qLeoA0c
TLV7gmqjAcPpJwBLo68czRXC9/4KlI9zn00yZl1W5G47OWTVYskViyCqPfSc+8MvyQDEM54tOS8X
R+sC2L6lvGOpWcjmq0xhAgGQmpddjedtexm0GM2ln6m9l4RaiQ+3Slp5Z98SLgJ5tPqrdE1+QfHT
fOyfzq3ffV1DMecutH9laOZ8grQ04bXV41z3IYGRHtWzvZNjXj+38VO7dH1CpML+XG9F3h2SQWsY
bQNoKrE1uj4cbPj72L/aZrNdJqy3+84MbATVd+itSwWv2OKTUs7vbdrTcpAh6W/DqRPVGGNESItM
fsvRR3Ght5gSybdTYxdKHz7pFxwnk5q9kS22DhnzCTbOFX3zCLz7Xly88x8ELMMChH3rhsTXj5kF
fI97CeJHmrkrnodXejnq3svO0v45HyZPBNHtYdLELxUVoDs6FwnppxPYiFsyF43UTyNpE25FEccC
cTDtc7xW4seQIE/siM3iW8VSZBpa8EFkbjagFE2otSsPjYTGxwrK71mSjk35P6RQ92QVmMGhAtJk
AXGpJt3UW3i15VezTAlueCbUpbThOZMCuic5rxvpsUDs/tTQGDy2KUkk4ecsPVM2t/hHU5kvE0p5
a/DOS+e/5en8Nx3onoh8WV1+d3qaJmc8GTOk6Qk4H1l4fSizJTsqKSRPHSpzCrqck0P9SiauOjy1
NaF+IzY9xEnY33QQOFlXyWVVMB/6cue+UaIFRiL4WItqHuhWVJKuQfhJ0tnCQuAXb6434cf20zwq
04IfNrK8yFdmATI1t72FNhgfYBgpbTRTw7F61CY9ZJK1+cMBmRhoN/+debAk64cAD90/2s/IEcJy
/9reLFDxGHwImmK47/sVA9EwOP/HWlA1yAyPYyjhRUKPAS5bTX0hvcKLcRWO6woRx6qdh99/zX2b
leGQ3dANuHjaVHWnJ2Dm4UtsBOi7b+35BBtGnU7i9QjYzKmBlar4oXUmOmez+gTiMm72a+eVyNBs
j32CubePbCbnGZEwkTcKvcyHg0y+lAcZTNHjfUiifJY8YZPPF3xCWYs3BTAq5pBAan4wrDdcbKW5
cE4bK20HMsryj95tKwVCWGrJ66dscBjpAeaeCe5uTki4PfVo0dcRUCSEb5lnKtwIqWCPeIyXTIq9
x14CDJ89cvXg4/wlb5CZKyv3PznarVJwWoSkN/ueN/2ZGNz7a3/CSoKzRNiUOvZxEBpNsvti3I7X
fMxQbBCw9E/6l1puKJwEaRAmC+D+RqBd1/pyUAsTNnrQ3TVnCzkBxaz4bNMnRxp7F8dFmpMkyRdu
0K03ViBJqZoupQevmbOl3sP85EexJxhX2KF4FfaO8i7TBrfw9guOEGKU6NY0eUR438h+OfntDWy3
p3Gvnh3xfbGaaTnLkHdOZRiWtRxGrWyuihmQA2sKhqu3xb+Tb7ADQjBjvivxCA8+Y4j0BLTUVCcl
jTULdXcVbBKQ9Qv3td7l/Pjs9lKWtztasDrgvMZInQFyglkPVWLEOoZc81uU21un1UVVF8p3M5HP
qcF2Q947rIAasbiRRJK/6bYAcHXzb7R2Ieq15Ke6EO3tsLAFvKkTlalwRo24B7MPE2GiWudbwkmL
UDIL+9X3Aerr08PSOtwafBmNXYcQnrvHhpfihc2PtRnIaINZ6pN3WyYW6PJuC4FxgitPy7i6L+vv
3wtoupmBTA6rfBNqd59gMLy0H2eHrwbfrMQzieVXB+3ldYcDMVWS71c+G5HMImxs6ype5Cfzntxd
2BOFWhudfSMEZBUNrXwvA6k+9e9pw9yNp48kVF6egq2gx//N3UtBNGgKh27IhMAa8B7bqNHqpYT6
Ax8Aevjx57MymL2Q0qtBD/8d2YCdNR2LZ9KL/72OsbLiSQQ3ZGkn8qQCX2fRr7ibnrcQ4VSfPBxb
oP55apDnNX7/Sgiwf62LthBaM/TkUZ2fTrxh9t0Tc8GnjTaA8ILNCjbNQ5WLlWX/GJgAR9pyRqCp
em2ffKPBvqgIkaVjOYSO/gE+zUZV5jk/s372NIswJyrLWFNu4buJ8VUYIgw0319ayW29hdAK9may
CStATYWz/MO6EWKKUOz76pvVDsnjhApNkivzgj71vTco+GJeOaZhjSEenY8BkUAJYo1DK1//n4CX
GS7CfYdXe07uXCIwaMKzvoCyNQvH5nKxg953/3cXaCfA8Swbt6r+bTKPN2DuiffYuJ2BiaOTSleE
nU3M9M0oSOlJeucH3wvrMA+E8KvIEY10opRVv5N9MIj3JdCKtsKDiUVSktGzly51y0LVg+F/9kaT
xsxzrP9u1EHW1XVKccdANpcKENWHvSh65I1FJhuECXu0GhDN575x7YnxzL35eNmrqoS5rtXAR9VT
rUWwW6TX9GFqMhuHv71yxY005oflJMS9COwjSfU84TzLpHQS3IWQ2sjRCkauCj8ot0BncugCZvY8
67HrOBtLVRHo+O5TPY6DpIZSHYEtmrfUoI1Rum0mLPHkC5plWKPlNStqJaaK516DJx3Qt4aJk/HQ
QQN06qrnHappPpwn0AP76KqeWwyfQ2bNpjjWljt+t/Zmhr/xaSG8Xl/OkNMbXmkF2WItQeaXcRpX
Agdvs3//VUu329p78MqCipqEJlfnjxUcJGlb3O+nZjQFLlfKHSmoRrFvxxufSLEbctOUiqaYai2+
nW3oR7329vIcQx1hYLG07/llFIZCRbAHpX1yDef9U68MuMDECYduKmihDR/EYi9QcIyU8I9TiOkz
V4djtel5U7wCsJvO4J1Rmr0nZuV/a958YOUSDXwI6gX3h1zYQ0OuSc2PDiqWQa93JUqbiw2wCojr
36vrwIZBmBEb2HOC5S5jIkLapdfAQjqJFJebHkl2FmIvjVmsYAh6FhGDC8g7a88fsWioM0qrMugj
UT2XP6UQXAJPwzTEAZ6KmqdksMfkz7V5B8aRFQ70/l8FIb261L1nOjvWnLLSVxN34fMRpldtyKeP
StgIXNqx04RjKda8TpDX7UF0tifEyBz+zVnJ113lhU92FPc1MdSgAK/WvwDH7RDqbncLlHkqfa5b
obZYxS6N7iJyudFivF71Pu2lXhwcNo+2h1Qzx7Pq2EzZPVE4fJuWj/ffBVl4ZngBzd0/8JHgjb/m
43myaKwA9uMnuvjjnen6GeCyNoWJyQV0LtyndeH6eLUH3T5XOjKAz3uerXAX/jNfTwhmdwJQ9XpH
nz1x5Pf5BU582yucl/PnHhMdI+7mIcwBlqhdk266r2iOVmr9Y/FocD0qmRkMgQ38kuTnc/Fdontm
OOUvgmTn161zGkU59YUDHtBVdeagC/FeyPALiH5JgP6ZjVoBsvQ3aPFfSN64ymKyrQ9DuaDrADFt
lBL/Yt21OS86MtjWMZCpavkYEbroKCmIkB0mpikq6lBJ9SXbHsm00QZTtI+5OqfU33q7YILQsgfn
jvctuVUqGd8u9DleeojZXR/2CLZC36pW07tPdvGspU0yCRiiB5iSC20lQhM/FrH2I9Sho+uKJrwV
O5+MZ0k0ywttmyGRGCOOFNF4nKifelk+CRO40V9Yo3KiePgS/mXvuyRZrYlwEKrjtOsINAq/WzXe
Zsfv9EFDWL7nDUoMOzWlbEKEs3IOVebVcYk2QuGz3a/ewp7UwF8jI5iBZG/rgaXWVaiUWnmEjtLU
NDKFl3sixehPALIo+oOeB90g8h+EHqXYenv15i8B1fao3JH6HNvewyvlm3+trCn/wTXSuTz7EIXa
MQIL9Ffyj4JPwx6qwei1WXhLszRuvvbkhLrBeZf7pAVlNYIAkweEMkYUpFHK6qIHgYpVf7htfWLV
tgE91z06rpoc58Zef0TWh0NrsqXmQbu8A6eGv5pyLTw1SBRmIH1sJeNdchijLSs1S2GqzjE7Cz6G
AgFcEIn/l9oGDDkWB1nIyND5szdTpVrJ3Css09o3S2voHDLUi6+zdHxV5qywNONpqqlCNx7lJVMW
HVyAmJIkL/0XWoChj+vh9OeYvbqOjQ+l+FXnkq7x0AXUtO1tAJmJCUepmXIsLxja4ZMDAJNI1QCX
dr8hBTAsbRYfeQGLaVqrdoxuUGJUd5uswAc+iL//pZzdbee0W+HzR46ulEaOB7XcCjmggppgQzCK
kYLL4jQCKlmhEQewwD2eUUkrDpCcdSJR/jacadJginGPsNhbgIbvS3j4B2ljcL99zpS7zc36d41Y
NsixftTbpndlXpB19Gxf10NS8jdrcVrPVpWk2g6Dp+8yLRvOchGsPZgB491ie85NR2sDmzwP0H7j
Na+lF28ZlZasBspvwIQGyXbSuBMLwqrt5p9ht5RgslQVeu4opL8qI3UTOwFzBmmy3LgOD4B//GmP
x18QbZ3u8CqmomlZwfduuc+KGSwfN3PKJTyzTowANpRa+QpIYqAFvgYbbFnKE+mWeOs3ioDAurG1
CmGTSnjJ4+Pg9RoLwiinyYsoBANYU+1vOVMiHzZi0371UeERAXXl7JpGlmvmOpaxnaS5HV4nZxgE
WtM3rdd1Dm2UVQhDEIRfnPi5v5YqfGE/I+hegKR/UHrW/ug2vS9VhyUvq5tHtAcNQnhBR7wWn3k8
+d9pvHFmJ67gvt6KLHLiq0fsS18P5JRJRxCEC4wF50S0yaQXFyyHn5YHQ0O6IPQbIijP3g9T2VNF
Bo0pZoUeaTVVQjU/4j3wJEDNvDpstJa3w5UAT0VuTVYBBv7N6Vie9ZpR9evsmhPqXQTJKYtayH0S
Q95bK/2TqqSajMx7Tvej2NW/wuHuJY1kA69dU8GvdqvhXxaVwxP6phY/CTBSzzMRwlSjLoNeKl8g
nU6iAcHS/KNf3LeDhHuS9VUkMseLv8J17Owt3AFh6pcwdaR7hXBK2OLopzwvU+JV6nSufmtUMUcz
YCzcfnBLsulFfdT8Lh1OtkonHNKRgXnzcMc221B/7VtHPRfCsAz9D1YWtcTB57pOTUhHbiUx4j0C
0X+fAMpuJFW5zgYmwFg3aeqeV/z+giUoxshN+eWiA2ImEbz1Sysh2NuVw3KAHtgFYXZmn//BlaBr
8FbsTVuTz9NkQlR8vSQREDF+gKlscFr1gg+cc79rSTvfRwppi5PMemW71cOatYHu5Uq+gyStFvCs
5FOr0Xq4JI/+epGBoocySRw8/mk4iT8IGKL6RfIXVSv5JG1A2v9i9tuoMwMJDgZhJrfKEU297W4u
DHiJlkYjF4LL0LtCB/aOzD+mEv/+vuJUIIACT3v8GiVVRQuQBaRFDwOWGodgmHhuRO1B55/Xoci7
eeKfilNVMLm+Qlo8qDA8RWJVFr44YqDPVSh//6bKh+fWCw97Yo75qcegdX04F6z59PQlLhSsy7dV
3k9ICQJqVb40v3XgOer7P3MnGONVwPaxaPk7WmKRTNeDbxJIdD7Hewn7BPTN8w+eH9QGzxFN4gBp
5l3KIOwaLn06oCLZ3YsXjeBzwUIGfsvt0K4GtlwL7/URZn9QpiTBqlcpNw+9eI9xXLg2aROtMyW9
2iYw1vObOTDnDKPUkNHzc+JIls/7SfE4LCTKBe/BTPWZFxKJ9IAsKHyho5M6wDmiJYqNdfZbm9F8
6EwPOeNlAAkqGOlyi/8Y56YLBOIMjnpvOFLooXr1qHK66ICgwdgeW37+vv6Ve8f+7ev+EiCmmfxT
3lAt4jQwvpzav6n1qpKuiBBxal39IFTx57PfXJsqvRyDG2dVBok1NbIBrogNPA1+AywO/m7cCmuv
MTXfxU5gyd9+EmCQ7JoPhSvAwqiQ/JaqcMtvnAazsH2UuPIyahQS8sCzEeLN8yUTg9K8b4RQQdA/
NECxwtXnUUVr4WambD33/EjGqAS0lsc45CQoxPc822hFuu7ZXFefzfV5Xgug2dHKmfJsTejUEsuh
tnNRZkPHSql6/4afsjmMQB1j72X16eymluOkrzvTrBEjrMhzbF1ay/WhsgTTr02alJPffCcF5E0D
FD26iz/RSes8m5/rrnhJykvOMoACIOGscTGKYBzIwS2T4r1wZBC1qfVfXtM8EOl/u2gf/Z4oOMNo
p2cDMKygQ2g+TQkRR5uZmhK3HOXOLk39F9PYI/KzrTvG2j0i8ixvxxKfgDQRjSui3d25+nhMEqxa
AyiTyj46VszmZjZJ8YCN1wFnR3ANCuuKvBIbd+SJ1YwZVwmoZlEuCfgXy+ekIpzaFucYUmRbSuMp
wQ/Yv0SiOHFELoZobPFsq6VXiWYy1aJqyZrqkz9Fk14IGjWsRvU/eCRYBpHg24yyV432zW5zjo0S
ZTByOCy2psOw8/5y6oLly2fwUUC8ciRHRX43Ae69OtcXF1V0WO1sL8k/DvMRBwrjsQM94roibglW
nYabm94LR3hDeoWBIicD7a/Trwbu+jvs6zFH+XXbHMFfVQLjg1k/wJ3f53Ja9zmmJhHQak0uirVC
zDMZv4IJMSh1ENK5zb4awFlE8xt5TCtSDIdzEiDJbUmF0SDY6TNw5L5mlUUiA29pX5TLPJbdeOOR
8kmdMGWDEY8VXmH8VJKDjFEHkElidjv4WhFzVkKsvVJNvGjVx6tydGgLDG4LwCrntiWolUr6iS5g
URJZp+us1stCZZH4MqFJv+Hfd2Sl3D5PpU2aVCVhqguIT5dvuwAW6l4UfL7k0w3pwYfCQCfwMPhC
5jMkw4Fio29p8b4tGV+Le9w148sIPcdQ7ub+LLqfXmVJWQ+/6Br2cuTqAr+g9KFIz+ORjUbjDgy2
s49zBQ4ARVBfewYX/i3PDOZlTCDadrQ4rPe0hhvNJUqqAvhQ+tYLFt3RNQLNeLdtqGjdd4tdK5R2
K6l4BRO8111zorFhZZtXGo1Opf8nyW84zR8A6M465dvxfkZG90kbtkyxZJSiN6OF8zOB80GdZ9+o
+WCfjIS8oM/AVkxBAeVD/PtqUwMHRbbFyno/dTZH4b39qXMZi1W4mH+LMM+65lUxDgDMRo+y5qxj
khTPtyD1Ig8hzpe0RPYeWRfSTiQOxb6ighHVh5dfz2O+1imPJdNoJFccndBk3jqWK3Rqas9nAEp1
CPX71+4BaayF3PXlKiSOsdrcCoPUslFx6ePX/n1sOIfiDQWNvc7syNgfJR9xNxiGpSB66X7ZsZyM
nBXcbaiVUtszQNLmf/v2jhhxzfrrDsc+dkbzADCV+cuthLN5xHYcaHFT2XQn4Yff9zxajxnC/hYy
EjH3B1CxgbIW8KJYXZq4XNlCmMGZLslLUnZewYfvlJcD7G0oldtn14MZtg0mKs4q0BjYca4k9zS/
ofrDT3+/Vnk2dpZcUCQZ2fpPFCz7pFP+cVbtobZzupfAPLN58fX35gwNQc4q3P2dnu3j373Kru6i
BhCHa31u7BOI3wkmNEZLQonkA8vCl/c/bgmoCER17k1HNZceef6t9XBiEXF8p84zha5BRXXbImxc
/NYoMWJY6582Gbc7D5XeTvlSqq3Qv95wM4PKpO8QofbDx9ooD+8BU2SMVEM5spZTxDEGQrfoGGOa
lqvzUP2qRMGarO+7ypCCM+5CjDTcQBnwlG0BNoqw2RODPigFFIqpw4RWboZ0a9XmvF/YQtVses+a
NZ2G7fLyWM+X3u17J6CalF1xCTShu4ihh9EwFPJ828o2XFRn6z2K5tUQl1KAnfTd4lZen0eyj7vj
pm3011iKIg+h+r/CmuLXJ0rOxM8BCGXjVtm0MyHEkDpUjyKp8b84CoLAH2Vx/F5MwBhRgo2z1Sbp
RHan0rf2m9gUTKuCkIkn5tZmNoR/7brhVD4kNVoTFamZpp7FLG6UtSU+LPEWDL7uOCOqKAfj28/B
DUZsPD51MNHRNmqZgUTTfXFmBaO8AjXNzZRM82iqRltM7oLNQl4pn/Ocg7BqNU9hnUmHlmJn0Xaq
T7B2XkJiT+AGXsAWfKrJHyuCNPc/F7NIsu6C6gsGixDUCw7Mc6oguHx6SlOZ+QZ9QdkoYOrpJKVf
62gAAzn7EIE1PxXagWmiskzGWmqxPhEdQNzH5ZeLzd3usHA9W1UQcytV2Jt6Ib0HUrcHsdqhLF8S
oDkt4yGRrT22spZZyCRNQkyCUttN1nCP0TM3q2LYZvJTR6EuTX9tCuWLgxl3Skf0mmob4xa8vKAE
MNiGTfOGzY98VmkXz1DUS7wmL4QsJrBzOayrPn7TRoJqoQSKUW8CO82gLQwfK9TDgLgxYmZWT780
CA7WVm86sBNVcv0/UeQm2v9YvBBu1IEzFNNJCPseaJC/6EGjtkqTN88DIkjgwxWp7Nw4zajmNG4E
KbHcIincJS/q2DfAq7dyWYncyFs6SnyXVgcGzG9qXNsR0tagrLAKAl5RJW8FZw7SwRRECTic78U4
0my/J0umwphczoKDG/IR15H/RmB4ygREZne/AgGdWDR7cBwwVHWfgJvMcYhfhdZBcLgXjkrkVIQf
29RUQfYFYdFtJWgeyJXjyOpwBO2O7Cf7jBOIMxxb/InxiNVtmT+MCbBjJ4unsQxUu+6Kbml2P5fZ
PnqZESVfL4fnyarSQPo38IBC0P1+ZJ8+aL/4Q1R2Zsm0Cd4r3yBbNquKM5VGlqWpHRTcjzJPUTnY
5e1nGAUALPAz/3sMxGTf43lBL9KVmiHemz6D7I/sxawNflTL4CcSPsRXHpV59VBDM0Cmp/3GWopG
lqcPVXxvlqAV28ig/6gY7iwxIHRok1T+qfwR3YpEDlnDqvs5iMMCmLmrgsgg2dmpwrtzCKYHhrkY
GTFuz4pTjfA09RajbWw0xsU/2bscyxb1rk0MU+E+bX3YalmnTh10a7v6GFYsd/kZAipeb2O7Q90J
VXvgkFPPEcplSRh/VRiW+gvXGX47HOsolmPZMYD8fVg3kcKGbo0/8AzpoD71JmVOdjsnz9QMQaxq
ILyzsIWHV/NNbaEifDY32PUxmpVQtOgVJS/Dhy3t/oH7FYIEPrCKBUcdLQ6lEhrX93R+TEMkVFht
xbIgC3cOgFmpcGGmluaMpMceWIGzE4p8JEfHu7A096W1awrMVzUy1kPioA8VfwLnSjowHQYKCnmL
4uMlz/o//hqwnrecmrIfxR1nNmYyPOJGjPGsfVX1k1RtcXTW+Y0bi1Ysz9JevI5HmE43BOuY9kR9
d8p1nAAjhk+LG9oPW2ngMJjfNgIOM5Z3O4KYNcveM1L87x7FsFwOy3nh3ucOsyvRXxg9TuHRV+mL
I+4xKwbVH+qCOyJ5GCsN8BpIyu/x4yM9Ve8aj50LPt8kAMJeMM+vfWmK26c/w2Xhrtp7qmC8D8Qn
pyf5Ic4YXGQ491vboQOkFBUY9s8KKs/Snd1cl3UIotvwF0ujpakrtwMF2XuvFwJ0o6cOFEqEJ4k8
XzA3CDd/lXbfIJQ5QIcMnAMUCbsrlA+ykHyV6s7odqvLOmDzxk0xDbrQVEzGDO06LRftRIV5nG3Z
D+oGXWttSkYV/Bh/6T0hYwbiV+WazPRbglN+GP9gw+2IedIEJo5D44EgRejOLtolvlQBdJ/WKZXP
D5OiY4QsIh6JDbTzKzKNKC5RdQwH/Z0lAngs/gqrSfbg9Udsr0gLelhE7RLe9f7QuGjebyQy4C+e
U33NLQoYxxopDVBU1Eo6oYhLwvM1YiXyHCRPEkipcRZtcxeAfLA+JqWVI8mRt8vcL4q6ogvupN+Z
Qf7G+lzggZPUej7Sul/GU0g0rVL8I5mKTga1nYppQtpRjvkpSlXylP9f/NOEFOsFnGHABjBBcpO1
94en2hXLppxPhqWpwE7VjsScaSntxrK87dIzErYoqRDebX4FZr8175OHqpqwze0J1DCaF1XsPc0d
hghi5GS2VhYs4iMcG+BcuiVdBI3M5GfzAdAKAzN4cVJ9BajJjQrOlnTuOyqUkz+H3PMA/1tUTpo1
KVcoKhzkzxAtxTgwXSt1TtlWN8zcJir9UgzbKaguQDteeeGpOOnytMYTrGkOjEOxbRB3bxG07cSE
8gVgENWetMMlhFBOUs4xoqAmqmfC31naSnAPAh58GmvptM8UbN1caPQDnlKvYnzAFYbJbtvKGUAT
89CCKm7LSGlpISxojtizFUhgKI+vXHtlrh0ks5YPT5nYARvSxSEkE6XDMW1O3ZgItdLr36OWYtnO
udgkvqAorkBQB9/FhbJBg8UdAexjoJtUW5izJgQ8LK2LMem3A20ePgMJcZGAKhrIBaNocNb7MWNO
8z6k12vmYI0epfAVLJneP52RQxYbQd2Sr4aKYdLTbROKhBqzc7/Xx2CH0uoFnMIeq8EBCyr2SG59
wZCSafiy4L0eQnG1KYgdPQbUSqtdoa50awM65COcs5YSxGCa/klvPaFeQnh/dgjX6FOeXUWSygbZ
JjgR9rYGnYolo7Ns78wSDuY1jZ4a5fDxblBE9NszUjuwP8Tb8rYiGnyq6juJelx+h1L0gFccg3ic
WK6VOgKGeThIgyTKglytQOG/i9VUoTqzFfkAN4dRAMi6pKNgpX5SB5D59ErxcFd5hlPEI5JlHpPO
4qIOG0ny8vrppWj0b6BsQ9I+XyrDfg1Wfebdoqfl9QxLvvFjMEYMZS0pzuSMoap5dR29LB7Q5aLi
NqxFG7plevGhWcxU11XZvLMSEr+Gq6+Oz66/MuVcdHTZRGG1xlLFBCIwHzLIl1z+m2C4BkbZsjr/
+oAypr27kQYhBFzGGrA8eNQy5YsLpC673VzA/9bUuVf+0rhKt+L22tPYSZGokbOnZMlurjvUb8ES
ys3sGLU/eDkFbd5TULrGRwY8UJQ+1tHQf0oxi/DK3Tg8v+u0oruwsxxkAl9V9FvKQskQKHSN0hjF
ctC1BQREZkE1wZFXxnqseMC7bhb6irKlAB/kdxWo/44FN0kvATuxx+t8sExIFciU6VlUlqu8fHkN
2AVtChEY1qu2ndnQ1ZMJXUq79kUcK/yu48Ns1ZbbV025fUoPIhVsmLmmwrh4UYEVaFBMEn7KuwII
gcV7P5oNoOo1iwrvaxim7FcbwdBog3ZPvQ8SzJMFEIyUZD5pkpEQvr+PsE703qB7iHdqwsYeJsX4
jKfotqZ9pJz6m5P8N+rScecZIt8hey5GcbcSZMXmUNcYMSRQMyohG7KscUkujZvy1SsK/SovL1V/
4KJ6ogXPXSpHRGegpO0FYMcYOKIzbPKMJ1esGg12eojpk5GclaAR8N/d7EmNfC9Y3ZpM2pfRcBeZ
BqNYJF9DmL6rwiNAhe2MQe/A2xGsgDUSkzx96oHSVLn6HI2uDOBI1wMNkIMvjSPMWsbJtDFe8dMt
mrYAyNpD+eEVlMD4QVrVfdWzA9KkEpp6xJZ7tMmM70XKx0O8Ygk7hC1ER0qr+ZY0H2Z87v3cRqV7
qvGqLkxbOAWab5oLHmlykBVXE0l55E3r6gXx2l/Y+H1aDhI+dvcVjZbd8BjNA4IMPbJP9b1pZuPA
AuNOo8RCCM8Di+D8rEzUY13zchjMbtgY5efJmKJeV0ovfdw1Zg+OKsE97u1WSjZqkQ11i65dhUoA
fqDsnQhAwVeqgHf3L6Zz7tQrUUs9/KKM9aQ0wdOVICNLygtGQ/w6Ju7HHBPlDBIhmY0/EOsCxbEQ
/tvhHfuopDGVu1urCWduvVFV19sIMRQHnl4RVf1kfrlzm2BhAi8qbQ/6Ay8Zq2lSEKOgpSFV+0P9
73w/QXBDtj45fFQjrdY3XqDJ6Vr1u/OFJVQRarSAiFDKdqWYy0whzBTZf5cjytBt9VIbDCintohk
5AtBKmcBK7mSqstJ9et7X0vB+mrHnjas9B0K10V3GIWpWVIoY0J3HCtaOHhPPfGW+i+LLSx14GMm
2rzWQyFuS4NbCipCh0/xaZ1FGr91ZmcF2/ikB9HLF3rkCK2zJqzLZHoEaWIYHcF6G8eYlqEiN1kI
gDBGqSQ6tU1ZZKIZerwcOLY1h8/J8YmxZVYBqSoMriDEBya7lS5iPI7OTi9X/szx16KWPY+bHnB7
YDjgJbgGqJzWJIlf/uJ998xIR8z7zvjv0C+7r4aUnbsZc1+Y3VM/NlD6+KNFFbr1mO1E7pjdlYEP
n9BcqD222dsEr5bEXD73Ny5kjEN07gOpB9S+lDF5gRWPm7V9pWJsjeq6WupAgNC+yqqSKkJbUOYS
/iYws17xpoiAW/8OD39vT1fSdQoyY0ed3jmtQtEM4++WnSInpSbvbFu/wxz3gTFv1lmC8wTZbDlD
h1ZKkF7upl8YlWsitEyz174qnLWnaBslkF6WtjIjCNkr/YLPm6KxmnrrP09pk4ejLwPqZQ0ICFWs
rtPYe2kHeGiXP+OV5sdIG47tXo9KuvWnEH+T6XMtt5ZlzU1bg9sW7PF69XfMJ3HhB34EI3qwCIVS
lw3uQC8N++zTjUt3dAARCcgoN/scmk9+kKxtE7HtA6MqHg5TmIW5fpF6AEdyOLsAPwkQAu1NkFDY
mU3Degd3vyO6MnlIZ2FEQQfBnOOZ6Fsi5GhEuAnjbiVWWGBo3Yoox0FnknekNRib43fwcaferTaG
r9t3vd/2QXniPaFTb8lwtSmx223KSucm0xccMdtLqI7CrceAYIh0ukFttzmRlw+bNRrm+e/GER+Z
eTA2yI24Vn91vpqHG4Q/zYds8qq/UL/ghi1j8Rn7nYf2wvfLugxGvobN5gjeQg4LyIG7Mf5z20s7
KJfeemOC1O0lK5VyqObQf/Q9ynW6mzjEoXxXjBE1qjdVpsly3PIV7M0M6sUP7vKNECzo2TAw5QMW
eWCedhvuwcg1JBYK4tJthzISo9a8rlc1xVWxDyvng1NkkR5yzUqQr9Y46B2DtdLyUomRdPrbrGP/
buV1DuUs46L6SZwV8ou01tKyc1K5F0fbiVfE3RhEs7yGcAzB+cfKoLZhdhiTw3v1cDy/xU1rsiNw
f30EkMVmtiSs3/SEwEyYC7hz/sW9vwhU1rtahJkHqOivKXoJN9EPesRnQ5lR1eNjgICSf17Ugekc
gpphzSSt9mhS1eItQ+I2zIgwFlv4GUJoluxJkjUYuY2vD8Nv5yKp61QnVOv1c8e43q/kaRNaeN2W
X7NzoMoNl9P1Tc/ioBkpJWR9oSTss1PS8w55VLgcZD6y+SzsbxUGfx0+lXF4+f9N5G7PZj+t3ka2
ohfCbEYHhM5DkyMjSb2taFUvXreHHYfBul2JqAIvEgpF/r/jodTDtyoJga3pWrY/1PG/RNEdimwq
28Z4zXN+BeY6OG01v5gG/wtkWOVDrxO0jaRord25XxFPvaysO/vuWSuTsBJkdQIgdaIl1BgFsJzX
6UH7E4fvyIEXPTmAygc49pZd7Dq7QMRbPHDBXfSES1AVoSRXExSirk+A1muIBHjNRpb4XaEPKm1B
eRYqdeEmMwiJPCjaD9PsBv9tYY9UHzJWAIPxeIdyXFnUVfoXHM3vPhIvEomuBTEeoh58O1XRoSNe
qS94uhN5dFz3flseKURk2H+IMwuyklkmmCuY3sYJAIPgJi0MlfTnVMyJd3SoVwtVJj/SVnyMe4Lj
EtyMOtqX2Hdc7lzSNjgJVsJCTYm5Xf8bSz79E/47095XayxHnxfqW7/pqfVVZfah7YsFW4wzsZ8M
gQoVBnMYSZ8m8FbdVYvA9B7B04LMNBHlLt52p3wgbPE5Y+jk7hRMWC/9AhCVSjJcDnViwXfZHo+Z
G/YiWrgPm4zeriQxXpoXNQGjXaBb24VsVoLPN1NlsDL+3CY5HUZRQFv4nRjwL3Hm4+hMYkZyYwA1
2tDNslkiZmG7dxtYXIjWQn/HCmo4rH9a/s3fwJc3TPGr2a7zczttixavlru5Z5iugfm6o8kUufUu
9kUxet4zYjmFWvlW1nKM8H7hMVRSplz4Aji3TECbTffPpiIaPIAynKx9+cr0p14LKdxpjVjLgBB2
rC9wDxnjeYyKBCw7ZZBcBgog0ScP1N6R0iS5GeR3mWijOR8XH203Y/oAIXFMJphDrv6CaDxFbE98
iN/BMgBVYnoGGRYeG5BtPQiPzHMrveUCG+Y494O/vr6Ji2cY+sHCLZz87uIZjx2VNTHG2d3aKRz+
iJxnE2z5NLK82YN/0RVe9bnGq4rXHbn8h7GbfZRplDaSnUB6vRJsBuKA86z9WaNyzUD2mcHCX+HL
lXiTSkyFOaZi66IxwAfReKPnwjjoRKCiS/90ewyZTdm0QepkXRjTZzhrh15WdYAp5S+nk0L63ve3
PEAKtXgsyyBlhHEBfbqX5eFX4txzD/XZ3FJ1AhcZUF1eODWXyuZNhmcvxgYfe3zJqRzJMUa8gf4b
cSE3avwi+7Ydzy+6/mjuyd/Ko9cMrGPeMsgfHFmOKLSzkfvXbWs9Sv6XyPSFIM9qE63cYlaXkjlp
2PTeD3B+LA2dUkCuYfZ/TE+1xoTP11ROsSPZasX7L+eLVb5oH9qNtcZtArRTXLXXZ1YolggHA9g+
Osy/sFGtfNqd0c5sszr0r+UAF5cVL4qNBRf4GYoyM1CbMgclDYrzNoYSB6R/Uwx9Jw6Hfw4jbHcm
Tt9lPGAJ8oOcuWycYVOg4G5NGln0jklrHhCMNaoJ36h2OcPb8o6VjXfpamfTESfNzu+Spf/ZqB3R
FwY4koNvH9EPdnutgZQPZYiWICfaf0qYmILWv9b3QXNVUK8pvTaAwjKkP44oxrFIlYL9gkOdez8s
v3jpY9uZAVr2c+m0mDHTPhR1LaR2gYJptSVYUNo7QlFYPi5bEbvaRi5vbi0vCn5j5mhpAVy+ck9n
Ct8uuCqTyHqgffW4Hdcb8thta2cyBQHUFO1eEfY+AHhemQfYScO2EpStcCGqNUf41gLwLaiUzdDE
YSR/WjqTp3KbFQ4uLBEN0hf7Us/zs1OQS8D26r0rhkCT8ST6fTRzNEdeFk2yfG/lv3BQsyMoshoL
M4Ky0dsrW+eHxFyQ0yuYLtbzKpY4uLXqJRgCNqVU/rZ5zMfcmv7URgdliLus9824tdU2pRQhsiYe
Tuntpfpttd9zEhmw7xgjsmGaldsdzgYl3Y1/mQeuy3nNbdzSETuciZ1fEGRxpXPhhQqpnM/XmpGE
wyqd83x4tUBacwQo7QWiSstbbHGDIiz0jXsnAczw1//C5L+gsedi6ZLpx7c89KFsEKG5kMF2eMYx
q4eHgb1gkVO99i5A3o8kn6/g/CrguvUh9sH+WcpqGYJ4dux0ts9yraj+AMukks9zlLuWMBX6rLT7
KzxJJA75FMGf4NAn1uyhgf/CZMmUrZrYb2y1iWKcN98HwqypevTwAbmdG0CVbc2RJCW+M2MtIdTj
aOrXZeKv1Bt6OD1MJbNBrAd8h7mbgjgnLFmBLAp/A/noHMa+0cVXcApXTaU7hbjzypJl0ji0cCoH
bk9k//HGE/Uxta+nvj/nnlusFoQozgjHp/Un12xneLqmKLk2eBwsBLAtV439fkC7N/D5hG9DNjQu
zegfsfTGzhF9tdGfyNSyDhDWZWYJsmLunoQB5DRc/2/H2kSl911FMJSwou73xdZxAwnPnCD7G6gt
uCrlR1dPaQrz9kzrwaz6G8y6B2Bzih0Cp0lCr1AFaQHkAWZpzAowjP+ZYf6NUZZ7xID6ThB0kSVD
gCdHpnDWLJx+wlS303dQ4GHTVTGUQxpJ84Xy9wi7rj5eWWM2VEqDVjOPf/CEeNn1IE/57c+Q3EMR
x2oyDF1M+76wrl33KURogShz6QVvYbk4F4xxqg0hWs1DA99Fnt4y4HX1v8LGPceXnt6cJCw+vmNO
sHV3MPUaecR2KabsG0Rfp9cEargg+k8sUZm1mL574fkKV9dBGqk6fqHFOoS6PDtKekBd8BEOk3m8
UyMTbk5JhVawh3NDml6FJskp6wgsRVnDfXpgPXmiXHVPQwuji8Ow1VXRx9oMpS3obI0a0pW+NXCV
9YHbomQ4OJ5q5KRymmlVxl3aIkXgkHbqEmvO7ENjs9IWiiV5xszYIRtzC//WKxxOFSigYC+EUjix
ZxjoCoeyOBqM3rcWTVtOQ5EUD1371J+zwcg/S8f/2wqMzTTxz1xmpvZj+eVI7lw/Yuig36y8jwFc
+l7dg6uZKkopUPe68vTMrmF5RwDfVXu1+bxNhKu+/guH2WBU5uX8nkri2QOrEe/V2G1xEHol1W0C
3tIQHUI6XN+WlpcFNv9er15sro8DmN7cQW3FsFSkURTLHwmIeXevcApWFOXwO8peR9PtNLG1JvbK
Tp7DNfEdJtNipaDiWjPo3GpHmkTtdCa6D5Valx/AMz78ZWaWbOAElgN3rEbtvPCfKz6sxmHB6v+R
N57Vz0M1PrxOKzjOhKofFL2RiRYwTEgo+JH6WPHGf4J/c+GBe1wm32Fp5IG4hukJIp8tjeInNvBP
hrN48pflBMWWH+Pyft2LpBluk6W+zkQLuHt3d8bxHm2nQVaDerjYO0KQQ5JxIHv2SqL9O+z9ZoI3
rniTR3tsv2l2H+whtewgQy6OdvjGjHCUjcQJGyf75siPuxZC/vXmJtbW46tF4oMult2o6EP+y2cf
vZru7N2U0sA3LlvfyG5fOq8u6fBg+xfUAB3zMQgCaUxGd1Xfg22gZYOF6XmRpbx0vWLVrhgDsdzG
vIcJBDuNELqhqJIjUPPRTCCLc3JDnNnni4tuhXAAzk5rPkkXXY+LlMb1pwEq/p8S5v/3P/9zCPLJ
80vX+RblYjeBf6/JhG/1m+H0Xe3TnWFwUT9GFrJyz8RRCE5h3s3gYId1K4/hA6H1Q5atw79h3z9e
ubS+/hXAHy9r59ljA06PmynUu9PWkWWt38ZL8NdwKDHNx+sxdw/mgf8rJNT6hjx4jIN7j7rXFUQY
qJMOAvHx0jTWvIOB+KL/8cFR3UQ5KdDBrQXo0MBS4s+cv4ijUtM8f7sgr3Bs4zlVh2Ej8CxSQV/R
8EHdBrpyE1T2EuRa4hHYgAyb3ruJ/gZ8YgSv2Z0+HqIoX3IGIdXzCT1I8J06wFKhAP7UGeIWNuje
o9mI3Kn4WKXUyPNqyhpWXe49cSnRe5jMJyCb9xnWyv0rJg6LtLrcw1B3uDF6bgp7hId6CAjzfGP9
xMBRS1JXWjmS7YW+zHER8YV14i4+rnzG8dnT1xJQG0hs8eTfC881QPjW2Lstr3g0xPiu30hGMe3b
9w0Pb0cz339ecOEL8jMAr0jCjKhbe//KtuiGNGiBEaf9oa/wHvDOiKTPxZOQ+q5QSYSvDqiWKpmz
k5x9YHksrJtjiK1uX0CArVH5MJTTcNAf7JWA1OUdBDi3gBvFbhG8OknO7L0KU+WPAhQzC7xFo9hR
FbcBRMYG2y1R/VAhg5htWWyBB0Hfffcue/e9TrJDqbIqEimafuhqDsn0e8dkpTkDXx5alvJFCYzq
kQDoO/LKCwLjrrLPlGnBFkmSaWBx2q03UHkAv8TPEHyajayAV1MGIchOEDRowKelHvH87bJ40Ba0
a7zd9cBK8ypDYI3g3C3R+rRh1KOmJZgeVBUai8hwjx75JboOQwYgWLYwCNpVpHo71Lg0imMFPtOp
Gsv+W4nVF0U8Onx+BZyrzG1TIBL+bNAthl8lE+9gooenJ/XxUQVh8VZBiiQh3i5aVVyQAEujoTOv
jKkdCW9pnTsWsCdgeXhzLJCP0Ky5fkid9YSKH3Mzc8jJU+69/0mmRPCVwQPrFn44AfoiBqDEsCcu
Z+1q5+W6YPkOum1U8IjmJALa7tfZYm9iLZrD4O9nSpT6ds2BhmhXDDNyyemWg6tv+Wcp5yI7W79p
O/MWRdWlyCzrPrxzPYTagEZ0qLeQryZkVeCZtRy2s0Qb9AiqF3t5PymG7h+aNrKAur58vOqMSYGY
4kCaw0FudtHU/bnttt8wGZB3fVWLaI22mXtQPakSkerufNrp4nm67H1MqCgzNOdDBWhJM8Ci/EMm
Vj7KUuViRdlW22rnf8xrQeTatU4fbWMX/TigPn3dADKTFcUJXDp1mWq5c7GVc1nkAus78IpF99mx
SnndcHLSV3TKf/WESSJTr7vPkwvXr9KSudJA5WxeVKI0YOurMzZEdN+232WaDYf5b/8oPL1Sq36l
onajOb3fo0jSfBq4mpVF65XxCvxIfwwGPfQTfOjyKDvPgSJrNt4/5gBMdLYaqVnqsuXQkS6wbPTg
8NIzpdMi/nA1XuZAKC2UdfYbMWxW2wp4uz8VVgcUIEwcza0RByOu9ckNXFIDmw3nwAc1kZGEzxDX
OXnQNX54Nib0zCbijLjvka+du5iwOItpYwBfgMixvsQwOtjWcdbvm+xFUTp9308bbeUUWWv3EN6M
9AA37B4BL2BTZshZkqxoGigl8kFlwKfO/0gqHKnYmyc9jSukHsi5DEeGqAd3Mtr8YToqdXw8I5UP
0NpUBMcBzt/eMRvEGGnZ7YCBfVU1V08r20v2ZxwnIwwbV51AWybEeJBCbthdNzayU6HaZAiHSjE0
+5yxGlZYa3OvnPAF+2edhQD5hFbrcuOUbSIfZM9D0grWcHfkmNNJxzz/N7RlvMSGqVEecwcbVxiR
2rtkKKay8by56eayNW9vV+rXf4YfRPcqecx9VIKjTiWOAbe4J7BRMVBDeTBGnljkI/Sj1qAZpwVo
HzByUbpqF3zu+zrcWueFRbgLSNm+KDwhrlYb+6wotDUJ9s2YwI9wQHxX26VmPKkOqtdo0d7NvHv8
WYv7S1YMOKDMNfjQYJcGyC2S3jPcIoxcOgU24nd1DUy+uarrDIwFAPsffSeEdzuBq8wM2w7JIu8C
rKTE1++2p8kXT1+tqgTbto7zKoGaA6f1S1jWlxx3lFo4bpu50BN53AruITYfxi8gwznK+RoxYRcH
ZyjUXQu+w914RDd3XkIoTqSrIvX3X16i7reBiLrq/U8WtufT6VDukFiXV6tOOoLPCqlTHBiIohUh
OhFsBBVoHvO8rlsX9CcFeuLxECz6kggYc4r6dCis/mHI+fzxeoMmGM8PaSJfdzyFstijp/VNsrli
sEstuZorCh0bLKHDpfL3p0tiAuGIcx82SltEBb/vAysuGKn52LHyValU0ce3KPBq5uOM1VDz2/pE
mcBaMV1qQCqvLkCGYGbEcQhUY575cnwMBTGV8NcE18h5ZjbjGVnrIDQJE8JK83Ud+bgHUdBasU+j
/qSaa6VZF76elAu1XY9xwjGtv0lKDGzXyrPZpVYr94HG4sBFWVIg7syJIM0CuErT7+cMLRn8S30t
Kp73MLbe1gFE+SjeXhANtGRKA4MuBixrDlnKraBHtNUVleD+6CPCjLyDGkfdf5/jpE2075rhEZnh
2lg5/L3EJXPfcJJ43K6wOHHVzakVoQUJoemvlY8OQXrzDRaTwCgc63Ea0VhinsIAFe+aUTSV8x4R
ejF9+hZ9GHR6ODnb3Wf5FQVhK2pX1/U1pno+oW7JKUy0XS6Yuq3flOs2WLp2UCrkC+tsp4PZJCdd
q56JouPwog45AZxsJXTgSROPD550FWkPZJ4yyPA+gQVx9SHm+ZLK0E3S4gm/ofuUY2RIR330QigF
nRUIOtCOiRI/r1Tw00Cm+lvuUXiYpg8gkXVOFy9SmKVpe+q4d/uuN5y9JkFGBNhgnmwV8oPY9qqa
aCBD05RX2SaUMqDzUkGm1ji7/uC/z87w3N2AHgdJRFr7LWiOaaJJu+L3oD178Pb+JOH76GtYSTo9
1i2enVithtyUoBIYRl0JNT5OWV+ghBUFIVI0IZ9O0HaTsij2/+fcFuJfo/T4WeTjILMeQcu8Q83A
Z51QHGN5U95ImPAt+XkzS8BmAy/l2/bDKcVQeuY+UXIT0XofthxahTXdL0ctQBXHzSA7yqNyKvdq
+wH+8ljPljccIMtpA0EegmgnSA2iXw9T4QOVe2QJIKcgQXD0qDG54LtWALkxo1Ms7mUHH3cUHZW9
RfFXEbNGPA8B2Odd4xk15N7mV+h3k5a2yTslYhi76MxaY89fJtZ+TbKq2Gp4z2abEGwTPmqG3J6z
hBNx4RrmnBqznULgp+4NxR62/iHMFLlrW3NRIs1AvTwyg7eSBob+s9z6givVXap3mnN4t6x5kMNg
kgIoZtH4rK8OFnVQvyWFXQXHsxjU+tm6r2SqU5DJoPP/k0oPWz3PlfMeCszHIKUyoXFxTn6Kebmo
vF8Gw2Zk6LBvjQckQ8Arnnc/ZdRVRKAWC+C/ijLh4pfmq91d0aQH/4cY0AAU2W6eGnriIY83TjBE
B+pq1p6H7DcTbTfdxbzjeyTRuIMkZbk0ibbO4+n88ZJOGLrDUS9KRvXSeD7E1ECwykj4rkplMwM1
X4i4Eesn3vs9jEeuCuZl68fjkEJ5TsNRBmsetp6NnXanm1HwtUSHFet7nK6Igl+7ja2kWZwyj50F
3iG8BQ7+78jkdSMx/u13uKDejnOHT92/4YwHLdaPJcxPMBsDwo8G7FYOyMAzsLvvtG6KkcXh8O+C
qf//CTtKiQ2aqjDamkacNi4KZtsphFE0zV2Twc8DWWocJ7ECmuNoCOPG20jFxahSNdz+7RMDWBui
chCsI9BnOCP+znE0qYFMgA29e/ox0TQfuf2tSlGZE2Ftpx0D37qR3YPWY5ULBLO77D4Rwhd7pfJh
o53AjPhwn3FIoe5UFRttcfPU9GFwkvON626XszfCxwoZRrWTBZhGKh4OAhD6w4Z92so3eDo3jEZj
8Vxzecqe3ePNyU3VqTHW2NPwfY7yWgJ31V4yPGDNO9R+T/cyPT8ky1/EdwK1DjY1CLtvVjQ+r6SN
gPR9mUPfoRexeQ2su4czTYsiti4L0FrFisHl9t5fXuGfdyLdNgrWje0j2+armRKHykADYkKLNSYt
MJB0oy35b6nBRxJv3OOK3XLOvaD4Ruklh6CjqkBIdybQb27xPtwmAENxfzSh74BiJRiXikvMDgJX
vp+KWT1CwBW6RiWdlIMJ6aEirjQFoRysUksZ+JRDvaKgUUiL+ZTL0gngU08t+xN/jkDPR9w2m9Pr
Bmjvoz4RG6LVm8cGcf0qf5S7mWPvlCQftqJEIGLsUfClzBspPOQy+HIt0LAny+QAhtmIoK7eAEjl
MXzEggkFOSN51qn5KAi3a6DDk82jiG4bHRK6FEm6cNhc8bsf8qwj5TlJeC6hqANdIBVwZEmqtKYW
dtirx7R+1aXr0JnC8MLUPTnpwlQ9Jcn4sp0h94mAMjSx0w2naQOk0oMr03xQhZlzdzAYtoTFc7u1
wbLQp6WSTdMNpXl267Ny9aE3PnwOfXE5giX1yiiTiCOa55YKORk5cgeX03A6n2+H/6oDLyKVPMVl
l6O7DaSSs5O43iiWVMaq2FF1Z+ZAuC8dzV7/fjiQ/rZD0yarbWR3CeOaTYaay2fwPja8sn1gyKyw
HYWZNeDXkLrepXx/Kb94rp75OpcQqrGoaO9hRZ5raCiGp7q0hj0BYHai7+cYpAZsoGClcg7JgDwq
9HoDwO5y3rtZXIiGDFCbYaDLMz5nrVfbE/2yX99zv6hO0W5JeW+Aduw/AYQDLEBtNOKvAttq6XRO
84jxTZqy8GW51HE8EDABqOP3M8xgJm+RS8DvSwtfAXgsiBd+XARmfvHYkKog8euCDJ/UMrZp6+9L
NxEBu1YdwTPIPeRpuMgRadSA6u8AGdXGUDK97goRTxFMJfrhEo1vE5rTxJJBUkkTJujp9nZyf9xb
TuYA7AZqD11s0ovw0KOIjhUF67MAovGP5p7b/QUkX17ecB8NIt3SVjux1CYUOTZAFNZx94oaz8/7
s5hqDsWvk+Bu4pP8g1hjrnfuIFKuJD+Xiier4beChSWCKgsKTiyQC5ye/+YcfK+5twZ9ZMkUA8Cs
HGhMhoeaPwzPhneMPt5n314qiGAK/H2TPpRZC/Q/mmKoMMcUNFOQLxq2t4Qym9Wgt6T/0uYeHtAp
VZIoq9MPwBX4kfrvgwrOT7cs+foeg7HV7wP/MggRAwaRGOx0aLFhOjOFl4LjJVu2ETosQHaW7g4U
eye+kXEOABrIU5/3YKcEqLWnbKVp81VtPE1q7HHcqz00TPyM+SjHYG9xQljlPYkvd6/AkQA7c9uL
lUzMYCn4b7MkVmYhwd6jjW9qFJ7/fyTU8HoVomeqzgjreRO8EBy0Asb5tOvxWa6dAa3kPZEwFgqf
JS1qTqSmKmEfZoPViGKM4J+Hlx5XBKtZHmUJ11C+BQ0TH3j4XttsP+5OloLuULSf+qYFCUf1W/jp
a6aqTy5xq6s7wTS08j8Y3wP7W1kmfMYvQ4upNg/QytPV1HN0bkXHJxq0tq2BKv17xWIRe3Ep4WNS
E9Istcv2EOVIzwtWg/5Tal3Mr20/DyskoZ1zhVjN5ia2voNZ/8jr+WNSgQTZ7xTM8N5+2g01Tv4i
R9xr9maeorcj1bHLdj+r6ds/uJlfY0AREKH/p11GZ8HndSxfqn7fGy28r4QH5tu+bkt4XpcffrJb
XqyrG3M3krnPP1RffkMWAWROCV9BANn9UaVM0yS0K/DTLkcCFadOQBGcNk3acHNQm5ruUcmc9t8v
BUN6oAIt7GtCQGSAom7Hjaq1woaV0fKACT+AgilrfY6YMwcA+E5v8/yPqPZQGM57YJ6N7Tm5Pqry
bqn+i17BdvAvIRYtClmyKtNslC5R2G1tabmv1sXovtQoPoqd6QVJhs8KDOdDedt5SQ5fE5goOj9x
6GaV65FBXgFAqFnpy5+VoYG6RbnKFUPHca+Bafv5IrFSCPlc8bfDvX5IvQRdUNCa0mlC/GgNpsDx
wufa+C7b86THtypeJ9QZHAFxOB6qGhu/GfR+vikGk5JugCNNhP7Ew9aTxfY3FiVPWFLlCgdqqZXc
2GbF6ou5g0FvOr87GFVDtcnNTTU24Ha/RN+Ey03P5lLmyFJQZycL6WaM0mOibx742BTIQNVx6ins
KZhFZO9X/PsrtuYGRNNCl9jPiXpe3E7PcB1f2wH08kGyx/077PdOIiKGMamRzu6WPI7T0VePyZb0
HOQ12LEhx7wEIlvabZJ3VClqp844njW58o2nn0/sAiyB3S9jhJdk2o8gA9hzDb0o0t3H8nRTeTjc
CQvd7BMxz8tKndsYhcLPiEhlI+dAzQd+0NNPd1AEY6Hw2eaCjjpxtDUAcxZN5rLd+Xp1OyEU0rCh
w2lFDwSAb9k9ZUIEiONAbl9Y3DAv7mnLZEV9zkUpRjZA8oqkWlm3ezedZbeVvYmSujgJ7pMTCijk
bv4Fj1m9wE/pZwoSNY8hyuZoL3yykXCKoFee+hZ1jLXILpr2DcosGSMAeOfZMvGxZpY+BVnozB0/
iO+84nTBKXrpBeQf4rENs+R+ybnFKFvr7xy9xIrptmmWTB2kbqUe1q/Rxdcg8NIukfkE9M1CuBMm
sI10Z1oK/nXvtAusD6QPV8X7oiy3pFeuzkSC/HK4G6wfgPWCvxeVFx3zfexYiCZfWGjMofIl8WmU
5uOn09wW76ynF9W4BkdpomWVCxVyN5OATyTObGcc1FkbzG9ddiusXnHhqdUQzL9R5PJxlTs91vFu
TDd3x7FF4fFD0OJWedsnkvAs/HWZGJhFkHfe4sMpSVrL3/hcildQ/96bENIm5/Mq5edwsYtYMPio
CjIe5IJnLohd/wn3OYCMu6ixlBYTsGj7+3NQ9WFy04lQ67QPLH9Za0yt6pTD933BdgTXJaZ4/42/
hhAEDRrPOn92cgIQJM8bbzAFtMkvzFpRokwgm1Tc4vpUn6Nqq8BGm24+TcxoxuPfrn4iYA/4ck0H
vJ03N7JaPy1S3BTjY4+8DBaEJ2kYRib/+JNhWgES76j5zura/easCPezQtki2EY6HSUBIdn+ab5+
/5Jo3W+Oreg+VyIXr8tHReMPVvVrytS8FoVsBRXMnhRMtx5nuMc47qARwSurTM9r1RxM2R2pU+OA
U3SXKo5WdEPTRm4asJHUBH3Gyq2hzTUtvJukHfauHN+t1KkAOtCVFsSa7dwGF4GKg+m8qNtYmt9O
nOYWOCef1K1+Fg0ozlT//bUbD0b5CPPmBL2Xi6WO9iMMyExp66UKycno1JnvEaEAJL+D9m6QwI5h
C0q2xS/GPaf7311Z3iEkZrWLlaLAuQzH9NHMUBUY1s3ktH7XjjVyLLzkt0wENi/iD9pn/ARzxDJq
OTDRyVav712Iyi2GYC8Q4XDUv3A24MpG2WgiOhEOKDI3v8L95qdCRbRvpWbegJSFbZADQto1drbe
tyA8jQ+LgEo9tLP/iDAcSZ/XIoGQQbHcxzRVMFASPKSPMM2YdWLGzrQDyiN6q5XAlq/eCEYvqYMI
a07X8SVwDAFkjhfV+8id5VjBBacA6wtcWV3MbM9XdRMLyKWm9lG2Nr3SnPenbemKMWj+7dv5L5Pa
tlJi5TqweukRuRKapxcmUK2JkUwREM//4zTGRpqVTX8bDTofA5zcVpRxeDOKG/uGD0vxZzyea5tf
NyYzT0F2p4BVgSjShadeKbxTDiigV5cn7r1aMfo48HBc2UcyUjYJd759n8+V9eTfda2Gq4Uzf/9A
YcX4T6JG/gdJDFFfTtWTVvYHXHNeMywY7XX2KYEJCbvuHBbjDclRKtjw6B7S+a8liooaoaAs0HSJ
JNwZv1XtzW/MhXPxpdwf+2S/V+4vjFOZapY3wCIbZaX187HMtfX6AzqKBrQ5VftyWrf2c3R4dOyQ
n0gSmfRJA0/m8i+qQjIiJd6WeV8ZLHLC52PqrhFhT9zsUYHhjOM/vBv5lXspixbK2AXjQlCaU642
ZtSNm5IuhoQow5L9hv4bDDEkWncltSRE4lXbL31EzCg1H7pPbxW2rNAj00nEUWzB+ZUC37zJpczL
oXNobR2OS8KsHPEKuyS7lgVkQmA/esphgJBFVFvK0bVJpvHAO4SHliYQq6KinpITCFBb0A1tkqjn
1ks1u/DQYPzkkj9ixDUBqOzixQMIOcXIG/B5znzkqEOM0hPS6yYJ5UGqf7BqdPc3423JoGyNLVxE
svkHWLXfFbES8FOuNVVAdl+wtxUdlKDTpSHdcWqjXOcKadbPuOxdY/dFGjKxC+kJ4n18Q+IB7MN3
29MePlTg82wDGe/q3i8VxodukkvTBdcJw/hhlY/5YRasNPyil1dojYC3RbuMUFoehuwrnZrfLlDx
pzMv3LKCCDfpPRPH3JvJXB9qaquHSS3EgU7VL9CSgpPlazto1CTdTFrsZx3uddidOhcaNs/nRjOl
R7npMlmUGinf4n4PFhV9k9QgyYmPAG68tG0/ThiPYZFNBgxjSKyHyfMKBjC91NJxcLfCNCoAP0QE
hvHWvfeJco0jhNS3J8L9QAwQyO3EQlaupaz3Gi6csFIkZOMjBSbyGKkmdpZ6+2MCJqkFmwTf51o4
zw7N3qXhCejQN69o3nVVfIfW17lQ3HTy/ztyNjNpGDRP4+0kQ8+i+lXXUsCS31wT2nHmC0qpZRuU
JBKty0pLCR38GaGnwW9NcHmcNnOeA2Nev4S8qOzoNrrrkIXmJcKgubWdT6jtBgThIxZtfLmeJ6Ai
CKXN1MpwsvIFRYapPlQm4rMFvIoZ1TYFCFWbvxNnEQr9IMx/dYvE1Yk84K/bKZJ3GHEWF4+cJSRa
ErRwQBlT3ab1uLA1WtCHZt/mKwq03Wx1zIUut+DxJs6I8WUNVOR7WBB5BvYPlPYo8vD6d8qSZZkd
as8oFf0cEeO6x9/WoMNVX2SMKE2gHL80OWmjK2r/BC44sKTDBJblCzhZCNwbfpzFJKUFgTYpXqg7
Rlv08DQa+X9cZb9slpwe3G6Gdd5AYh89JDf26oxxXZh2HTxQxY2KLO8GVDJXtiOyDnoL6r60rXgM
asDnfKwp39xPyLCtKyOvRxDy2xM84qKNNZ+koHCAhe9pJK6hiwKeisPeB/EdySy+5D/6mUvQQgtW
iGR1jnuApVCOsbeXL2IAUGhSNtVgvVwduebFNPHN2igTtfsSvoimyud38eE7IfnQ5MWA7fdsquM4
ncO1OGURyS6iJKM9C1QuqAQbem5bUarspRPx12wcv9qsC5J/PYeo3MbrPBJuCEQNUV0ktCKWi52C
ggQ2MUAHx/z0zj6EBmsLBBGJcnQOO8KGumdDhy8bfQtIkkJ5XzjP0NSGhL8aOlnMCsYEvnXkgT+O
KatnxU0fUgmhmmaOFMZtgc99kgGlGjZ+IqmI9bVTlcJTgwaKrWjA6chBvFq/bnTJEKRRRQNpvImp
0bNJt3uxQoYgXAZQxUhe7QOpqbVgiBWj17ypEh6UY0CJQt3DxUOnuBagSnrHwzPoJ8c/5fBe04ck
Gosw1sLHsjqC7U3Ko9AGJW04Kx0l8X7ndROUXyqGaKdOfCzlNDQTVEUMilC5xTFjcjYOefOsDdwe
Jr8NRiSqZc6dzc+tXPOzQg8BcAsE4M9WaZIxTuvZYUUYUZwp1YGfJw9CA3oXWJCCagSOnIbwNtwQ
Re6+31thx9/iuPmW7ZgRY/NcOqZNaeuC3xTwJt52xZyeaoUVWYYPy+OCjEXZ4jJnGpNy9sdK/cKU
bbuCgN5WnoxmqXdgrg0Wd4hVve2kvd+kU2IR8HiJHjt9rX4CqJnk5kfvGamvM+nAmshV54DrKlQ8
7WpouIPWWndcL5yomfon0b7Ec+ETT9VH0wI0NC7rJCCkh39EMg78sl03O443Tz7Hkcze5vh9KBDO
dnjzRlXpHOxZrAA6CfFBilZjEtHP5dPYONSaecQ6g/nNGyLYSHvaRIXAeJD5/qVtCDsHF7A9nR0K
Drf3p0gLulgfW+t+8K+FRZJyQvFQVJxIua+9El9QLrh97cFLX5fl+4cwiw/BJERWJRdfhB5ZTOdS
gtSPWftCHEqbS3zIt1IzFJnDJnWu82uKX0CRpLj3svnS8EqsLN386zRqQI66b0jbEli7Lscf9X+h
OCA6HGpiDed0DkNCbA1xkPZslTtBUooe82JJhp/vs+XN1nWbUi8WK9uZI4NzZ9Dq2RM4DjufzZNs
mxtjdCDhA4KhJomj4T1Qg3tyYDQbKvmF9jAGB/BYga2jiFAdpkOc+Ns8IPHIz6HQHOcrztFyvRCi
FhioXj9/4rWOGXRllkX48WLrjaQCmkbWvJW67llDyaQWGed7eaHHf7xcoOEjdcf79wAZLeWiL3yx
S/CAGERqo7v/2mkp1xt+n1r6mIXKyJtsunUET0JVcMdhjBCeeHnXCfyH4xakiBVanKsHJJ790Sr0
zW9Rsw6k9UTZR2QX+FUqWOkrUlmhDyf1iugSlfz448SWzbX1Mxuu0ZLWh6kfwWE7dnex20vsVtmg
KHnRDDWn9MORGembJL1dkULuj2W/b559MpG3TNKUBKtSVp9Ooy1stRW4YgSb/bkQfExppckO7I4J
r0oTHoogBtL5VZsm9JYWwmZXfnLPKHbis9ddC9NQyPmGDCZm5MIGk6ihTbfazH+aPHwO80kINtt4
jxu9EYUX9qT8q4k4wX/SXBCDR6Z8XLs+/rEI4JfePnh6yaq8nB9nkA4ntxXzcCNhuD1+L/jBbtCd
pmBKbqW7OK/RYzDpvp9q2JX9rhbKVHZ5Gb8sgA3Dujo3jGzBC3rCUvJz8bL3pH7s1XaZ9OghUoHs
WS4JxI5nQCOJbVLLMjjSKXON7cJO1Pc3GjF6RFk8mR+XgBlqSaTBvqB423ZiTF8wrSynPX7NSIH3
gc7BHJKrGpwYdKbcXmObQU4A8bXExMiu2yu/Mfd8YeUoMNXUH/zAaKeXm4ujY1vCk5ICDBuFfHaw
bkI1QBj1cBOkcT7KG1N7ZqvlsiXI4MNXzFVk44PebVdgfZjnmtGeBJqvDa++in6kYdL8tdLOBQVN
Zs4CQZqNLUzCepbq7OxQxEdFzDQB5HnLAHOyUihpGBAmRFTA/bus+/CJOojJBVEU3nDS8DYz1JAv
SooWtNmkFs5Nl1xUCAn9EIA04T7SilTsCaKcck0/7wujIvv9oac60Zq0MpV7Y0KfSJ0QUSu0+uug
385byHAy/P3dgq6u8DqP5gSmKePz7vcOiZHGLQADC0D/cEdDtkpA8kWfI3GmZQkXev/Mht4eETcr
waOiL6WhZUOwKzFVp5K8pvgs9gtHxF+pyiKEQzGKu8tuev3VjhMg08syrLyZ4DiMrjqxyFFUgh9+
Njn9E+qMnVsba8GT+IoFrXDdFfmhVXwO7zxEAcFgu0C+bTUOoI7L0LQallUJ81+L15CC227It+b9
sbLa9H9akdIa/Fi0WrR5P0dxROUP/Ew9RzV9JFp1suhadprm1pwezq1zXCdtP2GFTBObjyxDr/yO
vDkvfPHvUu4vlHg/UgKvNAfKdaOjk/OuqfT0yL3/yTKX1OdMtKW/wXPRyV7LArjpl8wA0FML1Es5
YqGY5H2gWJ3wiefkcwdpRZjPJcPjstPcFcaijlU/kgqd1ri9G6S1CR/gUaqEv6Y2oEXxe/0F/Grq
LdvXxg2nwqYplK88WwBgaPdCVAo4RHLWElWU07bRuXBTyVfnklQ7MobJkIC5H9ikN+VWrSIp52mc
11N1ZkDImcfE/kORX5Lt28Y45D1wZ8h4pOkdIjkxQGWWjNM1W8t1oU3iPDnh1CpuIZwHFLf7ixof
rTeJtFtQ8yjei2kwUd8XBY+DzerbszWllQDy6+JEVk9HofA0+yuDrMITToRlIQV7WUUfReB9NUg0
qDfcSMFOsJ7UY0vTU/+1XibQFX/vCKWGAviB6BlPcymztvH5CXb+Wx/W3tfxer4E00ik6MtfCExd
Ha659vcqPI/xGlt0z5+4bV3xUj1QDR0cXGqrkadDdZd9KbUlET8RfJnisytXBFpLiE2azE2vr0zg
J3BSAuoTglyQwWJmx/UGTF03Kjhrm/BjD+bINzGcTz6iZUawFKJRqszH9N7Re7STH4Z4akhbacz2
WPdFL+ZHCC3OIBWC0ZwGpiqhdGl6AEEL63w+Y1EpIGhDV+WXHyqi9eGgm6t3BKvpp+djbdVLk1b+
yb1r94x7qdPAaiM7BZT0YVMXtg7yLstxvQUb/5plKzE1d5YVmGicylDmSQR1hkBpPgcne9ee/gSi
LXFpYIVM9qkhvzr35NENH+McVoPfHYFuF6luNiCSa6K/lDKaHDqf470ANgffWP3iqG/6eyVScB1H
9vKQAuGs1i0G4dWRjjmnymvSo/BBp5ISUY18yc8I0OF293wkbGPNO08umfQK5rl56ufDMB6lrpBd
T80locKc6ir7RSTOPLrTgITqHDqtZZO/GWK5wK76XXndmAjKBXUSc7QYcWiDkN2rIKc5pezK+18d
EuEEOsgoQbofaC+JgXMUQYrl6dtVGw60PLeH4km98GrGdChi+KKqgwFi5K08dk7NYIPrjNIlajR+
HIyNe5tKQ/2wWsNCnYeL6Dw00D646lYFQlB13+xugCZJN8FHvGsN0Zp+oVEanoppo5YkIDJ/dbrK
7oda8XQIywVV+cxwkaEA4ebx3QhEtrTdxNXrUs2RWRuSCvARuW5rSCRMOR8fZC4aGEE+yg0ssuKN
Y/t1CKN+CiTterAzCGwIjCvXqzEOq/q4uWG7qecZWzz5PuFxfxioNam0cnX8vtv+m70QZ4j9tNZG
edrJjGASY8y6KuJyavJiJpc0aPS/+ipUdJX0G6bmEGmXRUUJMvuVmzOd2Nz7cG8RwhWRXRKnfcKu
/gpP2pRt4G1fZH6QyZfdKTyw+URMjlIHZUTxVYexjkDT7qP6KBu/jUzcPzg348Y7x6RhOA6t5oOC
XnQns6IXUTtwI0m7drKZn3pLrI3OKJGICp+pFLkmHSagBnhKE76kgvGZmxmVaJTQPZegTwzYHjZr
uA5RwzRTtkS6enZvnUCdJzoaZ6RxQA6RckrNQi7xD3MAzb3N/WKBxNI44lBTli7SxZSnk/OiG7YP
yJ4DbVVwAkeF11e/fCCodQCQUvwp8LBVNXsx7rI6TO2ksV+ygjHi+nz5hruaxemLH+pUCop04IZy
SUgf3beNjZAESbz0sioCnXiZAT4Z8mFxkdVyYpddDsQz7VGCpmYeCZU7SMXM4qGt3F5qByGsp1Zw
9r3EK448Npn3ldhd9gmjIyfM3uRB9NWuYaBRc5MpDqqwQHm+Zts0C6PoMgSCJtelwstWtQet12hK
LRLYjaDTffDIH/zsrQ57Ia58ITdWfLV4Y6s/YXzsA+Y3imvb0sTEE3zDK3ToKu00lB2kkaTnF5f4
taspno5af1PcRV+zLJgCr2ehSSuaSUppxpJ8VJBPM2wGUW8oBQbfMq146Zf8tDIj9Z/QT2eduJnf
3/EY0POfuUn4tM+l0bEZQ5Ur4Qaa8LRh7VGfWikvF/RjaCfov58pShzfKumemcfNlBWonV1qpVMu
ghMF4xG5du32lqvUR7OwnzQDhppT2K2k/URCHzBDmS6MjYdauj3XFhbBtGx2nf2Ae+cVQyjIWrIc
fHHjbv7v8Q2pY3e1ovSos7BHqVvY45ISng8/Ini6+qiS8LJYRV1A3aX8NZnE8f2VMbd4sl5SuEFm
HtdBoNSRQmOqvcDamr4i4RTTPFIO0mlJwV83O8SmyVR5T8p9S0wQRHPwLCxFo5ZboE78gE0Yj1fg
xhEgS76vnsAcdAlrk8b5uC1WR9aZuPadUtr4gb7A6H/PTtCeDXtLDYN3pz+tVkBAZH1ITq2pISFO
8cna5RK07fZqqUayVhXkCUH9hMrf4m1sL3VFkov060mzVCxP/bZVbVVs2wbG6U5ilA4iWnTWEbgQ
0qszON6ZdFovk9vt4JesQFFElCHCWqAx9hjUI0G52d5KAUru0VeH6Glvtuaf6IvbKFrrUFA7r/yW
7jDyVwKD91gj00Jig/FetX3QQ/VDESiwO0EclQnVkkLLlYhN1Yk43idE+pibwvP1AKzlzCEPb+TO
p+mHD8uB+o1sGdJ++o3XtWYajaeJPxvlJcVTyMwdiefkeiyZuazIpbbrlMmVWpRR+3APfGteHFhQ
Asx6+DvI57I9ujlHTtfED6PAC8a8zVUTpO3ljbWcNZMkePrXbYAr5zw99Nj+ssG9IA74cPMr/7kV
qK7FcsgHSTEe8t2P1n2+sQ1UXcxkcGcpkrM0GRsg6mxuewsxcm+1/vHmH2m4exxZOMQEd6/K+jZB
UFAOqzfGWndTy8md1iFmzh23877lVk6bIY8Q8wxdAaGbtfpbQNRJa3vVv7fQfaiX98IIMx3BOIJ0
/OuejAm+XOWRH52K6mZ7z62Xl8sbigZNQ/2anyohbvldFQaOImJ5q8doDyBcxGxjehmNyvphi5dk
+1sBImVPF4U9fo0TG9QH7TnOxcRnAe3F30GHjT//a7UU2RsQ/0ikooyZctNEQQ6yJYN4CVELLGs9
ylo9JvtIaXf5zc5Ufi8HFp7LoWkMu9kPkVw0R6KkWZf6tEuTdhxyVr/EVev40OmSP6lDS8ItSsMR
2iXPGtv7or5EsoJ/59P2qLfTqZ5nBy3x/3C22Jlhns5UGPXAGKSOdUe3bC4l0C5elacBo/L8iuXM
coB3lwLw64K21nz93TFoL0iB0VwdrfLzmuG0WXBQJiKeCtImEgx3PD+xrmLqNewC6LRaiEAkXm0o
8hWB2kxEH0vVL4Go92FkhqY+gANJKecWMqAzYY/P5QSNiBMLrEE4FA17MjG7FuytbVH8/xM10/tu
6duZrgbO+DsJp23lTydv880Vj7h4Jy6rHYu/7c9X7bRKpWZImG3NyQWmt7FAbPPNiC8/rOsMBvIz
Xjz4PtBFKMFrTT3YghIC0mioKUw6SUO4OFZ2lTM58747kiswED2Lf+0kOiEcZ9DeD8FMANzOmEMr
20OjaFdnrAGttFsiGLIgzrDoRwlHb/UnFaeyH/KXTiQZ3yd3Ex2HxcUCbkqTlKOePhYDj+lSs1IV
KIkSwY4uEmxJqLZCQiY/LxvKO0HAm44QyNv3DeuhRHMIokUjliIQLWFg26OakJiKDPPBS2k6BxFB
ygFeK/lTK8MldfLHYxXp3gKa7MNpQCImiRkpuIFT4SRQags2nkpsDNENW5RgqBkGsPoyszhsN2YX
MWL/PK9R4IBe7k5LZOqoyRjd/nen6IY+C3Mrmf1qpdB/5Qu4snUbb90uWCa6Ff370MNalyTyhNZi
tFx0/b3hld/+T0hFvz02XRxPBYfurdG9KlLvKg0yp/mJnsSt/xaCuCSJnAeVkyCl6crHIECb8W0A
W97pL3q00gCsVDynZu67Vp1PKXiR3EO8LimOb0Y6/IBLAS+OVa8/qGU85TH+7wgU6aMjdJmNWXU+
9nEBKv8MLDUeLPqNE+8ASuzQ2HgNk1r2+TtCkU/LJMTRHoGuFVwZLLa266FrbQ2cSZywALi6SvkP
zEscNtcQ/ZaWYk65hhyWggsn/xREvK1wjROEt6snieQOcM1u5uhOEfSyI5aTOQ8/kVqSIkWFMWHa
frUQYwvxAHzKqMNx6z4fp+IYLxL1ZN5btE4q+0OBRVZGw9SJpi40VfB5IEFmxftH7teTnjPFJKnX
KSczb9ig48bRSf2+TwUxSzhjmVSfScFMoaMchNsEUs9kz16FgvdIveRao6ugfTtxBaLiryn5tVtb
p7PIuHwFoa14AfZljmlqK6YmaGll0kI+6Kvs0KnsD9bAMNK16pU1vmW/ZAKSR0aS77nAsZ0kNGrN
4ddjO+3ti0LT5O8CqqWETMuOJtPlUQOSjddNXQ9Zg3MB3X4ExYxiJVrD/Q434j9kc1S98OyvTTar
nxIikvUGD0Kdla/3jM95mIeq7gXardNcgePOk3i8trgThUT5k2saz6Cul2F6OQZQSD0OHkrSrf6F
1tGNBOVXENu0Wa07IeLGwyUAPsqRBv8UvyuXbDIAbCfI/WRsU/xnxdEPfuAhEax2vL0wY5kJCrPv
JRBmocusoN+cVaVH8Mg5mJKiCMfm6rhiTh16MXUz6DV3v0DQZsEH++GzIh0Odwc2SECEC9VMSqSs
SXKkZiqSBYcWRtRShwHLh7eYYZt5WerAK9XkUWxvXPIUrl8FRPKzjsnZxaumvUlAQ+jN4mn1UcWd
7CUNL4b8prBaRCDODYRNp90bz7oSflGutrc8yKVmJ2kFnJn76RAF+XorHLWDfWDA9mJTX4rhJtEh
FhWpHx98pOxoglKL5CFxJxJrw09MGUalwiowHhG0QXz5wV/caOUbGgau4OTzzMRobzHbTQ3lhx0+
Sv94IlECn6gvCGjP0Ad+wkWWptrAH07LY7+yFNhfJmgqxh1bYE2xaksIbibHhJ0cHeUKxlBIXp8Q
9Fdsf7R5x0ipvTF5LGqodCX4ESmCOUcJtGVo43J3qTukBpOoBjPCKgsUjQdkM3i91Vv96Hl6VYFh
Hgp7vzRfLyUzCTB6aYPihZIeTCyedel9GRECBd6ifFIYe4KGI77OZCaAnUtHbxOlC2vjdDuP/V6j
qca603tlw1daLzrsmmR5SgKaB/LmkLCY5/Oo7mGwvvefXrp7tf9Rsx42yrhryFmm0Fh+8Ftlai2Q
/qaBur3Ot/0Aj3OoGtQb1xIiNSUGwwnbBsBJ4VMgGA3Jl+9bzdJcEutzrRIaj4h4oRjEjbXqb5yt
4YOTczgmmPKUOok65+/F+imO4QCAKDONoCizVe6L7m0EVDx9Ru3Lfy3IWZ2TDS9u+NEZXGlt9+rG
qn7yl+4BvKc/cUxPg/IbRqlSDN0CHfmXWYhL0ZSHxdJ+PlMLz/iFn91z6sQgHGdTtYJMmuYsBK22
DwlF9HWdYDAz/gbkSIr04mdN2b02Dk2fYraXj7CrQSj7aJhroO34qdjOWgx8Pwx9wgYjoW7z3pSw
4Dy0YOA+B5Yaz/mt8Rx5VCOUbhg+PGhe1QzarD0MDYwiBRYQk4Vgcz04XBRYZBBhEEuQEOk9yTWr
OorTLqTFIEaZnn8Zm6oCl+7LKXF+HTZkcEUQxYCzzzNiSkl7u+VHZuiSGcnfxUk8PHsmCrGGg82t
cdNOOVNb0yzkK3TOVWKyKlSFg6bM4yDeDgrTqs1uuwU6tCJUwPgmORUeWY71X6EAAAPVmDq7dwUR
XLhNLi5GQNvPprCByufR5qU8z6/pDVL8wuEjuVsG4w/pM/+Oe7Zef+PTUQxSWfC7WTMZ2tT/Ton9
5VTHRKG4+ZHNcry37Zq4N3+dQBIUfVABV45XNDyAxa07ame5FQhSEVTLmrGWZz6KExkDe+Xsl+8D
BrHFyjCGn/0gJEM2QHXz3St6z0Pkzua6h2Y6VPszfEL1yus6JC7gClIxSZBdClz0bH5wl9VTTi9N
Ea3ARL24PNC/dgYoER3DlwYoM64F3kSQK9oM/sudmdAUA4fy6c8TfYCYpnp4kLS+IVG6Ikn9BSoM
lhsGHMW1E+4ryjCiD9kyndkN82N5dhmcMCBCPmpHz1YDIk0rmqqxrw4tAH6DyVbJGPsqbdP+G85M
gsSgaAZSZGz1ZmWtYTvVaVKdkhfsuS892WSMYM1l8yuqPH2e6IxJLf1uJTsKj0IJNdRd9Jc4LbLA
+2KRFYZTD9eLgCzaWmD8OoI/gnZEAKzTNukHmYD5aXL3NIGzaEcyt5FLg3HLA6X++1HMbdZHCwGl
D+OJvruKb8OzNmc/dmFB18HutjSGrGHYQSb9/eUko1pLdrJsnvenP4rogOmtva639oG/ezYQthly
A41pCYwo3KHKZT20ZqQJmQ8nK1+FxJCdb1jbYg9prIYox1lHd9PwKgjYcGKycRAoxE+OXgHM2wpn
wd1L11TfM0bqXF/cBxm7+tmZpeVv+fx/pR2tAATTOvoad0GmkW1sbjcwiD6emHHw63jDRgqFal1u
OMji5LLthaLj4zZHFRRcdRix6ZK7i3JG+PhhwtbPU7B5p/jaCFAJSzSxaT3Y3IKBcpQKVjW4oKm7
HJZ/Bk6cEmjukyqRhgXPzu+ANm46T3Ju7ax4h7P7yWOR8hvavYfa5N+93Ga3kXhR42s6XvcjMkdj
TX+daH0DLQmot+yUD9Ht7R1mxmUHJ+YE/6V1aZKdNNtkfcF6nCgNmXg3bCJ6yVnTLxRLWqrT/hbw
0hyfQUe+NW7OBEqTsJapuZQyfR01SHYcDW/zijZX77Qg9q8P2VYblMBnUeSzVtLLv8R42VhCm+gR
MqinyNn/2Bkq1xDOEU+PCqUuIOwLvsxlgnADjl/XF21eUIR89PVDo+SQ67zm13Ukf9OB8IFM9ywj
ov7s8iLkHXbLedTzhb30ikouPkZWmPZ1Wse44VG9Uzk+vtNMmBPkYFmhmyfrq0A18teHCnS2mYck
svSb1ZX2Nv8q6xOAcak/yQc71984p+CS6h6Z4Lh2jY6DsHIS4ely55rs1/Osxziu356Tvv5s1RRu
rhnYyHRIt5kKC0MD8a7T2c/tmzYjDbZYUN67XCg3OWpmrPNjFjV5QE07vRNvRGibr0NMmT2YpPR8
aotVcOiVOJkykwCT6oDsVPIWU/4a9SifKwIrvFhFp3J11AEKv5203SDdCAsocJrQq82t5SQOiwuq
3ylaLNrjaECeJcsjfXn/HdOWvtQVz0ncopCQcyMoTqixheec7aOXAjgtrRx/j56DMPp9DEE1o173
LHHUWxBzg0fbjpQkDJUO2ZAR7+cx+G3OY6IFTDJGhIBd1vDSqIFcejwkS3kRkwUZogbkNvH7z88z
jiTgYqsf/inauMYwtpjEj4qlEh87QS6URoCBbRjC9LwC/XuT+SV5E9heP1QGwl61y5UELEKFahB3
fKz8TD558w0aPgTXp8Q0fwXWM7xlzCIYAIMRZpgUFu/2YIdxd8/t5i2Lk3x+d+EJuOQ+ZTWgvH9P
mIkDKIrryrpUFMd+uH7Bk8H84MpQFBj+JJdng+HgRPNqsd4e9ySMzZyFFeSO05g4EF15sjAQ9RaX
NXpbaqXLAbK9Qf7i7ufKWt6QXkkLEP6nofNdXWTAfoQhfXKW8DLzEhFDAkJuksM23ARC1TakmE5X
hycmV2/upCcit5N8AkQ83pJgooYSBm5mh61ukJhCG3mOhRfBVJPPblDyiUC/qVy0GJQjgS+H2J9o
lqPO5lYFsOx2Oi+/8ImAl1uVTUQXfitDBJSSFYoasiHNXJZGXPMp5Nsd8TlnEX2WI2wkPlxnxWgH
PlIr74PgHSxzQxtb/2jnqlLN7HXz2pq8e/vlS8tk91jZ1woOve8RD02CnruRYVJbuSSTkgKbWqN0
SiGt7fueLwcHVPzVOANess+puiRPJHNDRnkhO2Y1lmyK6mfHrPh7fH8rrde7Bis/I+HhCXjnHABk
MJW3b3wA1LImW64wDqdiHv1Bcr7TIFJqhjk1egXd8X9Y4jxNiBx1a4uCCHrEMEuUIhyfgP9cx7aJ
VowoFOAXLq7X9cldbvCQrfM/2Jl1QxMsxX6M+vB8jDagDHYN773yJ/UKTn0D+lr/XL8/HqBhebSn
pLUjmKFi4VLQ+biUrNBdX7bkq5LJABp4U0fflE1UTT3f1TsaI1oXfdrExeK3zXoRdhEd9DCEj6Eg
51/KWCePSQtDAckkalmhE2hsjqtNrO4pz20sVD+pHWpWAzKtXl4eVFBd3JteU975eCHSeBXkKW4M
7Gh9+N70xLwzGCmqPFhkuhBArDu7G0/qepY/MTid824Me7JL+xcI8TTp7siA4P0IZlTuPOyDcVTk
xBRAHIGQovMu4GhSyYBx+3/LgmelWFDZiXV32GXzgokNJzAaln6LxX6fZaJ7ENDmi4c290ozFl9Y
Epp21R+BCvhZW6mtmRZRuffNjypSGvjnMwQZVTY03zNZl92E8CnyIPXZ8+BVxHN9vUI54Rjc9Gup
V6CrKpr713fMHbyAsNP22EE19c3qlmyNBpdIonNyeOqnVm+bxzPxQetNZnxJFKkMR3yicsTO4NTE
8sGO9Ydt+jYjk0SV3INZpxzCaMbpay7HzBMqBZo1Ku4V3wWaLxylTkHroH6VzNn7B6sZrX4EMBv4
ZAe7xilpB52ht5qTr0AQrFWwt4/a+MO2xdWgZ+VSdKZ+oiy4TBNI8cSXhXqEhSO91elXwtI6zuJW
SIwcpTpCjoUEskHm26ftZfI0GT+aiSvPvlKwSKfvP6hKCXMDtoyf/E2BTUqPIUj2mO1Xhia/glOq
nW9XkNs5wXhs6AdTgPQBVfH8oHNcQzAFHK1Hv1ajKjnqmspuzhLbdp67R6Txv3XCq5A9Q8Lhj+c8
oHTOfRjiabbq6LvJe8L1x5JEYEv0J5Hr1+iTX64lUiLCRQcMlEKv/cJ+xt6tXy+q3/OZJCSfTxSL
CSsw7Nh/ZwY1ziwqzl/fgXVsji/SkaokLCNWbs95SJAq4UhmyZVsO3jg9li90Haouzh5Q1/cVFep
8xzTUAQuaiuFaDsY7HtHUM3mobcDFcbXwfHYhfZKYezQeHbEsygcLcOdtUdCgkyDiardsAZnCrQ7
4drC2O3SQH6jPF0XEWAZyuJdqZBwiAVEH2KNq8k4CBjZC8geH9Cf7hqRGBxYIWMg+oQTs9jmgWdf
2yn2p47RtNAxHaSPeg0iIL3CKMrcLS+giRZ1lJs0CC4pFm/azt5q8TISf/Zpn9rrhwZgA5aRSwFP
yKioCFtq6+ADzTww14c8Lp0ZNYRh9CHl2CGubDmf9wwAhx2hETGJdQruYdsY/GNPj6UbbMaxa4D+
OqDohN2R3w5jOBQJQn+P2PwZOIpglnlPNNJj/AtTzRMJHk/JsBIy1e49kZeXHlhCfNxfyBE0x3pl
1CmdZaZhqnxm/dQp9bPQC9xD+ZpB+VY/qdb9gmLb9nqd3+qnc2WBx+WSATLuIFa+43I25RzfnEWJ
OfWHyxo7efXvjSxw2ZXqIc9KB3LEaoLiF7u50X2XnrCsZFn9dK0bGb8cRQZOD00r+N1255nEZEV9
oaWmcLX4z7FqU3paaXl6MxV18bkLHGByeZKDjCkTbptQQqMM6uOuU2MqpeMuxDPfZ4Ekhl7dqXBX
L2BzV+XUCbLWh6WGqVZAyCmGvA2/fph+h8JBo8RRcceTG3P7aV6Cc2A0EOS5y/RFhdZY5nMjTfZq
op/Ln0K1vUH9Vb2W/VlVBssS8KpIQHL0sLypkLe7xFK+H/0QtpP62D5M5lOOFQtfjBdIydw8tFdA
ABgI5eu2nZ8+77HuKpwkZzTH2cI3SuaMR/dZXa6ZNn9CuA1GoxILAsCSrQiQd5k4gUvKMc2FccYC
Mr03hbsptj/eyjEqHXcPcrnL+M4TB1Yo5f4JPV/7Zwcb6zbcy1UAgypClnH9RhPckt6WwFwcBPrV
LJmIHFmRuz7ErJN5iz4zXqaTaVzkfk5mnvyWT1RoO45OTMLQIB+bkoDGQbUbP4UOcW00OsB3V/uc
cP0Gvc7SUrK7daMtCECR7XChi+H0mCvldNKvmygEtZktwpfScC+6s3s+1dgGmWZzLWVDN+4Tdgds
Asqk3yOMnvGjrSj0D3eJ1p7XIBe0MHg0vtGW5XbYazpughul8oI4UJxrHmHzflhI/sB8q0mPm2rx
/Ty+CyUAqHbX1KZkLH+0D7z8n7GSiODpchmGwxl3HpHXdjr3RQfEes+oMCCfIzXuO3wOaY1KFkNP
cPryH0x1vsTGFq9TjbCfFht8uHu4Gj5ICYLZYCklseh6mSeFb8Jma5mLZpTz1X9/uBpEyheZk43x
bBJNUggRIJhCCStWEcP//M0OqlTu3q4BWtnyVWZeZtGKUqoNhqGplYC/Ag0qsHO9TYUQ6NKPt7KX
hQq+pivSJopUCN3TmP47Vk5qoGZc0xyc78s9Mu5+xAoqyPcPGBFYzUGIweHIexJkmrxctmtF3loq
UuRSx3b3+X0hRPfb5+ODpGjVHJCq/YLdYl+El/1yT/2jFXxdMyNvV2gobCiKjrWk4wOiMN4mxPkQ
6PmTt5D89Iu42kCqz2BqogblTZ8i9s/NWemB8n2RZm7FpFsgdi+4lnB0Dt8PWvmF7PK5QdrLBWcX
sMz2gt8iKonBXXQ8twDspRQwBAeYVQeQXnEQh8GJgkvKc4mApvafhcSoDwzISvM07jWXMRsVdWB1
ZRIcn8Lu9CDBVwmXYF8T3FUy0bB2bjhEtF2QH8p+czMY/dJdxfa/lXPwNsoT9WGCGsZim3B3s/CV
1eNEB0JKTkOhc8tWPof1UFnredqv9sdXowPg+KvhtveWEVZ5cOVVDK1xGsNRSKjGwx1CtKFjlLra
8+i393iu4s4NTJMCH5/V5r06yx4eWdYbhr4DtfMZv7OKt4kv5NBKCsLcmZcXrZIj5fd2XAMUZE/8
Y/hQJjBdYk+cZhNhSUJ4ZIKkxxS8yNlwcJd6YtvXjWCphOTfPegoSQPNyUxAORSR5+B8xUKMjTKr
9sxzKD3sNnuOQ8XcMiBhV0s40PPLi7RHRbabVrVnGJEQMDt1e2i4ME2GqFk4BzRUjTRtvxyDGPLu
ZD5yTw59+7oR1I+X4KrCkPqApSCBlnI5tKNO08TgXjHzXw0KM1Yekg2nA8cfkNMnGbZBKsroxjyQ
VcSti6qo2tJkOlGF5rrdwNEgiz7GNY1FCaxkffJVucKS1MV/Utr8N9lXxeCasiRyPVvlXiRiQNtz
lBUlaYTR0e2B3I8rSk6hswauPEQNclOqhIWmu4ug+/5ka+safA46aqk4XEwdIRaBsRO4oKhCAFJN
pXf6k07TVClpgFbstWqp7VK4/egK1k8ZQ2acPSOYgf1dPau8j3t9tz4YNjJ2pfV0pxuNm5apMKo1
YKs5OQbc5Dewr1HTUMr0KbVYMnxzyvt6xaSNu7RunawfmM09MaoGi1MP3/2GhHXRweF2qKf+/Ndz
Mfisz+LNP95tuJyW7Jk8sSkUqP62ji46vO1Cl+Ry663ICl4sqOvna4nK0lKVkoS0R/KW35BBfV6E
Mm+Mg7+f4zO1eQ840sL4ML+ngD8Px4tT7dAy0xv7dnkr9Ul5OAgkILv0ZK/OWCbXJqYjxtw/6kk+
6zHskoeM7VOoo3jDOXOQzBK1ONsq6b+J6vkZ7N5Cq1llskKgAbra5A6mdzn2n2uqV3SOY0S2Ih0M
QnU08Q43vvptOCvtkwCKEdQnAnRvP5Tdjw79gEIzAwg2H3LgMRMdM7yMQLCE+/Wnoj7L1rAV+jL7
WWOsYSUEqVJ4+l2d0K/wFcbCLyb9oYxZrgj6Pa2Y5s8PQYA8MvLm8XYBhowun+YaG3vjPWvqgnjm
tjqM8kyRrOuKFpuQfbEFJroH0ji1pJTAvg5b6ccCt0uvPONP9K2HKp71JKdMIYLzH9iuWF4ZTmK9
JB4vftW2bsK8c8fl0smQVpatN/KSugEAFvLxChvc1zN4/BfNiPdbo/GnO4ngBplIOkDcvvdNxbes
onHVh9k5F4TtGHhmYyRZm23ZKa1pg511Gyz5eTUskoqSSIeny0yB64RhpOw/i1f1m+nGr8OjZ4Mt
kgnPkKrnltiNYd3s6iQbkNzvL3bRigqIjq3wYrGANPz1X7RVQ5UVllDjM9mS4O1ECKbGtXw27iHp
09hP9NVW/RGp6RxfClTb8WdWP2maI3YYHhU2d3+/bFRks8CKN0sO09vnDkNUhJia+v7+FGxR8cvO
mfqhbNIPros80u6+LJgd0rkeZDubBFx+QDTDfyocNcb+Wf0evyGwTUa+0AyxFbt+Z/YMfFD0O1vp
M47uhMVe7Su26hVj3zD2924eYHgEN7/9qESiDXhMsPyA5qJ6mqFLWOaPEOs2omS5roMdiocep1cM
Sk563kg563ksFt0IHF9J5IPXEnK7wPpASn92BF9P1eXAhnGowXYocv3ZbTz5VsVrXc3177ejG+Xj
YGRxFKrh9jd6S00xzK6u+lssw+AUqUuudYtneghEAcoC19FI3vhrzcy4mK1cZ4YMDY0nOoAaALP6
4eO09160gqycliR/oGwD4ZgLyOQ2DBxEPTYwotr2OuA5gkk8JMAggkYRhuc4IawF8WSm7sP0VPUs
rpNCi8Q4zzicvuwZqtMMDwJMHjdZ97f00lG9yxg/luNsXrkfEyOAWrwUSwS5ieFpg5SD2HeTir3r
5IeF3LPPhGdtETBdjkReMIb9wkU3q+aN8YT+840hR1+OPgynsNYLki+yd67QwSCptJr2sof5K1Fl
7hth9LHeebeVd5sSGr8qYNrKgXldwiyGr9ilyvo0it4kMBSUkcnUlMwqvorEEdwxOQbsngyzt4J1
j6AfvB+G/sQMaItz1YQ+Vai+LilQ1n3To6kwGO4HnKHl5UsBUTrAoOedQhcC9NACBxml3kFwWzYo
dWHmWD6VdKj4EO9yIKcXlefkOWCno9EAKLakhOplJ7qFGz+KBGuqpL/+PzWK+lv0ll5TS0IvB/Xo
kYaU0LukP9IHM1EVmiO7KLpRetz4m03zfNMjMX1OwfNs9nj7pLfx/5+ctL38QlL7y3+Totsp7q2t
danFVVtQGdKh9Zv5Nig7cYpDMKc8BHLW6Er5WEhf6XILaUvg6O/13v4TXUC/MWoE4V+DOcgGQGG/
GDOwFaDYdKDXANslosD8cDQ9v2D4zGb5Q47mtiLz9Fw0F8gJmt6fYSSH6ytfCX8nPuZuZGDCyQnm
souoamvIIYwj0FDMzEE0iHMrE474pARQIsCnYZZqz1SuF7SOScc+VvEOIA/TGYCBdGMAA/CWeZca
6oQJTXrRAxs33hF6ojcErG7NCrmL05L+wa05E92voX/doClzNqvK6PCFzByuXGOv0G5LwYJVYZ0N
tCulfvr4tFKIZepikOveAO3SzkZ3hBHD7vZWgobgZfEK3h0IImPPgM8SK6fvNPePgZP6rarp9AdT
wlCMzGsoeEru/p2N6jmyB7JQLr+MKYwOHXodhRgob7VHq0/v0WxkIJZxCktcwV46JvIBXxfd54AM
XTxWs0UdHvcXNxBEAGtWv9pHCi3ubV32/CMzkFZOblPeyKtr6p1EHnjj0GT3FzdeD6ybqE8PmZKX
99XLv1V0V4moGnatGm2x4RgjTQDr8WnaI5EM1euCs4Xcg5QQnj6r8i67jLxO+rpCOgE4XiCIlBp6
V9bFrzL+hER0xIjyTbx0G20/efKBToHuu+Skz5p/Fqx/PFV9ZiscOskiDo6MkqHNIXLDCI0a7BJH
FlY/3/kwL4S+eFFIEc6R5zbY3uDV9Fc3NCIUFf56UrMZ/yAqooBt+Lo3+RgLzyAXxI9EBeepR2HO
4lpdlPxQVtswtqYj9mjku+1qhhIXjSh4SfpjBVUD+/7DANf+tEf/vNWuy5lY6iUR8qMeC6XQ61hl
ukjDChLTbIu1F6tHBRMyoZ1sVNKvZ0g2el2ihW8MLw+TyM9c4cDrQyAGkcbBesPG6SoGFxfiK+tl
YQd1s/I7Fly64kyY2KNm5L9y1ULqZfZjkXyVuHy6gTOH65KhyQZKBhTbW7me1nDvTf6XjDA+T8Hh
K1H4jGFHwTo9XcVRPNx+YRXzdt4Q2IMaNt4DWWAR9Vcefa8u66MKHQuh+fnRyF7Fh3TkepVo/Plk
ff4+qRGzbAmHYBAKtDzedjYw3Edy2+moHuO8MWEwfKGmQGjWbsRf4m91ZHOq827X7jAghIJzDgH8
+ZY3Cok3G3gFZ++ME6Ml7ukVKlft7RRAm++dDD5vQMgzmBpIdbU6k1LuGJxj6hPvLHMHUfiltsti
FOnhbaT5nGOig8Ayh5kkIQ0Qa0PrH4kzDjrTJngJagn5cMNWnn7ylTNDbcLpVUhoeYbNAFwnNUWL
IvDUejvjU844JoV1o6dY+fVDxuRoC26b4d/L+g9VEITxMIyv39NXXJdwa80SZ1IPeyq3HwT7jhmN
LZkJ5LDNGnnfr/+Xe7SufILlOmvYYGCjO8DFKtBPYGrPWWX4dRK0oiLCsA8q5dSp3M4Hy2kFXFGu
N/fsi6MKwUafwV592ohOq921w7vzhM5TCdLm18nTv4nn+UNcvZsGvep7qmnPWnMuFXc7A78RVAwR
xuQaTL5q50ksfsCY/olZCkzpWLyh+2RJ4L0kHUTAbZCRVOPQSC8pbSmIzsrc3XYVuDWLp1vk/TaU
HyhOEo/w/FeafYFfgH1jTOYeoJDBXbN6LhcjB9IJ/2YjOIZ1Ir6kHFDo31a+hUs1pcxkVvx3+jB6
oLfyTnZqai77WPuSzvpd3JG5/5afyDNH6mExQvYjtMysh87y+6zx3DmCeSI2RSznzfTT5J/VJ16x
NHlLSljLtLhQNa/5SANIaAb+bTqx4xWLMwGeGEKwtklA6NHifClrOyP6bsyRCfltJuez7R7EgHdH
R78isOSR62/Kz4irLyNWKYyF721HnCWhteScTtVGC4XEtSEa1cOtz8gNlwvmqlq8syOXc0a4fLc2
zN4CqZU3GUuIZWhftjn9fL6MiiebfKBdit7zr8F3cqL2Ot3t6q5S0j8QAgeXjI72Qcg62lXxu/uo
/Jt08ANctIIcQ4vXK//LNhqQLZvX+InJ6JWbjTyaal8lOvKy+al3lmGVha2Rfgegbfmi76bHbOZw
h11t8xSB+sW0JzXSdACLkTtbz7IWueKf0OD7fYIwks1Uzn7Mw/SwHfrpTDsNtqtTQQkBhd4H6FXK
wvVCYhEkW6o7to2ufWDL6SI1RDVj6AkovPE8iMhOaXNSj4saA4OGDtruC9zGjslikPucSrofLm0v
QLpivL2NuboAUe+OFprk8HxcT80y0OVsjp62lmmfG3pLeMwTD8H+VmLrR9ozzgRz5n/O/tlHMHl2
uoifbtjeqYnpY45LepAkp00lCFhTzr4Y05y34lHUFV1mdGK+n3NQqQE5JN0MXNTQQQlnhkD/bkNq
VIxGJir7QwHcffvGHPvnZbTcCD/XTu+IzCHRsyZbv1TQWG1HlQY/IGOYKR+9Q8oyp2HSyObUDrdB
Rl4viK4Oi1b+TTzUAcAL5uOUEfb3Rf0j/58v5pJI/q+HFf/4c1tIc5FMXb7+LVogRMJhQkC3Ej1p
JYpGxhnv+4kVSO5xpczjSX+RXiSoOvHDrgjbSs+XoM4bvbBEAv1Emem3IHhf34gq4njX2LiNWWwm
u0c4EOH172UiZ0SfwGwXuF6eYwzGEmJDtiP0pMiC2CXAFR8XMYIefpBAVTY/tEoStJabGvqjVFZT
a+5BqmacghXjVoVF4dx7/6tzoWfcpULt0AxA7I6ojFraOuMyHherE7gjSeS6Rj3Nn6KKRrNQThgb
L8sLXIYK+eUykMoo/GNV5bbaYDs98gSbyDdYJocViDQghDbYXZYO8ik4vFplIH0N+DRN2yTtqHUs
wUfOYhPDGfKqLeR7AWkbCc11CNICZuNbhf17B8z20f1Ek4yvSVTNN+sNLTzbxZczVJtXyLWrD2Kr
2ueOeYIS3PKjuX80aLNxFxyuD6uzqvvWrzRLDp4ddYy+CeN1fH0BfEAkm3Y/BtmK//ikiHffd+VO
MB92vHBKEUEDVes840gNPxsHHkhTLrIXTODcmTQ0eJtiCFaYXQsjPnn5/eAIVgolWvV+AU+eb7K4
iIuQxhCusiQBPwwEM/cc9qxNSL214YB9lUx5TFb3G3dFAc5w2r2rL56Fd6EwJ1FLn4FwNdn3g/xo
sRgg9AE70lkLEfTpCNkVx8viJ/n8RfKqx2UchiiluuXFjV49S8mQlFfWpuZW8NwKj9Estr6SuLwp
POsJJ07kA8BTHyiGnantLJEvUqy3X19c9jSks0tGt5hAKLPHRUQ0KTUC76McBFdQHGJlQgsDeFvk
F5eA4W+bCKXMRey4G0sKD0RToHHS1z+62mKW0YvVlCsys5487QUr0pNSS4arnntXqys/OG2L9tte
Rd14oc88zMBoMz5uI7fy20gldMuxev+q0ynL5978rVxwKGZACbZjeFH3Puytuolv8aXoQG18P4N5
SIMwx7BVen2rvjpCCRv5euApq6nk6pmYLAaCS8ecioqbq+TNKxpFvwzCof6E9NP/9adbI2wB1c3B
weAAialVo05PWudTZSFNg3d4gEMAjSiQYiMnrRfK+m+tJTaKwxqmep2HwRcb0oLytgNl9eHTipJ0
szf5zFfongT8hkuPINYy7xTx4/mqdeCw+KMUoMyDdCcKwBOUWKxVE9RPSaa3e4CC99iYy6/pEJDm
RXvt7GJktvTRM4NWlmqD6Q5OO4MUs8jlFswmWDex1qgMs/36wSrUvIJK24uch0zFCVRTtsS7T1++
wcZNWOFLV+o8Av2uaFdPrapBtSu0YcKUFYKjS7Bkycy/B3IhQf1tSczSvdD06qAqUbGiJlmt9cqT
D/gbE3v2978g3qjE6z+iv86fIxcwqiBKNqoBiJrMqNPwWTDTpdO7ZId5i6l+mxLevofn+b5ktVLl
vgHczNIi+fEj9M95QEjtD4LZPPJTbgRV8Jz0Q2uouWGPdRq6wCLyatwzTD/kkDlwic0JUpZ7DDpM
AHoyr6D8lOHQUciV8+wX4OxxB19X1AQgpHoQkIeFuDPQlET5h28N60MtcB9wLDgK2ogV5hi01wJs
4iKhPFyzH23V6Hj9ES/IY0Wi1YLGVnVwMd+dN/R4Kvi5nDPF10mG2iW5aMC0SfG3/ErLVgLG2AO8
a/rMZ4TgX3jBl94n2kJ/c6OBzUPS+aRbnZRXpjjkBQEjBtw2NFOzCNnrRG7zTfAjj5S6Se4Pg5mq
pyPaIygt9YJYlQeZ4Bki/4K5A1kQEPV2r+ONMysK/oeIY7NnNR4RZesV36XTrTVN8V+4huIAoHLo
yleHk1ow1RU9p9ivV+rccEZm7hGVs93E2bUc/XeKYj5IsgIoADuUZfpPH8WseRS5s53YMipn8XCQ
Jby8dKcaYCHS65DHaAHccGZYVqhr1OAvwcn+qwUIuIRdWW0A38yabn+7FJ6oWih/Im1apdQvniVE
bPTNqtD9ZnhmgYNT1M4wGeK+JtT383X2oIWn9/OdqrL39984rN1YyT/3WjVrGFBLqoMYekxH3Pum
MC4FyTa5+nmWLtiUVmGH1nY5UQkyMe8+vRBmzLNOrsId1O13Sl0lM6HaHGFx8KZ0KSYDd7XW3KeY
VlSt7Xi0RYx6oxh46GKTJJoz0WgWeSFje6F46QQf3ues8jPESedeoVZtqIi8kXA2RX0JAJ/Q3iIi
Nz2Rzub5bI/sw5+60Kukz0hX8Rb+dgZ27ZL3/fsid5rgI52JByOBx9DTylnDOTimJqevpeZmgNin
vRIP4zuPzTpQIZ2rXa7T7GRf/3Nzm7vOj6cyRIKcTxIHc8SLAwn1srLd6OsydrXtbgW87E76mXEB
fZplDiHgz4nV91hpbGbDGCiYjyVnwH7R44y+qmGuHU6i3cK8+R3D48IHhtbxXnUewXrDL+uDWzqd
gdWFYbRnu4uNrcibOiBR4vJPHopD4KKJ9W7Kk52LqRIhUjup2frQcjsDxgtOk799DJmTlaFtKbaf
Uj9QW0Yng+JJW9KSu35CDkB+CFtXMgRwJkDOlAc7FZ0RB5x6SgQeCDqwkNHgDOecfNsl6/ZnxfTz
qSY4rb27OwOt1SdlmICo6Tq+1TQd5L5NTZ/8IZmWSLRsNEaA5yIq/7LFg0OBi1/JWeVjx3/w/00Y
EfA6lXOYoycmLh9bOK67XC+iFBMGvWlfra1GB9TkZxdCcbUbJAOpyYpc7if5WOxLfj01i22bhfbx
gnhMDO0fp+KHXb/qxN8WbOM0Qxm7ykUHRAURYI6CWXYlByi0snVli6CvUZqe89g2HmE6eIu+3PKO
FvoQ/sucNCzfp/wbIFMZ9eHKd8KNaxSumAzeJoMRxh8EYkvIHFnHGJ0dfaMakRcK2PYsjqLx22Y3
A7zU3abY33Ym6N8RMmlhdRedeu5Nf/VmlYygKy4ATye5bEfAJcTNBjK40333QOAR41A7O2qu5jKw
y0lyyiMJoU+40hDVntEHXuuLKhOX6LqTTTSMd/8ZRy15S2AlKer3hgjZ2XIDZ6e5UxYDq9z0EKuy
n3QsRfDU11BupZZ+pIGE7zmUPg/U358s5B0LbsjAOepddfSlBhztoEj83XL+LTxtCfzhlOfFpmba
9akJ8sXR+xuWSexMjIdMvu+ZAi+O7mf20QPl9RDpcsgOKrT1A9E4mrr+s2ko5ZVbrihBr9s+Q0//
5hR9wM87JhaB5x93weHmMVAbhyeMmuCA+riNKaGlpREoKJ9aH5Vu5+/kimPF+rOiZd+axYoWC+B1
FdgcwxlB3hYUO6OC3Y5oXgYTYcS3+Y1chilkBEky8Hb+KyQHjy3IKY03jk0LxjHql6nfbN/NfTcU
bjwMLiAkCLt0yc0G+kLPa5u4eXkGHYoSiXfhPStbqHfGCZ6Cc2SpxN28pvcnpp4ZB0yw+Kue2TAh
nt01cNOC9jFe/i6RO71k7ktk78fTsl4K0W5j8RN8e5exV8GqS4ftYDmW06qeBkOBJr1OTu64yKDI
btHUi9oiSR3KnEc3ppuEVKv887aYtXEZygD6wH0kfErg68EH131ipGGs/z4wz9XTDfxEawI4Xx2a
82tPsuFCFCD+W9Byw3PGiYV5bc2ER9AMg14FcRSYZbJN9Wz0t9VWPjCkOIDOjOk0UvCqO+VYdi22
ncbhTH1FrEUEKpRMBoJPqj6XLFa6OzX1unb5sjnWE6DNY5ta9kOMsLnWu0xauhhin4n5Gt1qpCGm
f4Adk8bNOy51mXoVKbMIG0q9UTtr+LRfNH1WvJNIh/nrFPbfmixLGmF9UHMEdaUPKJ8H0q817p9+
PQ0LL/uGXDGO6tWB6BpOYP296oMTVPCzGB1cMBnqAslhvqTYcRkhzCv5odUgXwsRzh0ZAQ8TbhoU
fZwt217uvYZNFFHRJ/7i514LIVia9AJiuXYztfj+iBONkNAcW3T0sGjJErA55ZOKg9Bf1p0X00dB
3NIZJFV/S7x2zlszK0paBSbo2y++7lPljX1Ih8Lj+zvIPWw5loxm3B9YsD+q6Q/Ph9zgl77bK1RS
Ff6Fo7VlvHEsx59rCJqm2D2zOZCL+WHfJBmHXRmUZ5FpogqQNg6rjWDRrL8pZ3gak+BqzwkgJXkj
qow910x2z+023DUMqGe8BgTyFJ5IaxMf9TUHCoZQqeVtQlie+aYD5uUBQ6dpsw5Tf7Y+FbWQnyEj
dLOogNZx2olnke0Rcg17JEdIR7BrxDwEa5Gypxu2s00EWhfsV2wtp3SD3blm/ARw8AKic3cjn3g2
dxqIj6PzHJbNdIbXpMYwMLYThU2jHglVjnsEkVsblGW2+1lQGLhB4dE71t0KSuCQ4VVkxsefOwML
1ysqRs9GnJuFKLyHWdc2lLXyxUf923+Ca/X4Itp+8y+O/pDct5w83huFAKn7TuQu+NZ1p1BDLwQq
af0fmxSJ+4f2TYInSllD66kpM0CZWGDzf4d7qz0WhQucEvVvv0hISnYaWw9Rpty/UAP7PS3LWRIT
QQ5JTNyeIq58hm+4wJ30BXYMBI2Xg3qaQgQx8zowNIjaUvH40Ak6sWCuNM1Vf2wVe+Lb3G6Y5pDZ
HI7YTGKOv2SpqY8aKGZK0If0EvEsZbg0bbOdSJ6CXz14XpRq+dK+Jjea30NrqlLYMUS1kEjUvAnh
x18SCwJJ/944HyNcBbauWzwAZaPfNSTLKigx9Q52puKwjERwBfVWcPnqRCgMPgKpPa8k3lycrtil
ZIcSBVYdiFLMU9kuOowplEUQsYMf0weHDLJg87gheYReS1BudyWbBkHjRRbwCDsWU6cIyJbwbSwD
5lNfdOZgJa9JpOUj8f4gpfT4BbGbbkJvGraqKAkhzs3Ts+ldGdT0FSgIBjdYrN09WSa+3Tc7OBbe
ecvbxc1dL5+5ETvXIzA2cr+KTBfbiUad6fme22yF2/xhi0RsMu3dhJ0qYPrKRGzIUg3W7EJWPngV
BHYSlRJJDso0Nd0fG8wtg1JVjAIC82ayYxo13R9r8pQCZdS4+mI4sNA1ARCU/183tbpBvPHClnvO
UY9RrJwW4gk1+JiW2kKvBxnzAYq2PSvv0MqA6u9FusFSN1e2CdAQf/UCwkUhrDqWxt86SoTNN5bG
xpXABLFvQ5QVYlxeVLzxqZdUXXj4mbuIVldlsHMOgqk8+9PGA2OyWxAa2SH67WFoXMWerz8h6z3r
An5L+4DDNZb4Vjhpg93+TNg2I6pbmQSUK+p81MYVIHEVFV4mMicqY1/KauK+flGPqhsuWNxyW4rn
I1Z25UB8dws1kPXc1zyFTy39uuVpCqBM+bhPHXPgyxqbnbTOU75XftZf2RsH1scjxBE6sBUbX5NK
V1eNc+lPN3mqpQoW2ksvvkg59mVWlLuFkiFDVcpz8voz9RZnmoc5TbFphEdnqbYnnEdXyzzU8ECA
vYB4DwNgAMyEABa+RaveJsDgb3zvl3qe1mU/m05wlYGOFbow4zXb0yAhcVD80wF1a7tk6gBuhJYP
uH23IDp8yBtsMHLIIs2vfBUCze7UZR1VT9Oxw7WrDm4ci1KJ+9FzT1EmA759l/MeYbXcYlyDYr/K
sJtxKFCXZk6ZhOaXIF7drFUaUlvk9mIiLVGW5lNnLIBrOG3a5/3KPXqcD9qQJn55fL9IMnj1vrkI
CObVzK2STq7Qu2Qibs7tuwpDygk5AAfFw+yrPVVHoNHscjLbB2DfYnqMyJah8OY8sKVc5MvWydE3
ptqClMjcsRk9wK9JSQFNqzGMntiMRdbtXhUOyegT6MWN3tvOpNzMc/04P51XDJh5eSQdPaekiYJz
Buzj/yGuZ04u2403d1v5alGZUA5lvJW5jwtSPcdKu+MfHPU8xLcvA9LBBmUQJRa53/S/kn+82oCR
FdYgdtfGC6pVUEgFsa0WdgHlng4PMIamDjpO4S6vbFqEMSRMSeM6yo8TfMF7JC4K1xiJAXCHveup
gnMA43+VYsCHAlqlKMh4Sqv2JJPQDnXS104bVqovNHmOm9TnT+wlzlXSAVRYJY7wORjSFgHcRU3o
ivz2C7qBEuttZ0fkuAaPmhR1zeTSHo45aqx3TrwmOeuz60/kHoJJ5ilFb/3aNxKEqgg/VIjSU76m
lfoiNLpUuw2HzvcC3Vo5o6hj0AW/PjVP+yzAZavDCSOUW2+hfLEuH+fdwq0L86LQhHKcpHqC4ndR
XgwJex2lE+KyEh4g+yMQiVr5vtBYxEfqbh2YYyPZ4TOkpn7oMW41pxrGuMyoJ8sEePBNfqZstAQ8
SneUJ3r+2+lgg7rymcjmmSPVCwM0bGjSWa+N3NjJMs4HZkN8LOxzzv1GMJ0u7G4d0QFsmFak62es
xNORK1jscgwKnIz3VT7BBVWe2n1MsK59ibHdfdgSWPcgFGVTQYMIOGafZNzGPKucnxCbmisMVk3h
ca2cRHezdk8hrivQGuGoH8N0M8sUfa6O0h26F2IbtzZBG+z5eqfUjveMFofFbP3haRpV5zFUnjRi
Ei4thHZk3eVg8v+Tjw1Ce8hpALiIlt0Gc1HPO6SLGaPrfAVmwOvFqC34jwDoyEcIswhwMSyBU3k3
wu2La6cP1U9oTh0Jg8JTbd230NDSNYZrjepFyJasdckh0H3E1De/g32tZEyz2CGFaXIuGE4Ih9fY
9ejI0tq2rqwTUPaJrJ7Iukjoc99zOtck0UOLueST1uS19nDbvujeTCmY6WYbvNkxPULSJH5oqEe5
0ftDZ0bYzJ/POljzkM+6ps5qneXKm6+GVGqcnYtHVjpcl1qBfjD9xHQomvSJBXLG5P5r5eJ5QPGC
Iwsv7socXu/gj4hDVoNlCz8hT9Ueh3k+3tkU/c25nVIB5RJTCbc/QjvgENKRNL16LfVErNo0BAvG
wyk0zoWZEmw4zFsbsn58Tz7Cc4Z9mKInqEnMh67VT4vKGpzQAXUvBF/0UKPEruqYmravq+wgRq8K
Dr+m8o+fE328tJY7q+BTo+zD/hZyuPvtpiGSeDxBdFTHe3FGQS3pRSFiTaIrP9zuszYfFqVJT0Tr
nq3n3y+4gXJxMaKM5qUHd+1wBVdDG7uBA6NsgGxitG369YgrW0kZQxYBFzqkLXZqerIRO4H0O0QC
Pts3v1hiPampeijLO79oQLdd1l6spHl7HL3/kUZMXQDpmJ6m1wKXUa6Ft09qrsPN6b2+w5kdXtUY
ffw0tiEGKnvHJrMDcdu2cugS5lkESst3zl5U6+nkqE8Xn3LDEJVs3qivqICps9rnJH6RofutPkQB
ZD983pPpraq21ikqm0liMYzRlLGafRODv3dF3dUH8+SYUkHEnCuhMhMwqvRq9LkoKbqlXYwZGrbp
WHxfvSvGXA8D/Znzq8ArkXPfSMJ5Df3vw1CXUalN60lt2gRm/1WWXHCPE9w339hs93mA8VQoWARg
rSCtm9x4hOuXwac51iaJSqTFrHcO0eqYgb3zAEZXy1AT32WPgVP/e3HkH9AWrYu48NANGXLN7tYN
JN8kwypaVxkEoSNyaF1V7IxYqeqTWB/VKz9CALwssg8aKsVdb9ROsc259FnDTfI8d9KzB3KKiWxU
j8KwqRMOhyMZGxWIfWkzb2bpUY2i5J4Zoy6EJPhsI69DMgyoLCQlfq2Up08laE7fHNclPpCtdoe3
yMvT3HApkyUe+W65vxCW3tOWwaALqCWhKsIqFxbcOBb3bQp5sTRdmJxxBCnWIEhTBDNxOHTvNVaP
rkMWY4yV7DkcHlsUSR2LedLOICcfLTOqLLYLD4CxUIMm09WUNMNbdtfGRx7u8UCe3kFGcluo65pj
os5/AfRAG3CcahEwd6q+kxGauPr0P80DwfAyq3FtvdqMCtUzoxSn7Gf/ZSgkUHxT7I6vjPuncS3W
TZlaf/48A8xtGjiPoJEF2vfmiHpPBvP2HcvojwBEm57fClNaxgspSgG6t8sWJy9f5WTLhhHHTu8f
8jr/4G6RakctY4EAuXz3lmHS8XT5X+mYvmkVA/Vo1W6KEWRsDBpowU263bS695ESwX264ZTvGrlj
/pdLBKLoyg/v4e11VZuxiEnQs8HEOCnwEFIygnagseISp7X9YlELqWO1Xl5kdunfetXoiz1/6NMF
j25+P9+MMuzZBqjlDIL57sTythFCQRUsOa9gfM4Xnx44nYn2MNQcGooPVytZ4ZurMNXmsfcZRvMO
UilWNeLoTG3wojSqnu5BnOSXRjkonSxado0ntQzyK1qA0JxtvuFy9zFus5nYi0omxO+y9ApPyZKI
9Hcqb8cy9v+qJueZ/LooU/3kRPK02FO85dLwIbXwc/ILiWzR2l3q7koh8Obvat6G5yJBX1iwqfwq
ykW++QjPRvzXFgwhOry2XaqKo8EitKy8ZhQgOxjZ0ulKoqloajCisvOgdMjiP9iA/02HWCgsFdNi
jRVCIWWdsuIA9CImrDwGsikHLxpqaNyZOcFGMRxmYou0WCJXwwEIuHH3iwJ8mDUJaegO/4zLJMQ5
pc+EPtG2zMYKlIy214JUPkI+X9R7Nf7rdfiMJBdyOWtKmbztspMagtYQJTEELC6AVtwxZgCw8cgj
4LwhktN1bMP1Vgieo+ac1E9NXsbhrSwEtSBk7Bd6lEQecfwjzDyq5L/+NatYDYJU0K0BP6nhuIxO
YrOl6d8q0ziRoVUVsbKQmXdA6gzc5C7eSAEFdkGcwHy94NVXUUAU8KL2pIhsWo4z9B8TRc1yRVAG
TEsb6iJQYPVQu5HkWSw0i2zkZSRtHdzNbqFEu2iuqDPPAdqsVdx3dIG1pEXBPdD8O6hYp00phWEG
wohi6ZaBzt4hJ8xaD/LwkxcBOf8D54HPGsisVz4mq+EBWC1+Ib+JPtLXiqMW+F5gaitXVGEoQqPJ
h0G1s7y09bCZ0vfoupmb4ML0AeBhpt0AyavtHS/+8Io1K6smanBLcYqgR5juQtthUWVfpqI9BIds
Min4OGzP2JqWdwK24n2cT0cpplecM8oWrelqsjzizB2tnMZaPJIyviYBt6/U8CqDQERlDCYmKDXG
PdBIZkeP7uABJTDwtL7V9VeWcIMonb0Tw7AfnEXYfo8P9ckHXTORbCB1UuOQxB2CEBE9qdZIgwse
H/PBUkS45RgH0z7NdniRnujZZ/IGADWRzxpl0S91VMhLPll4m6D+3pacbGeyciGnO+kwscvq2XL6
1VygBU/uVvIbPnXzk+dMTQihQ48Geu9shDN8Ze88a0Q7odWgMGqb8bmO6y7iBQzbiKj1imuvzebq
hI7AFIvYbUhkzoFAd/WCfDmqo9jVrf2Ea2fEdUERAJouOkGAmKSjSTLAvSSYYPySBPI90pnqwFJN
JiPSdwJxYwA5L08nYl9Ojp6FRg5dopFM6aUEpJRVod1mfAgcIl8Lxb7lpb3Ic0m5QuFDOSDh2USo
A2vq51A/lF/MbVsHjeD9JkBJXV2Hd3P8P1CzQX8/0oyrY3ieD+h+B0s4yhplKcRhi5mfZc+CQCbX
TAKn8o3fDMRAa0qY3PItEJE7D2ssrmSrqbrSjb60/C+QQSx0Jx6DbosKxNKiEgQyyA8+pIljGc4q
TE29Rr2DK51P88RaT0lwLyYjpCW7MTsNgeOqslhgIb2VvDiESq5RaGD4DYhcq398y+awrgYV982L
hXLKC3+TQKc9lqac6YdFGylHk9/9YlAZOA2GM2DQjv6FSDNY9G9Mhxhk/5KBNMmKf6rAAxEAOqe1
RINCFWdXfmQu+x7jMHCZTm4Ui0TAnn4XtkkZPx5Hqfk2+8HezJwET/6s2Utsz5RF330x/tlu+Add
6YzRRTz/vkIal/c6ZSqS/ED0OAvQtiFLKA+Y/JsF+T4E6Y8s8f0DSRjXK8S3ZKJhYe+8mBIv/KAl
LgVXyWAKrMnmUVAECrNL91sbkYVKbUE/U0VIu6AOJeTZeq7YON8SA03+KQgiIuv9ceDuuSajYKO1
IpX2a8/wz72PztiTarf6PZ0N+l9bDYwCBXzOxwfpfE0hDucNIRNQ2fWJdHVyC9lptW1YAtIP0UqI
jG70HC+HLsYZdqFuVVpZw0pESO4W9dEZ+YnAnicGshtTueHvRc/mKqcjMeWE7rnd20XDypIEsYVV
Jiz1Ut1X0c9gPkOadEBAzyDP66nVrtFiFQot9UnX1HubGJGJ1t58aXG7ejTHctpfYFze8fbYK9zW
wRQgjWBnEK8MzfHP9rVPOfKL+kuCAOT3fQmbI1cQMPXXl40Q5CUi0xOQSGN2sT9gd22d9BCPUW6F
77bM4yvl1a6qOe0udtEeIAObwAefo/s65j4YzycAA8arl8rs4aavqNvL8oZ/RkCc/rEOCepAAxnR
fF+H/ZPmvoC5dD5fG/Li+JeUWLHzOxlNVO1GbsSlP2QvyJdgMOpqJLA/L8RXuHalxsuYCF+Frd6W
HSni7fgNkZXFQGW/ZQ4/Gztq/JsFrjuYQuzKN/k3C0Tek2AtB07Rj8zApp8midqVdmbqUYZUMvHG
YGKhrwFMw+vefo5R5eJtU7OvKBZBKtqucKHUL1P6Rw9o0oMyk7lUly6iexdEbSdMnB82/iCCBaFk
OvPXLsKvPXofz+twJihTFzVDzuzOCCwMHjer8a/U1Cfcaum7A7lA3a+kao6YCL+uu2cgJ2ZN2Kg0
yL0qCa9RSH/LN3BPUdfiUVYEKJHhZdz5pFho6vpILRw6jdRV8tdCGi3DAulj+ujuxeYF8Djws9Xg
cjR2jrRLaupIXzP8zsm9vr4m7/QRSqWQEap0OEchN2Xq7GCjX24mjy6tMfubw+vVFUXbCDjgGwBt
+5TvNfxcPw0CzPUZPyMaZkOXeW9TqiBc+p9PV8DRSsJmT9PLtdhhSPJUdvuj6h1jxnxfg/KZ4ZpU
PQKh0T5KXB0jaHe/AV2DBaKrCfKO7wWe7j/oFzMMFN6b2h4XGBcTYnxllcU+HYZQqA+UF1MNB95q
O3udMbTNImAPg8kLnRl7ptG7Dgzpa3zDayzAOlT8RHzJRVKzYb8lA0o9DStYAyoM6J4vkzNiwwri
6lj+9ZX4K8YNEc8oJT5+41as3Eq6RYMxqzLW2W52Aj2fQ5RzQnmf4b2GcOoSs8zJoaf9huj7EklS
We6Ip9LOV9KlphfRyiS7DeQKU5f7gQmOBTTB7eMNW9kunj1lt1Jp/DF7X5b1lsxgohvc64rlygSj
KaK9lNcrPJeIu+ngCFdl1pbOPQ5GsLmRhmkzj/qmNpb8Xt+o8E6tOwPiVt6LnyTlfWGe3UzG5TQf
IZG7FWFzIBrh8+Tx8hlX2hx1QXIlkZQqa0DTonKzbyR8xieCMj8KhX7fkuBM2jqvPdJOKNcVzKlg
2bDq4uS71+/8R2a5bF5/IblRDb1Nany4lhRa1a97uglY2iF4GD9pf48XGzJEAWEuwuO3IOwtWnBS
naggnR65LWOpn7Xe6Su6rWhgVVyl3oi76LdffxBxoOvPgttsKoHtyQ4bsmU5GIcAMhhIsowHALYE
5YdZ7aZEG3q2fY1Ge7YbuLXu3AFTzMa8UMtwEt864x/KxQZ9SrvW/FVfTvRrilGFfzJ3FIm7pZu6
45IL6yNN1BkgpInN/MHH0mnuXI29nDNOgHKZh4xSj0bu0/7vFEPXLC6K6Och02hZyJVHUTUdz9U4
2OyYDXof4inNwQSN8xJSPYtT/DtljhGx+CKWbwWul9YyaeMoVIIkD247KylHa7313urbLpZK5ick
LXboQrVu2q+ViuAZaZrJ46VW12Yu4fx6lmLu3ovpnXFezFuNZ1LWLaGLE8qGWYfkADDPN9Yr6lHl
83ZutFtLG2W3cDD61R0r92P/tVSqJHDfhppMiTsuiTNmQbs+xPGVAPiruWfkr/zZXJ+ajGC2xrbX
4SOqtnRsXHBkR1h5EdQKazpPeIEx296h59NY+egne586Gfzh9RPe1r/s880jGZi4orjcegJpWzi7
cLUw1u22yUa6xdJK3d1bHACGnL45OFfV2J4g2VNfMAd+p9a2sYR1vqc6bMhFA6DxxCcV/Yyrp7IX
dcJhf7f4AFk5vY+nXUCytFuCKdZA6AFcUdo9kBRvixkGZCfQich8ThGUTNODFyh1w2uhE+haiodF
iTIAJnxBFh6UpO/vwlmmuXyrz1Jhc9RJLDCFGIX9Nvpq9psf3iFCLdhekHAIc7kjfzxGlkcZzP4d
xg3OHJajjeFFISKCtE+E8onuzLkTSN3gLOSNDb10ai414/wuLtjFBlvA4DgBBrzNJHwPuS6p7w23
N78JXJ5dzG7UPvW+hi+DFsQwTNE5aCShC4rGaeK08VbzqhWYrg6Xx8IJNfoGc//bJ5yQfe8c1wBP
WuLsQcvXlDTL/N3IzFXI3g+eO3uQY1S15N1JVDHIYT9LOlkSURkYejiVcSz9C+IZThS+H+KAFkQz
HojaVh+OjrbbRRA304rRcWypoW6plc+YBDKM8KqsyYGNVh3GcgtnnidBUFu/nopjzKCDAFdQ4BRu
VnGxPF8EXplrAQxYfKEsFqjSvO2sld7tNQZp9HyRUl8+3CsFGkWisjMmSaZAitlALofJtVaNoL9N
gOoIBC/piFooMvoF1Ew9Yo/pJuvkaf9Fv48Wr05d/yXkSrIiXw+QPiYyC7QIqTB45KyXoovMzKBp
zhczD3YPdejJwWiTW81WxzjABlaB5tWW+IIywpcM+1rF44KLbZWtTnxPQnPF3F8j9O6bYRIa/IjB
RR/hSpPlY77FMSO9Ef9rx/zcZFT9cvW1wl+MdkMUEH1lqyH7GYzIw6AshFPwhzQeBtV7ejyNnpfW
4iFerZs50BwoBwew2NN9nJCt8ubaNp1s1WDHdvrhokrj3q5Dc3T3LR7dn9K+faEYvGfHS7r2PZ3S
43Tzv5ttATiTfRKvm/9Ug1ehbsBrxMLzZy3H8+h7OBzBhVLKOVhzW7UG1d/2eQqXt7hDE998Siib
BsmIovkAS2VuHq6mAM9x7Bz5JKVGMUFy9g4RkLzN+aicO+6AOKJyWaGrm1qRbxRWLiFrE3Ppkmb4
4Ul39CDy+3kHvYRblkiu/v3ngsnHVqv9l+NcPXjDG1fWhxJJya9uEy5JCGwlAV6aJRrQ/Wn/q77i
R/rEibDJONZngNkjRoP5G+9hNTGblqbUH9DDfsNeFwdUpK50wKJHNbJNeeQfHwpnzTX6pevb/DkL
T5NwQG8Tut8G2OgGgOc2pGVdjIVSoi7vZHBbI2jpNnrr6+rKUtbAQOsMc5SUcZYc7zvU12zcbtz0
GgQzc4Gv3G2vjpuZA9cONKgT4tLF6UZsamsL07l8yksEwAyttWIKdU+gIXsPspK5H9LbJ49UuXNp
fxc+171sCFCSBfl6BTRTjw9rGdnjkB5pSHH0pV7jFDWkQPgogoVzqg6Vt0mf95MsDj84iUgyu7TT
66/1jQP7y1+yXITRKqlMRtGWqcsYhuOHajc/MSuHIvntEPy8M+r7NNTdAQrHz1M0vbR3kLLgcY7j
JD2rwxxclcZH6zxpLefX4TOPoEW941lWQ/FY9J6LXKS+xHBJHngUrD4XyzBIa1mZL4y4XjRhU756
J5cglKJaOjJkHCuStxaB26wyf9SE6JWaCZCWsLpM6HbdSHXoBZ0LNGQ44yETRGdUHAjLBbgwpkYY
WQ7cgXER4zsX7sky53zEA0O1fN2OJFRzYQ8s7wPy7K2fV1g0mHF/MvdIDQFdP4ezLZx4jjUBf2Hm
WmHvignkDJyMPttS6+blVIZkjHdibpKgVQkzEMjMovy/QXnTEbLN7dDWLkZfQ8u8TWJ3Pwo7CKJ+
FElSwwaNG3oryMTKFGWNRHAKuiPJ1xrMyoWAgMSLMBrtv6j3OQIcLZfKkvlDDdj1lhL+EokAXoyc
TZqrk0RoQu40lo996kBKZH/flRFL9OI7n4HMZriwEI7tykSeCfNidojYDqsKi4VW3nTBLalxgsbZ
IQx1ZG002dg6ybz+FA+cfyO+eRBqLQC5pAztsAHFomcWFBNrnaahYfdTjLjUN5GaME7RS+KObo4b
cwOoOT0wrBrAAGvZFTOzhIqtNG1cWF6CGFj4VEURViUd+cNnEEfDnry6D8ud8108fsgsRVA0B1sV
RO9vbwxj3ZTgaVxz/rW4B00RvgfxFb6EXKfWwmQe41eASWIP3CuyLcrt8pRkPU+oD3dL+ceivrVo
6oh4gZIcrWdA2LmpP1U9dVCQJYc+rP+XY4irRTcRJpxKL3jJ/gqSZ3yPQEtjItPevFlZZZh773OF
+ZDqUiz7tsVmM8zBXKtqA/c5H04jBVAGUYAgKW1dv6SEu4bjV0W8CIJ0QoxlmUikVQnA2M434812
k697XwKVCu4M2euiFSJdi1mZjOQpuUg/Y1sHmknaYRqar6uijLxjnCFLqPToOBdTUvjWhi+jKb64
DXBBPk6DEIn/68WS2RJljdaNGWalBapHOOaapQi+DB9sycD7shL1DDJQY/InjJ6HA/kAbtwl0IAY
POIgYVWQ71mH9vuJ4Z5yjF331FGzJHfVd6nmmDGVgypoTY+CzKy0aVPOhN/FlgJiSmvM02TzJT6j
hUa3rSxoP6FduKipUgj+y4CGIgpa2+J41hQLYGgMcuC40k57FMYveDKF+zc9MCDkM51gBgKulO64
pZOhseQ+WdeGy+6dl2KGnK/ceR4tSXBQ5nddryBYkncDiNPzDjbOStbKX900biPAvNPwwaoMFmLn
oXq9/W8S1+xcSCMWgCofVCoajpiuTPDaCyaToyDBzBdZUq7ZqVUsGzrM2Qlepw6zn32ZDzkTkxFz
7fONLQrnE8H/uUXTs3YbpwfVEcipbnTwvK3i0L5ZS65fQ8/wFN/wns6IUlGrgWirlPQPUrsMuUK4
XXCH0BEdqzdlNSUorR6LHtXTXbzbAtbcI+595TXMrbZnisLyFv85/YGhQaGTc9O+mBpkjZYc/Y09
3wNJh9GZ/30ajZjaQnG+rtGmV8OXSbMb1G0rdl/4RtvIL5MGT9cYM+fuMxk4TjGJFsftKp4OPjvC
XAolQH+LSQS+qqiEqZ96E9hZfrej4ehbe/Uy5Ek8EV5dWAuk//iTXJ/baTmCi9WSOGPzTFzvHJ+G
/WRVKbWcVILI+CfsPN6vIAfbwVMnKwWYUsSskrMJdxne6bbyhCQ44XmcKnC1hoMIaCbUzcI8HvxD
/jk1aHuaVaIdDFtJL5bw4SstJg1r6om2pau4wt9g5Cu805g106hjNfgVVpbKiqbuOWV3xctFeZTb
KaVvi91FU/BRIEBgOURgK1a29jkCP4gQTRVnjaWhAjK2iZOnageaoNLwAPQMBPLGQmLXMmVsvRDU
InCnca2M01d1V6ji84cSmJl32sWyRZYYn/w4jHv3sOqPjo3JeI8OjzcCfGxF4EcyByNb8Ngity7e
Grx5jPM43ts964LtwGif9VmD2BbTJWArLOA+nYv5cBqu5MXiNlfNst6wi1JAYfG3c00REpL8OUMq
GXJPxKUZC8ss+XF+tnzZnY4yzVJRcGPb1ZhPt6T9LKE6gx/N9ArxbuYFDirefsoZHLzFI7P3lFqT
QGcwLlxm1NeOMovxIemspX7entyOnoEAaicIBfxjZkPxo9hFKcIs4oE9Ub5lUT+GciZiTfdpIZop
pH4Yv0G8cRw9nb7lYScb6pFaPfrIt3FmyTNBctAVT5yCFhEGgEM8hiMqb5i/rhgWJliltnVFCNXh
sCS93lS5Oe3hgF2JTXU5kftIcRxFzObLy6/KoWcJscoo7OLZ+goFHypz6thnjEUblwfpMa/mM6JE
YxkUwqC3aT+CqX/zSaPikj58rb8bpnz5Sv0csFRPOlSx7v8V/OT1bmCCtaja+42eJV9e1uGlMxbI
pQKeYxf6gh3NcLoHwZ3+eVAtTzEQxu5Cewlui7gkgpL5gmMXPr9jZ9Pj15+Qif8cJ+2uf2NB7UPC
dnSiHon5hGF2CdUEqnsYwBmlHFnhizmQ47w7GNlzrvwUupKPE5hNR8Vam0WtdMa9mw0SdH3S420b
78MSH5+TjZwUqR4BdXUJzmABdR0n/oN89zOgXVJlOTmIk4Ci8HqD930AnoyavmgOScn/nByDyxAr
k1pSSDndkAyoXUCRcuhFURo3oyk9RjnXtu4H1w4p3XPAxVnkADxtne/RZ+52uTg/za5I2YL+qdSK
iBxxtIqQQWJSVGR1laIuSDtNhuLUxMJzCFIHyBvndslYg+wz6hgb+SyI0zcG/ySvN62hcOJz3alF
M6hzwJWg2Ibfntr4fxKh5xSRSTlXVsbNe8TVMHtFNmYU+iDCJN7/C5a9eY7NlwcO2fykPqH+62J0
aO9kq3LB9iWUptAaQw6Vm6mfQHvaynZWFojPidps2Fv16kh9tRCtDh4pcpyLNBo+o+sm+lm72SPd
ghd+FvhSiA8nLZhJesyBcY8mBiTUqvM7UKpfLSu5NXN3mGFAc3tOsy0xQj1bjokq9qBx6Mqi0BhV
s4Z9EapkMlUx70cBtqecOMPun7IbtM76dl6rSY1bwfVk0vAn+vQA+BBtswnPfIgsmO0JmV2v0iCy
bhqJid2oRj/jd+rEYMstnLj0xJLa1bExy2I+/yJnZr8U1A6PlwFv5YGXThW+JO4/lqSSjVXwYJlW
1pc5Zg6lYCZpN5m9gzmNkBC4gElKyJZXrEeZ5iA3b2miSy8mEsHipSzHf/xHLyml/xKtxmyNxHgk
D4MWkpWLnfyoQ1WWBSmae8W/u8FsVyWl5cDB3ophe2icXh+4M2D6HQwzZKwylTlOY3ssKzoQdHKa
HI6DGl7qTUvrmEXkVkwdKtrDkuwyf8+BoGQuVfVNv9bZNkoE2NKe32dEnB2FOjsVGcOpEZCT1KMY
Y7bG/n793XWE3KTlnUC8jH0fxWnkUFVD3MYrS+vXS8TezdJWdCchwcKcfqg9j72PgODRNZjaq8eo
fu2ilhpoYso7U7psrjhzLlpfL4jXEluYXyr3oJJq+zW6kENLTS8kXRgZEVvZwrAG6318qJxKEf/K
cQs2xKAWAqeDDg4IppzGHowZXcGQlmn1mFlcQg1AqO3PBgm/F7im0FEV6U5eL+jmW3gmlHUh6IEX
vo2f9Xl91vndkwNfaAIT8ipOny6+rpLmBt07gUaZ3Jqrw184tKPDtQ+ojIYDG43upSDSvcwXiJff
1LNB5Mxnsq0qJmfjwIbB3JGEfOlgZxFMSoYiPAa+0uRaZv4I8bndmtz2njts/A6WLZ/JMNqTIKZo
7Vkwca2gg2Ke5xKWvnKDjKmh9g4zEcMDbcPt6c3pcx1xXe7dxg3Sic68BmvDGyoe0A1wPW3EOljn
w1rNRYQ4F+VTviK0dtprC6jj97DFbzYKT0z4GD7Z7QlmMjD8P90L9u7epZpky97cMWmrFEjIoAvy
jqb5UfnFrOl123fP1X5D0WdHezWk0blRwm1IhWTht9779WDrzhOm5CecnNl35AFa3It/ravtU6uK
pX03X9hwPkzIoeTT2Jjgk5t7QLP9C6hTMk/HlcQc9ZbnP6xr2TRxKj4dbKgTGt7E4C7Dllt9b0e8
/Uc3hhKrVhWAvn03OEUn0lYJ/OtEkHVJHXTfSUVZxKYgd0K7NZGGk5EwqkniDqL3UR0qyYCQRQlz
pCyFfgZuwdoqxezsGdXFXOVtN+FcJCtNy0aSKlkDZzYtZP4Iu/OS9beNATk6yh0c83O8hEO2qwlB
pwwD606aWKEZzmrAAO+mnWeZHiaMaBS1+EWNXTfzHnKcnDYjiCY6MRoKci5SDZk+nhiznXBw7MVm
KbSI20d2U0R0QcL2rlYMDP7chEpTUdDbbojAi8op1XjAdPhvEl/N2qcEt6022tDo8FzPZzBoh6tP
BxeNiXitlhHxG1IB6BRiAHzBMYOy++0HNnSSgHsqi1oyWNnUQl5ZpOtUpvPbafrXBLJdAGW1We4n
zGT5vfIk5IqZQkBI8GiA8lGbuawvPQpdU7iSxmPM/J3TIig/ysPfESy88+4CTiAwH6kivkckoduj
0Vx/dBOyRcoyBqvBkRUbmGiDp2l+Rgxs7s7bnuB9aoHsD8P3Mse1y6TwjKHdk2Qh3k9fbX4G6UuL
bj9jUiB3GyQvuVWV0FUgeDUNrpbHEfjZ1aeTLJ7qGyEwRIpbaRysfdCG4/tCnFL33s+prDv/6wBY
Ibeh8p7VL1oJ8Azz8uALice3B0pp4kgNE/E+yW4T9PEKeCU0Vzjhyg+nC+LWwXZldskKuaVRvu5m
ApVTQHcBN0IkOlIk+hYO0AhJYPh1UECZaqRSGZP7DHbVuWe9gvR5N1onrwloaX+js6HfDbo4c+bU
xpVwTcocJmjNDs52Yj7vhMZA1JOvA+mqkbKuGJtv87izUgk7gqTg8U+SS5i3LfE/2plw6S9wPesa
k6pQjwoKIUADPPfRSlePsmdqfueRWtwZiZamZregExMIh12EIGCiVxN0u26nOfnqLWIfvf36eb0v
AApGTCkDPmwMiSoz/Sw5j3FR5msyWqxT5o7D7C6QemXC0EofX2R9CYbDEcTRk93j7KwqpeaWvjrU
+A2uJ2kGoz2oNx6cukjWXhhTIJ8hULrpDgAEsDQYoyrV7l+vpT8/y61Xx715oemgsPb539ZsMgYU
zAbUbd2lBh8VwS0PMW3RshmTBAkgEr5BtuoKbs0xCKJ3Fc3X3s8MJhBvPzBzwaKN74kWnnjOoxex
of1cZyJAnbo0ijfazoLHvQHeddJVSjJ5WlLWPsNxRC6kNsik9rluQP7QjrLYwEp0ek5KVy9Ia2UT
Zt9XlGGeiLh2kwhBApkkKxVgZF0XXQU3dVkQ1p1Wpx5TAz9NohEBfKZ/1mv9PnPlQVFSuxWCKBlw
8pHqPjf4OXWtORWWdiNy/Q5xsJDcxaamXC3I3ufvEkaeWPoTW4ABMiHn5sUt5vDhJTHf4jVGagql
l9Ko3JopHjBggII8xQ9nRXBo8LPivz8yHJ3vyfhlxZ16jPlUuJIyj2jztfPdO1xCfoWkfGB3X43z
72bEkX55qgra1vv6knc7j6L+j/3uLNlu4dOAFh3CUvnRdzSH1/JK3xbo7/dzAVST3cYeTe47An2N
Pv/IySecQY/Vt38XWTjLdYF4J87QsHXfm2Vi2OeiKgLzKf3EnsZyZLYoE4E/o0mq5itqP7P5hw/k
J/TOo6YzNV6hVdqk9B+XeHDUuhPZ7scKAqSdIIgjTHCYJVBlIm19vJ2jHhju6P9FJtn11SfJu9rr
O2rzKf0ybB0IgdDfRhsOBQyjKFHdN1Y+LX5gg8+P7B7Ar++skE2/RdDBDtyOnoZBNdna3lf3K50i
xNOsnUtCWdMgjq6JokyJEhPQX7sHcdCtHaYL4Gc6Mz1RwlxBJ8fKCpYtubLU4HmaZ3YDZ7qH/+nF
2JyL1rRFaEKSRC7YlhefiZhw0o9LIZvJDbG6GOweaDeUJVFppiQXN2OtRMiwBr6y1TkdoMsE8dO2
8ZxCxlyILO8/9p+3cph62xSSjAJIaaRMNq/JpLBiqrecwBXwvyMyK05Wwf+8/MotbLtWKY1i/+an
EuHDA28aQ8F3ScdgG5P084UzqCkcd1wHSoM5AmmK1NcD+EQW09zPf5GESGk8joyD8mx0IRQbzJzp
etgeW8W022aHs6i4gTX4psGxgT6CE/RG7Ir1IOp4k0yvGuPRfumndX7C0JdQf8L2uQHUN+zeYcOl
I2h4r8Y2iTSUuV5Vv9UyB5k7IML843yMuiehbczK0BfZ+VGpq8sARkGRmIkfOqsO54hT+oAFb577
5hdChoI31ugo0LwxhU1pSGKv3qGQJzp1uRotRhDpa+cyMF9kswjqIdrLPW1nfGKSUxQpDo1OL+C2
a0u1VVi/xX5v9zFMg/cpwT/3hTV2kM9iZw+pWBI93BrinCBdaQx9SAc1ibd2D1Lo0i2ctoLDj9fN
3usih9BACSp1hoGv2i9ASlocGSYfo8vDJ3opcDZUq9PoaZIihP2aq0Be0gsgRcx5w5yvrC5fY/3b
N1g1m3sRt/X+WL9O8BKwUZfdAjpBr/4zc2NVoIdjeF7X0Wki5fVwxqvxM3dYaxkUDpKYnV0NG50O
yHGfhu6dawULyW38rgL4NIvc0TNhHfkasr8K7vJIywl9dGoxI/ungSnqWNQatwgyoWkE6Dhh9nwu
eSUvqIY4BcVos6bHNAdgFztQHVtNEL0TkDleJADRXmTDJ1BrdbGUvrdXSWCWv62wL4jKZXx6bpBg
P++XYvKwbykZiLgklKIe2ckb4dU2J1s5KEKF/8youmXbkNH1kjQUqAFPqS9oJRJV/g2KdbNH94oy
RlyJLL/I1TmCX156OBpPXXLL07ASrdnt/EV3mmI0gpp7AiuYTTV5WhEfUaus3BoY8TvhCpflCeb/
7zhROlBuXLwmjPUOX0Me1ZMDVUnDMbDLstcKoGPJS+KfRyBZwe3az6loCOTyrgJxkmsZLLUZijgd
8GqVfNepnt2aJ6Om1KA2SIXjkEFcQrvbh9wbOopJ9G1Ddn07C71i3zkijenkazQK2atqBy3iHwd7
4syq3mCzCQXLZedBbP7WQ3Y39dl26Gfl1TB0wilox/5nuYk3TPJ/Yfpk+5qppjVNUO414RMOyLPh
6lJfIhll9oGbczdYqVXfBZq0ToYKst8cYi3VRyzwgXl3KsAqBcVG2bH1JjrDJK6Y6HyXD1KaJbgl
poMT4GJiA2LvQZ9nLYYjE+ApAbeZt5q3RjWbouSo6wFgb3CeTjkpdWqjYc8mKa0JTqabCVm/giPR
5Rxb/oF51EN4WKtlJHx4LkLkiV7OvhkfWO6NNEcGr8LliMJl74AUnamGiNfL82Sl5Tl8P6gn/cIn
BK50ynQGy8q661/q/QGWi6xtfrhHmT5sXGvjJ6Ou/R/1wf/aiP+sa7F5cruJVDvuUQe6xLgUEm0k
fgZHdLacY935L1V14Er4TpXh518ePz1v/SvH5yBfsNGTnMRgx4ErvMSd2k8/lZ0b73kZPIjJn7Kt
7pLRuR5dC689w73/IM4/mxZYAc9zydfRvBmasCnFCdmXT+bzm43lQEUC34BQ+fTP6kIdSxJx+7Wm
+4dOOj0e9HPTvsx+vPJ562yTXi8EP2UBO6J6557nfe7gyxNkt+eieds2FsLBeMJz63yRQcJlHjrh
yzMOs5Hxl3maulR7o/ZuzAa2BO9Q7au2elcxPHpL97O6CQ0mH33yMq/uYr1xdcUQj0ep2y3Nexfh
Xu8D1zqUDFj08EfxsIC4MeZiQdOzIE+SdJh/mRu6NtqX1oHqtUEUCi7+RUs8GWQQ0UvOVxrQ/tCM
FEpn22yA6+74DRm+KDoSZfwvnWJkcKN3ES2c3MUi5UP7bfGhNjNiNEAxLWit0/h2BWiPWzFSyZeO
eU/y3SOpowkp1/6NPElGc9Og0fMX7J2J1HvTVE0f6TzGG6Sk+b+ZkLmFgEwP06GBKgV38qt8INcU
gmWquEGa4ZGtUMjfTGGKCHNkoQWiwx9PNVn2w0cHRczQQsbbSERZrjBXzurhrmlP5t5jfHDrZmoF
c1hZrKjVd+6sY9vdoIkFY/CrgGBMUyRGxM/tO0lbQlQ2BDhikvmNUw2pKvE7w5v/pEIGmk8f8fGt
AJmbe3ZpkmgCVMde8kDfnM8LivAhoy/dzJgl34CFw8P0zRMOgxhR/Yjr8zcxP6TmvooPFSb20Hli
Di8ikNu5AXGZhLH6nGTOjM12paZCNLiv9dNLc8VQTRcjQ7qyHA1sG9PhqTmHxixya/NkAVni2KNN
I3Mqxli7EsrsST/9SwDWiKjMAG9iBtG7DALENtMga9Ajeg6bbFMs1IyklXockztcsvzLmagfrFtj
615WCcSTZVb8/vji4EdxACI2jg/xLK9FED17yxaJgF1pyDjehe0mUeS6NWt+7BgxBIIsk27Plo/H
q/IvWRTAESyYIr/pGBaOIqU7r13P8wp8lMCiObWFChSHiRtMysFQf3C+bS0V6gLH8SYQNbDZYwGr
NC72WflsRJB7mzWd/RilvtZ00WbYnaZj/2+kyHjP11ULv0Ky4VvM2uPBGPsK+pcWelGJlT8SCED5
3FFSx37ZLDSOdvYSXLRrqqYfVt22tl/XEEEdVyWAlBWlSRoTiF3CNILHtNQOhvTJamXHdb0MbIOw
i+Ae/rIYF9/5JaGBLHGb1cEHQttEUlTxmGgb/WfPPe1Q4h8YRYuCfXx+sQHnGUAmktomUJLqAlMx
7shUQLrytYEKLdtwV9yV5+P52XrNOmfe+iAUmq1YU/UyPg46PIVdlveOuLmfQgFdpr0qYMkXN2w5
Z6qeN+6Lrh2KRZTvvyDEec/wZgnSiDf0gjMd0xT62+uds5JBvVN16KDrOHBLFmvSL8XWgSNOX0+O
wrWb50KQFI3YXxEJlerusFi9UHPof6VdlfI00sG07f4tYqfz9IQH8jIMVcXLShjNSUzLKMEWZU66
E0l3XQwbsxj4hWFEKM7E4Vg6kJpQxwEAkGQGIcMN1+MMZCGvrFrC4yxljrIgCRdcJC5NwcCavQWb
I70mcVP9vL2mozHo83R3c6HQZVRkitEm9df5bW4bMpNqctCjLBqdquiGkLQSAlaqqlTWnlKEfMMs
W8JNuKiFek4Ahr57Q66yTugbz2WB+fGn7GDz3hMChh+hNkqV1HsHHhtDu/hyP3iMb/nxWAGA55L6
CDeE7/88W1gNCFWiE85KhgdXPeJFeCSUA9wqHviZOtLv7nfwatWNRdgietraJNRwxWRhVzvqsyOy
uM4zPNGsijMYKW2IoCa/YtuVBCEIEMfwQKZ9G4G4Hy/+jzKyVb13IIm+0Cf2FlhcezwlMQIReW4J
B0lFMOTa+aZyC5lFU0P9IGt/NpLaQ3QsD3Xc0NsaCb2NGwBbBnnmi3DYGMDsGoJMCOMKJAsPUqFV
izGX3MYt05aHIfY1gy0nP5le2wHnitMQLN8MQWA2xejusuTK9/ytXm0G9pqrP/MSzfvsGJQ7vGzn
d4wo64TW1Qe0Sw61WVsVrCZRj2mtOEzR8tjjSiCxKGm2saCPptb1eOkDGA55yXs3fn+wQccSzfA3
kyBL+fvBuzf3EGil6XGAG6c80EMOoUv9tErFDrf4qAj2o9oLhp7AGhYVV5JsW4lweWi/AeUd0npH
ZLdXkg6pouykQsne+w1NJ4HcbSpBg+r4F1PoqIV9FrQfWWEcOAgPqY22mmQ6cr2I9j/X/GElk0Uz
YAsbNDGTRSSINDa4Oi/hBNoVpiH3tCjkTZKQens1RDZf1t4FMsIvAPFGXKqGzIXu8wpvnuU9lCAC
2UCh/3X2VK91CnqqPqOVzCeE5EcJOhn4ehNWDJIHJsIPf1PTeRSkZNs0egz2YVk+TDPjTUhsvNNN
PJM6UTgCAtnqg3fgpgsOPFgUnzDKMZXdKuJlPgxH87TcOrCS4vnWBy0mz3zZxcMacnTV9x2PoI3x
m3nkgwQlQpIt4DZbFJnPk7Uvb8M5n7SyMeQZGwcUgEywxSkznwpS40QyUxupfO9bQNyLNtO3LXhT
HrGLiblrMxxzdjPzyKGIUzx2frf/zQQicWOVHVCcaTw/s8raYYqmqY2263qp1RXSgAJyBRGjEnkb
y/08yxmcECrbOgklbgwQbUtb/Ioz4QAVDNKgT5slAb31XfPcvVFN8X+/l7sQ+OZtEYciPgqrODZY
TAkWUinpj5iIxcgGmgq1ITrSqnxrUunr/mxbr/5CjUK1KkyuHZIryhJJi8r9zkx82pHnoC2+MkHP
P0H5cVFXw5MF2Bmy+qvh5+aZenPKGHjCgJmg3EKwBKzskaz7GsiZGqpDiDhuQukkezQNzP/4KQoA
IV37/+Fs6WKx1KqRQ2w4af7OmAUjWt7pOaekNs0+1mMrHvKR9tNXyZNumg0xVhWFfwIVJBey0vrv
ZrC3nvgRhq+3yMDaJ0NleFhIbIRnLgrB3M01ULINhyN5q0n2oHbDJ163WmNI97Z/TdYns4dytfh6
PhLzO9eUbQoSfO78MbmClmd2NLFX9/xVL09cKF7A9eh8FWSGRqPkMdl05DDbGM4OTQ7YnxAduvs2
xXO/Y3YLRN4fXjxQvNO2VeQ1ybLzzsThwKiHXamVeW8J2EQR2FNEkb548EFzvsFMIB85tM8TRpf6
wXwC6cksnmlruxTveZdauKcGqK9Ji6fLTM/+oAh1Z3RIMncreVpXZCrkyYUD7FMOwJB59NOD9n+1
mubCQ1Ip88ERZ04aE2GJCV7ZFh0rXfo8zvSEmhQ10J3+lAq4HQzRpCm0wFtoOL8Vt3QUPXBPm10W
ep5CWG5PUJ3G1tBcI61MRgexaJI9vXsGUASqMA/xhYO1GqziTbElT1urJT1p4y3ChPhT8cqpxZls
S5zueliFgPApd/c+5Uzrw8eiTvnopzEM+HiZKobyXlPb/Z2/Wqt24U+UWTdP2w0zwgAxtleb5/Zn
CofaXfa+Vy1leycJ0FM+qsd76VE3g6NoNF4AM/Me5L+dpU0ndzlSne4izKfHGB/jy7Inavkd1WzX
RzEuUBk9InQZHTJLlqMpQGndlmhnLeTNzYIuXzOA1H3cxYDmzOChx8dZsr8qrGnmUQqXRVMcjkA+
6v2nhOC2wufJZKbwrQA+AVk/DJwklSsxLizrPFE7b1zVccKKlaiLAuUsTFD5vjnL+3EsQRE5TXX/
mhFd2y6Fa8W2bHkDWYq/M+Y1LD17HWATR5+iLKcd0FKQ71Eg/Fgjc2Y1cDcJQB5HV9Slsc+46pT3
q4OD/VHuN+PJQF6kPB5sfONUWGLoCGW/7kWOpcQsWp0agbcytzKzmWbqyjluVQ2rT3nK+wzqbKNl
7GhOj9cENOcST/+TyftVL/a6AtZdwllX7IucEX1E5TQqdNTGEQ3RJ7NQx7ghJvTqw6pHd+FZ5Pbe
tJ41Y86GItZaYnnLWtaQVqP3nre4W7gETKHFEhbjE1x5/QkvWDH0k95N9vZw1u8f+Mi7v25R8M8V
KY5d0zdiKuxmubH28IzyuTT4mGlxqCxXddnwuYIrMo6VR0i0n1u/54i8ooAIyVOHc3NyJGYjPC1Q
U7APsV89/BuWNslpSRgFzqMnnfXVJ3U11g0OsareGkLn9FFN4/M+j+HWYf1dn+eqHDsKJD5oPiDX
eiLHHY9Ktv+34j431VAI4JYUGeMqZGe7wGjBwkMoc2KsH2G2O0pQmxp8bYrtykb+bhVJlQBx/2+m
BaeFwHfo363xYkljTJ+uUp2U/ibNrP26cfPJfcvIFYx635wOq3Mwt9QmhKHBqI/JiUfrdt5na1+y
2sEevO4dDLGKZ6ekTnhg7Ahe6pjl+Vz9LKujZlgwLxvXRNSqGYJlcmFLq/HG699clThqWYmxVVq1
zTvUi+C80UY6TJHHyEd+K1LjfWAfX4MiSIMWs8Yq4l9ofdBDobVx+GaF4926V9BWNJHUFB2js+fb
vlDVmz4IOtWFvH0JLWRbpjJAFonIscqosFTWzZ/8TUwrjO9cLtlAzS6Bvcw1TP1NYDylE5WJeNXg
xrEhSsshOpNWqTNbXcD0S4sWoDaq7c3UXshXXjNW2W/ASXJYvnYoeuZhqhaMAj0SAU2gYZZYN1SM
2ABMOKOhcebLXHnaRBh0tAmV7I2AH7lhgj/2V57elgkjIiuGaDIsPY7LO9Sq/filecvat9CF+w1k
Gl9pCZKlahxvyiI+z1qqcQFGqB/p6VS3hlGylvEsxM6Ki21BwSd/2AufBXO217/IimHhvIrnKyeM
WIisxVvSLsOVcmByq7am1QaBMk8qJ1U2++V3y3wv0+lCuaPxmTVdm14z2GGOvrhKTrX4D4n5k7Zw
nvTorsp4PjmkM4ix6keKMhuUpWm4En0SKkOr3BsdijmpIlG/nb0x5tcDGNirjtok90vyu+9sPs9S
cd24Tv/uEkxRgv8otHJHimDJiSpCwE8xYstsRm4ETcRj98fbBIRgMmyy+CNwE96JCDGO7mkLWFuj
cSU8zpcB0Lj3qi9oyR3xHGRVLKOJxY379H6780Lm8YLLlBKH/jVHQzURZZghjB+h2Ba9gfVqWINq
f7X4j6hiGelWjnJT+ybhD+zz1OUR2T9AFRHnnKnaCRhAjVkAwLnOTHqCuf3GSYtB9PUc8ZQm9N65
2vuavnFdyvWqKl4SGDmFe/uwOYDBBEhVkFdKJhGDUP22vWH4zeyyLZD/kNuWjN9MhqCT0RZYyVLQ
30RCOUJ3FY7eAxF/rH36t2SIo9AlfuqRbHmpy6Lze7cwztPziBQrcWGD0sRje9wlX7KDkYSQIzZX
6bX7A0j4NJktBQowJ2ushCDgrACqacYNKZFUve9xeHOMmQwLdwqSoo08V0UrzJr/IvMPVFWRBRWF
IuVTYalUKRnWbvDeK56xN0JyPn21r+jGFKQcYO5Ab6uVpa7p3AvatEidU5yqVO26BMMgnovn1DaU
i+s0gzIe2ynR5A7Vi0vJlzWrPby2y/66QymwPBIvQ45iiW7NTpP456Ku+D+h1GXq9MUZo2wD89wL
9f6Eyuh+wWoxujVqFmTa2/L+YFFVhmw0KmBUzapvJUDc4bXlqGXPf9i8mPW2ztb4RiJaGbXYzAay
ptyArf36KeNcJyIItRAvIswvu08XPQg4VtAtDC4E0OVjrrdkiQoRYFnKMECLPRRbAezGMoStrE9R
stYfeeiGmHZZASisLbUxYo/qncQm0qqdP00MxjEm14Kj3PuB7hNvo2QyikvLqYcgenJUdNh5ROgi
4evAPwMFHY+HKjVTPmbK4jvNfxSICzUo7DeSJBzkdaeg28KB01s71Ypxt2m0zRJu4I7nThjONgZy
UF5hUChdMuY2UQjEVzDaofmqO6EQsJJTHKBmjkXuOEqQCk5JcbvP7+52rMOuS0ysNUJjmM7YrjT9
VTmFfC/Fzn4MJ9IzezFXLUugrkM4siNFGMzKbBBTiRwOcN7vUPhEWsjPiIn0O2vofnkGGH54ikS2
to7F3WEAnf8ZekFSboeCHZK2Qr+iw//94ciEEPnjWj42UgaWA53GNZtlKyxfBUT4OFsjfCAM4DyH
kVtfRX1LS28YJ9jUTpjRsMoo+Ykz+VLSUcvPtl+FioJZ9ixk0ovFi0Ytdsot8OOduPItdku6U3rI
fGNW7DyNi/8sln0koj1SFrgVqcJGABQhysFDNVQlotDgb83qp63DRwvNH7oSQmuLB+TqsKvprp+5
0GvVtDLhyG6J7h0lUb0ZpRrHW+LSje0lbGFNail7iNHRzEs0ugcVUGnSwB40BnJXuzURz9mRSNqu
sJZBB/gHnRTI8rkPLs7ZjFbQ/HPUTiM0oCsGQz96p0rY78byKrinncp5F8cuohGyiiYwJkkz9/Uj
43/pe1W534T01Gr27HV9B91eO24ISGCkQJJhcoJBf0hlczWbnNiTW4JgzHZqZBydOVZ/e6V0RhDh
Bou0AxFE3FMWs/7RAmrDKU+sfV0mK2xf65xJwBMIfZZNbj92D9ZXNX/anYQanreFyUBORa2HQuJv
8BfPXbt7nOyu56iEG8UQcL4JwO20swrV1lfvXWNvlwwrdlMHiuMtCp0aO5lWwPeWwMyfjXFpmKL5
73OQBmPkaw6zzvWZGjizWsONH/sb/TR2+K5k3bBTEngg5TFHyofIJhMbgbkPWRsXZB34/MevkYv4
G8KvqRH3h1QfOCYe2ihaAQfJeCI49EDSYUxuKcucplqj8sOxzRfFXMX7XjrM9DtJpIKya+Fz1tns
t/jawtO649mjwOasGFLMhJ3QoKI8WLLLJ5pbtmtbDaZUappmAZoRF7gFqBzhkwzlcd0V47VfzeQE
rqZQ9yg5xGyYvaSOn5vNkATICcmcD9iAJ3/tcBjyIjy92AN+RPduEht//xKk5rBpNxdl4nYaWrsC
vkJml1aMICkqUoK2grWoj7nW+kKlMkMerp9mnmRnlv3FjyRJZkCbxJEpmdSHxKIiTB41bGOScOW7
gJxoQPklQvYgwf8Fmn7K/vM9TuHPqsUxrQCAtR/lZWdXUJnRvTfdXDx01pm6p8OR1c25XoWoDcJz
MXAxUf01UhXXti9WU7DGfpnW54D/wxEilqCcCTMDjy+20Agl0GU6aI20UkYDRbKnACwDE2j+gtt4
6+M4ZC0c5ef6nmfc7ob8IBr5CZXN9ymLEhcXS43MQ9o81EiFjEI6m0AEkuYWGsL4ykROvSlY5bSX
HH7BewIAa5AOVsx1FnEsVACnY7cLheyu+fSXZ0xEauPBeYPCebaEN5oI0WH8Zy/qBJIkrJFc/dP0
fDpNc6Xjn/m9WNwcpIMtcdtjkY/5pAVrwk0zLt1ooyxSIOkkSvXUY/VKRiHXalwK6S3zzj4cmzZL
vcpcRfNKUCWFRtmPHNmDWVz5a6E8+bCdX2LkW4CYgUDxzhmmOOOuDF4s8pwhcTV9sH+/jHE0hQY2
YVnxFtQ0N8n+UoPAegjBxE1YV3dm1Q14dgcqWuM3d5TJ6qcRbs+Pxh0FN8bJaRjqdAXmwgIGCrco
ekUbr+HzxQvgXCorZWfOaid5qKspO3YYRRIGm7e96ccDwopznHF1qiQpaXAo/CR6rm+GRVPUzH/K
7xEv2tNt7yBOuKZClKEjkFPF0gWC6Eksqzy30Kqc9RHjohwOCiFTXpznq5DoT2BcmMVtApq2G+TV
qvapFV5PuRVriw5FRzOJmouQJbFM7vf1H90h4pr5MmrFpqbYb0gGBwWX76CGHoYqr5COf6GDEbPM
9vykMqpOoCrxju3BqtTXqxQjpYXFtuNSFD/SlpVI+9IHq6nfTsYYaAlJrX+eSEauWmro/FbBkK7W
HwZZXMFgkjLhHwrnAm+9BYmLUhZrO4/mm5r41byMZWRhHD8juR1K/mz7LWxBrkrBwUAh2sNP1oNI
EjB06K9puvqgCGstR5TQfct1vHCM6ityhqXqlnHRbFvO/WjF2nBE86uWhrTtvSh1Cc0gOBiBZFOT
pOmPDrtXRZyi+XKkl7IEgQfrx0xnmsVBR0my+hyI4Wili7wIucC8JqfyuoNmga0w+S1bw2YojyCE
evc82mPOvX6n+6as8kgDUzPfyxHkeyeK+iFocuKTRl7lVayfbX0M4IIrcWVXAWxTVXeUyfOtVOx9
myVzpdwwu1VghBJwVy8ZMGtWy0UyQoM2MNJlxSWva9AgITfj21FGEpCWrdrlSTnUQFsV6C2uLpHL
Gu07P1jUcQEaHRI9VLq6VHV2b36csIduI59xQFhFGjitvEFYSYmrG+QS24/lH4IjT2w32fD0UEIE
owi3myo9ip1HulWXTpwe3iXBpo6//ka3+zvM2xpBKY5i8DCJo+CfaPN/Zmf//K+jLeMwWhtKnyGG
+5IkdS0cqRAKOH6zi7m9BE6BNts7kvB6UPYy+h7J9lh82jFkbk0mhGGjM2nO5u8Pf2Fmxc+zNqNA
A1KbbTrZCsKJhgKZ/ej2VKjg4B6b5JHFlFj/jlrL9z+JKM/5/LKOoqRdb130iSK/ff9QvIDVurUF
tI4T7WI19x5Yt88vu65eK3vibA4odVQXL7U3FebIZ5MY3eVgX4BbyHG4VFM5Yfw6q/kxic4vLMPB
DgFdV61wRp5xb/KywojSChgPpyamEUmpsyX/BIM2ZVCXrr8XrPYG5v+6vPWaI42bHXprHVKMLqkN
4M0RqOWMX9xa2oiblb4EpG2wbaf5llX5sbZxq6uJBzdepA5vc+FNL6Ut4NEjzJ9RB5V/Fx/+6Qyf
xpcvBXzNcsZ10a+z2wCwiRSPNeUL5JD+bvqbLXtsTVnZjkXNWMoI+SyU9/aZjc/KvmgpgP7hSP5r
NjmZpHl7MMGB3xBrbZeSfEbclsaG5Np7sxpuKvhU1XbnGFi6D0Id9dS6N5ImRpb0s9ZngX9wPoxS
FEiMrDks59HyF4ZPd3T/DseUwY2xSHlHi3mMHAN69gdVO8IuXGk6uGOWwFjpr5WIH+axJO7v/L6k
b48VFKqkd0ijUSc7hzfKiBVXaPF9vvph/hvvgTQHtQO2hXM037ADfelCIjfT24dqNtE7V1VaNNif
OR4Qp1kbQoEibIvWwWi7f5s4RIpwXfTlOCaRUtQ3dGTZjFVNMBlcG+742u7l+FY7Q1jhmQLCBA2P
Y6n3GdfbvGOlEa06zrLTypBUcY7Xu2wEi+x4e3KW8ATTkv1xJVMH4BWSbLHX/pUnLtoBzWFgs3l8
QspEAP8Ihq6ct+mVEo4pShgji/N9xyZYZDxdIxEshPH79nhTHQO0J6vpj8RMxjGWocYsg0PO1Goq
xr9R8/KHlvCgxy7h0TnDmC1XiQUAwKPIWejQDwid7vg3yWcxObvztQO9pVyalFmgd86jjp05Kbhn
8gBKTKx1OjnU3Zs7tmGcPjXKNMH9uKpoittICiWotjwzqs7Xa5dbX/p+88JddACG0d1t16KgKi9a
ZyX7q9p6y5250kvfL4G0xBMviuqjdtohdCppudiZQncLlP4oP+ZpQysV8UAUKwjjXpb6tEgiMd+u
8EvAW+Pe9/p+bPA43brd0X+6GYbztuslCC2rc/HWRLW1w/VQvmAJaszZMR8UpLPtVBVp2DDnkiJ1
EwFG3nkq5+V2C90/BOnzUS3otvtyoLh96QHwFLev7c/DePbzMixpBE4xSScF72sIosEKlZBluABZ
L7eKsM3FS8V2nVYBXUXkGSr8JIYp2zYLP//YcO6iiqyT1HvURKJ/IZjkyF8TwKqCm3kRHCaUkJEn
4NRwp+HM79G/Y1KQtG57o1sFW0SnOC8GMkBe3ewUk9sJw098I75MVyezNMZMd+kBt4q73PtnMQtR
3KycSCP5XWYsrGBA/zaFV8vho0TfZX1Al5Gd+d8r1gDSyZ+EXRJgmjnMFaz8z07GMgtfZMGFSwMU
rDYgiI8LjLtAHNOCmP0iAoIdms0CmiYGdWDQrK3PQde4h9PgcVm2VsiR7upIydJZg/UbZlfluFvq
dNpjvkzJFGcepypfSBPgp89z8S8AFdzhBQRznN3kc/hqMacaDwqUSN17Ktvqb9m3LpVhoyf8V+Km
Dp3bCc6eyTs2gNiyatVD0cCZrLlkZdu3opD+gA6FYb/sJLo1Xko1L7S9ts9ktexnwDoYONnYyDEK
NEDmnd7wboPUFsFIL6nLWxIM0rhjB2LFz3Go03hRdxpj0tyOjTLvm6qTW5rNp9yPpKDhRvy/6KPi
2Yaqmu7+x6yhkaeyrdDwq7cbDT8UZ77SYUsn+39DjYrThntHYUGjmiDzGp7+C2lt5Fl4SK8EtYZy
EMetd/EfD7n5O5ttfo581vmTMzfNInzhSBGnNTmrcyw1N6cSfWOF25O6JbI/VfZlHxE9HMdxQbeT
cogFSn29OKZNtFwknxN6V8+hyVRkMLR4O0JJgvUu/vQER9PI25ZFy8GBhtYIMG7Sz5ielNAEnb2M
D8pqfAjuqV2Ux36IrzGjiFIVJepNN2jwfksIH8y++ItwBziFTsWH1o4z+zSxP+jw5KSKN5NYMV70
lVjXiUudANiJ9rcb3J9gNKGGyJ+qSRog4QCnhexax353PWt2d7YZT24t/b30fSMdvMNcm4Vzbuy+
A09YH3MWvz7b+FPHwyaeKFrA75/lw04JHPUn6KMwllHiksMIdEFuy/CKc4vdO9fG72uyMyiquNBS
60j1x8z8e3AkmmO9+Lu9JMZjeli3SGNGs3PwXn/zA1O3cFHcG+yaAoskrqfFnuopNqT6sjPwqU0U
kyBSGv682phUuKt0dZdq/BizOk5Dwzr2CUHDksmjE+O/vg7NBY7KWYsXEF0F1u4MNCF2yP63zVSJ
bPT34BdrJCAfZwI32EKmExgzSI33SKAYHRgwV0WZJNyjYbW15o/A+gYDB7yu9BDdgWvGJxYP2zQF
QpPAuHdo13wo1F9YGJpiTbg7UJnn9bpxcMpKLXkIqdFYgi3TATfYVG7G+jbu+YMeB6QQEK5EjFU+
vDx2BJhrnnp5K38umRkZJ4ahWmpGv9gkj060ASuKL0wVGOxS2oNlLdppQIcpBJ+xtgkvRRs7VB+Y
lfWn6myRCAUnzE4vL8aMIbWdWBUlLV/A51n+CI9f8DDYI9ywu09Oy589MauCp6Snolj6sYMCET0s
8BxxQzXiFSRaewDXw1J4nM3nVkFAcODsNxAh4Cw25lGrrcrae9uxA2yO/AhH39Hbg2Ph0ifJ0rLv
+O7R+4BE8+ZgPmAJXr4omjB5Df6FH5K6iDjB6q/htYjHn7EqETI3t/228ju9GUNsc6ZgMe1+2s+W
01awk7v6U3MCWPCVpFDw8CrcljxM+VDFIpBG9ZoJKOQk/fiw7maNPsoDF7q9NQN89VJfUvOWCq7g
vPCRnEXTDh8VGoAJcp3OM5Zk0v210Mq3kcHl8FZ1ELamx+d3/x42iz3wfPjeqbiNkUMn7HOHIBXf
pRR5Fvs4Hm4PTnxlwwHqaiPLA/UfPpHGFv8IOi07t5uDZTBHTIDcIp7CoAkTfoSa/yHe5M1aY2ni
rjo53BxTcKNgdpbJnqVomTeiPFmS5cmemfCL+KLDZhtlprhMqrdGEvpzVDQzvBEROpt+YVbnxPwz
9cuC1d4QVzWcaFnXcq1TOO0kPTsBosRUgcFCl5XA6UKERcoR7TZLluMGtjbXl7GBcBrAwoOdvOqZ
05tbi8/8NQ5sMFYHkesBuDa26ImkoTrXC+uVuIXABwRUUnFaMC5nBdhn9CBnDed+AVM6i4nvBgv1
dFFGFCwt+9W93WR8Szgc114SIKKHWeY97NBNKO5m8cSlUU4zjd8ZV3pCF4heb6cPRodkQH/P/ckY
Pdc8F4yDNOvdYNlZ5kDfLcOHIPZkmIWBM6DmfNLim4uefaVyaO2HwTTlctMvBm81POQ1Ox5jvXzE
GwXLedgKUg667g054q18us6UgHn0wsbkR8gE6kN26m6u3hc1VTX+Nc2/nGljwdogZsG33vscCYDR
OoaCT4pU41AaLjnRaDdiOcmN+mufn5bXJzJIFYhVXW+7A+NPjXHsXvQrIs3Hh5rTyV09raPHfPpR
iiXaswgOVug4l12uDpocFIZI3HUiehzBwcVG4shfUkCVgHPOn2xoFx6Ce09uouGY86Mio3ViCTmV
ck9EL3KNxi7evjmFesJaJJVlm5hO72qiLunwC4mpXTt6T8Sdo8gTTZkwLrukJxmUE5tv8lPY1xp5
oT6UgPYEZSmmW+Osfo4WHLiqbY1p13lKkGFC07/cz9AFzfQRb6MhKo5YJgRzQqi2nBkOwmCnYTOv
TN93/sHc3r8Qgk5VQrTfIZnzCaOmQVQKVpMmU9IMKhsCWrpl+GPfdHnnOW3ZGqNvHNNykhmX0BRo
bYVhAP6j0M2IN4se85I49htX3Pt6lIPEYPa9N1Y1nQIgzrsrQToDKtirEhBg8nPyzyRJvdxesDSr
gfoYtGi3Uf4veKpBfu516hQERB/Z7DFBF2NBshVAAhBe2qzaudIJ/byS8SbXd4Bcpw2WzX0QeZbY
IdpMOK8D0sw6uJFshsquO+aQa9xM+UnWBtKRr91YMcIxgAWmqpLlolNLfd61Jjg45f0gCo46xhWC
K3fxWR4s09Yk+uXXiiH+FkamknIij1eBulZUzR0YT+e1W5fAeGEMtUKwI2BMLXmR7l3DMiOlnxSS
XUv7Ll1//anyQcxLhpqYoP7uvBelN+hFSeMvtnll4BZ3SsrtIGkVUGVWFGwe1t0WFJvKyldpUQem
uMWSkbpZ9yQ9mjyFBKZCHf7QalVJuNjb/c4Lioy3zILk2jJgP+pThsopZX9RWA8WSDrjRvKGXwYq
N6DQFsXylG9JAG6z8e/fp2RJNk4WIqCUSg65803KTjAaOM2of+S/j0ZVssdj+tQgG0dfd3HmbrXW
Ba2XUFAnU5ZeeFoBq3xVnUS7JzKFwIDNiuV7t86nvvGq2mPq6RzJxGGbJwfDecntijM9oKypGXwy
1wubE2J9GsijRM96g/EkPS6nYTzxEW2+tJrzA2QMMYPVhT6HUPnyT8vwuE3nud5VL0e/PHW0UAdo
Oyj34hXxObNgcnznjM47OZfvMqzK8d81+tYsGgNJAReJAipCcIarn99K5Me/FafUG5FD4eo0l5F9
10lwNajmIrvhTik0wNbzRDUFTl5HbafzisvQ5zzMoLesr2JGi8CJAkf4uO8j9NcNx2jZiZVSQ3tw
TbI5ELYCiu33uYciEznR3B0cB8mFIFDBkNoP+ZpxggU22C5U/UUDZOmFGwDtdCGhT9A8YY8RqMuD
BUxmRLQq/e8UVs/Hfab5Ur0wuc70PjA3PTG1+PZRcDP1Zvkc10TYIv3kQWi4x3uCFzK1N7J7+Gn0
D8HWKtuyKOlf1rzqI+Co+J2QqVN91UJ/EjHU7ekJkyAvYTsSlk0jR65nqMYgE/c9w4J6Xzus0/fU
ZzHT42ZratVHF0/wcHOuqJnp2bDwtR39OIT/gNTJ6A7yZZnlr7HeE5x+cvHJoXKWjAX1QlmKhk13
pMENNCRqQe/YchTN5oCp4X4r3EA6zgrFeaZyJg775S9b2C5c/iTvg9Xebt/qvo0SJWsaCGXa9FEn
hTaNXZKv95rKc5E74EK/p8JpHuoYFNA5aqDc6haKQEbwt4RcIIyUMAwKHITI3Bx8H7fuOGO/jmdA
HQUiE87VVzjY3A1pHnZPh48IkfASyqwA58UKqrI4LYiQgIP+v2dC5+YR3yG54fRf/5qHOqcvJy7b
CxTS6LBWOobY8gRbQITfj19xrMm1Qj/8cMbrDX787xOL24uHV1570urvQaststmMxakXrBQgZnlV
SyJ0PJ7c3rrDvMiWlGpZikTcvVoVDFEHR6w2jzA5LP5GMzQpdNINF0/VKkhc95LSp8fJVPqj0H7R
z8Hbv4nCQP2Ybh5P74TJNP6PQp4yJ6C5O7GBgmZZdkBiSlZvUy7rW0bTC/Tn6epgY3vCjkDcd78P
4pHVdAEE01Avpklzv638sPx8f8+jEt9RlQ8IPUNNdLKrJuh/hPnYCKGa/hJ+y2WBh5A9YiBGANDL
mUBD80LEtGdpp6QTdBxaW1UP8Jiugg4+CfwfRgQgY+bI8LQtrGj7wap8/2vLsDzrUkkHDCs9GQ2w
EzO6CI4GYpmFQ+jQHVdDpca9Hqe26jZFEygrjtMhJnjx+rs4nGAOWxob3ynKejs7WU4mhHVNcvdY
h6rxCk7sob5rq1LZOwmcb9ggupmwYiqnZuiBGrSTyJBPunwNDVHheykBtjnIDGvqR3y3b2uyNAjG
j/63U/FJ9OYVHLUNjmg9/CHXG001EqiCswAaqv1mmaqz3iR4gr/KKI+6RLrUB4Lx7CLr7YYGXEHA
RmdQHAUl5XAscZXMXJw3mM2grEoBMMqJhGG1NMh8hyj5J6lfXmenHyNb3j0VClHn9s86C8nVPQ8/
yXRmHcOIw+qSM39/FQueWlzVzjTepdAOGU8xBPLxvDwVb7w+QHGH324AbCLqgNPpHhinD74aGjr/
CsP7r/qjkExLKiht6coTMHsn94hjIORH9HNtyUAiq5izuZe2hJHsLjFrqI2/0KWP2jyeVWq/0WbT
hPtBLB0qosZumC0hjLp+NdEtSkmBeHF47qbMSzFTnq/vXNNJo29NNELOvlrS8F3sqGs3H9tcAl+L
HgFuX67gfW6ZjdaUKJm72m1OK9CXkSSrC/hK85Sybd0yfXAnEreB810mnR9RFlADjJAgTrTJvvBV
r+OvZR/sviB/wx9xz2g2CEQB+SJhYT0/JPWAwj2A3035sVBqb7dml80T5dWWo1OZo65SjQThQv5Z
150AokVvA8C/La/+ryES7z0C7SPBguP48R1u9/OUEBO3EeFxxquhvGlb6kMw84LRhCC1nvT/v0vN
92GNVInODEHF6drUBnhw50bKxHcbUCLonQimLibaxkBpP83iaGtG3qCKlyaVTxZPjkDthQVzNo8w
sGel0lgzHGMaefxApNELmOm/gRbnA1IFmzPfy3TF2OB9h/nttkdD3+6H7OIFy4Je3kRu1gwn/svy
LqqfZL8H8MsGXnR/sOOIhds/Hi79hEzWZm4PhsVfgZYJgIXZXPBM8aDjP4S6sfOFYusNcr/OeQSI
jFmt2w0aKJbENKhcyDxaOCWqO0QgoD4ri8SdmKhdYX7XT4mJ+4+i2sURz0aXJbPHxUZTjNhr0fE7
ahnq74HY8itocRCdyrjAGEysdsdQD7V8NLNYeAZRggjPs/CwtfMzhbA1a/8Mu1rXFc8TsMIY2NQ8
ikSdXPvTKVUx1r+ZNCt+htIM7yOb5VJAkxaiAHDnsH9ptwTZlMXSItT1TBifxE6P8AcbX2nT3SBN
VBdAx51HSPW6W2QABSXuNvJ4fxcKaKL9/9K4qBbxQ5Cd4VtEv1r0uicZf0a7CtOmwoHYvwWmxBrZ
CiOc9YvXNJhy9X/YmnhnruK/maLuBEBBED4sOqgqG850YflWyVcCU+ihN2RBxf6dROnapcABEQLi
mzAyKCjniNMchVFDhKQhSk+NHCTzeZU2ok3Dz+xY23ppCd3Z5FkCNQPlLRHRQBFG31RajzLSL5Qz
pATQxhbqPoFu+LnC3fIlwDJLpN9EAB0ab/ugijurSc/ICEYowJtsCmi0aLEu46SEnnz96RQYISSd
40L48KRUfPA8CfCykDbjO0aYSPi7k3LbAhDFqqOs4Eo1Gfmb4DbS66UHY/vj9i3GYsXlCyxkA6K8
7oyXB/mq2CDKaZrUorVO6PQyrIhJHS/d1Mg4xSBfUhsUpIn2ee9pcro5JJ98lF6g8f8ueA4LKmvB
mwFXhly+8LQcWes3q38eMLmCLrOpvHL22Iqemx5LVNjzzBYrChiIuPOY+bmZ2GP/v7dVJzBWEgWP
6YcinySgHsQL3XAxCBXCAX0kOAaCwvtkazhATQtaRs3LIKybgF4Uez0bO+Fbgrgv3YtWJjrq+SX7
FK6JZpg6LPmTQCQ5BtLPtI4z1Ys1Vl+KeNPZaotTjJ+pzHISxGIsEUIYzwB44Y5nyL2Uw/0/wS5K
B9udP+yVHjfAKyQqv4ROlbDTrDZPFXb8aYHSuc56aF2f9he/9XzkUAh4c6H/DESblKEOSA4TnH1H
8xKY03F1gv8vOpYhM5ybZhiBPk4HPKfvNj3OOFAefYI7C0TfL7ch59wkGRJfOUCF5yGziq+caGkU
qAdai91+/pg1BMwLHVwdD422VBHcLlu7wuY8UG8iA6FZLxNSf9f1FE/eJEP7LGyUcy9vJHUuJABQ
NktWDf4V7HnjDJ+b2GWP2o4QUISsLrSaUm0BtCPz9lnGU4xDt5JNWxtUmCKvLaf/3lwRDkz+RSuZ
aCaJ2XqZj3UYt8zOonA7qF1UsSbgKWDGBQmklE1LB3F6dkcRoBFBCqeNeEenrFTYK0feow/P3Rim
ypHb/B0XXNsQCgn1/n9/sBMtyOdKfyIpnPr9I2OYwa0ZQVkGtgWOIZw9b/MZxqLGGlui+mgZhYZQ
0TfU+ykBDXeO7DpG3g5Q2tlYU0oYidT90Uzug5Cvrh2f6gEsi7+Lq/GeXR7I4O80c4c76AHYteTe
YaCagFz4abrhCFuRuu2EBoV2WbekPps7scLq+wvpZksInwvCIJ4ijQs0oC/4ivJlkktHMl9O1TQ3
sNFaxBLX49f6xzj2i6rIs9FUEizzEwwSIh5176W2wRxGs7X6TiYiqYWETuINFnTjC+PIF/MQt0S7
5WIZGqZMyI5PScURdZKt1tEAzguxUf6GrQiQC6QxPO8J6Jhg7R8jK0f47gjb1RhJTPHPdvwPvp/6
MJwFI/Zr/74CqNuvDy7r1Wmn69CxUpuk0YYIpLU6bAAif2bmUXs9VW8MRo4z/QIlpuoXOdxf9+3C
SVrfAvr6GgS2ChngWSa9rl5rd93CdRnE8i2ZXGP5MS+QzsCbvXXiPG5ofIAg+KFK5L/CMECUcORH
5WTyL2CgIsBJZJKOmLv4c0tVrlAudWku0LXcXn4Q3UZ+g5/b7Tx6GuBfGkm7Sm/6FzhjWpeOPZjg
l7wY+I79ddc6RWoKaRVBFW+rYlPRNjIf0GczkEgUcDFglDvDFqrQDDCGvg03Cw+2XSJOD1OEnfmp
wSveMDXLSUW2MbJGtZAqP1cnsw5T8coMKb29MMdNdKXHsBwYahKQ5Lix6vWdUJ36atH/62AkNYBa
PchS11+1i/VFviyzo/dPc/M8D5+NgDHfpZoS9+JCu+6jLVKRbvepfugILthZLWyrgYWK8cCEcL4p
QiNdpBSwuoJQ6tYGUYUSszf07XTPOGxNiVvtszTliT0d9nz7Kh1DTUvtROt1urYGdQHPuK3PowYV
fj9bSqz3QOBRuN0XKu0V5KlsNm4780mjhFMElAvyKd4LNEzmMLYGQcunP+FG+VGIaUikaCQOd8ai
iU68M9IQXi7PYrFO0bgWSv4iUfI/lKYrJ06saZ3Ceb/OtwhvvNPe9AMrL8npKzNu9+lN+y6SMLmv
k+V6iOiGW5VH9dgQ94NT6H/ly1l16ksbvS8udXieA51XIjU/YBAbB9hwkVR8DY2HJ3xy8kji9OYc
fUF0G7ixVYa5t+ac2nyjbeBfZJaE+w0SRNjEwk4+b0spK0HxIT4hhctirlqzpNVLl0kzhCIq9gDY
sg+jTZyBRdBlVXDdHJR6D+XVRRUTKkAMb7n6Ngc/eapJSxTV9t7SaK1gmwgu5/TudHc7vO2FTRkp
PhUumEDDjt8hD9j5bGoqPG6j9TjkX88T2jGm3U1aIRe2CQx7jBNjwCmwZ8btI1cjxfBPgaQ8K7Ms
bBeTaBNUJmdQh0LE/VKTMHhBduF5wzumeXDU950WnvIe74HHl6g6bWQ+PuqmROP6gQ7F/ALoje3i
oGhFi3OKaFHaHgUJ1RDVKPdjBL+odTb5d4r0z9Ww3Zf2N0YqL4Aqqo3yuQ1fcrTB3I03aXR3C4hK
v97lIzM4ryqey9kQwdK9cx2snoJ1F0LW5jR38b9Nt0XNPjplsTORwb0ykwoyOTsFSs2mhCFt8CNs
g1A2ircp3ELNOFXvRmRpJeddSNdmJvY1OhocJPUCszqsbODn8PC1bT0OWtykHOwF7cf7bzD9nRnE
bIt5OjWuRqKpk4BwYFXM3kHhcaVq75HTC6Z0lv732jwfSLdHJ+0ITkVuuGRVflARQmwnXIWh4sop
y00xVoIS6o8oc3CN4RnAVnsG3ySae8jcoLY1NtTijErXDSgZlYLO0J9lQ+y7zmo9/wOlca2E6mD/
D22UFUBAYsA621sXCH9rRYQvtEkqpNsCDrjkIXMPmL+mIaSxIAuzUCegJmEAYZ7BTvML4utaxEai
jRHLD0Q8NABcjkQnQWiXPvz46+S29etBsaPI912yqHqipmEHN1dqGqG2SNvOjGqyQGEPWJLeZ3sO
FlSMTt9ejWR56aiR5ExWkcqGL7lkqOBB2NeLoUfy986XDp0q8ao2BxZDX5ADPTu9ugmcZslmLAqh
674tn8HtJTHePa37m52RnX8xxjQYLPLE51QWPggXwAeQSJ0wfbvvHGM2t8yvNzf+XYacckABjuzV
ITxBx8RstAv32gLnb4JFM9oBj0Fo/cdndDqTGwMAOj2zzeIkGETn+wJdILxcr1lW1dnOuAsBGN2i
m8T41ZDvyzBSyKFVEubKfd04jRdCODBgLsmV+F8Cy6UvNiFo6CmOq0Sc+9OF+y10a2KGPYGSbO7Y
9uEopFB6D+JXvO9/ChmkTn8bQwgwLJrDpcWT9So1BcZfyRmZlwwxVoV1jp9nz1XmOnM2I6mHH+jE
ttD4CUChRqIQbu0V5oLqqGZAV2P3MaS6/R+t7HzCwG4LprlnjciB8HTyyNIOb1QiKM96E4Elkn59
mxcQXF8lRgKmWUakpCDro5E/HdYVz21xw9RCey0jp+ehpfiMuGCjBWUcTZsEyKDeyRlWKmLH8ack
DVk8nktCSvezzybs7uS5aodqltapygOuJvIMt45Vp8iKreJdXQboZdTOhXuCEPr2izM4OuRWjGVc
Rpo/PmOnTm11foHeCkL4WKBZvh8rYKfYEg8K/G77wopN9DRt0FL+kDR4ZxA4F+P84oM7kS1fwmDS
fa44K7r0EQqpY08OAb1PFThFKabdaGqVsDByl+JStRPqaaVZzW3au5FON8sNkNNi1o8GZRS6PCYV
jOMIih6m31Q5j9yze7bjtXPpgwaNyLAdS09aOREihL1rbMCmz+tA4PsgVYzZJZoJLVy6nZzw+wE8
xPD7s6s5Cl2Tk48T+PsB7PG0uB8l8vzydN1xT3+0Nkc9GRbt7u1HbY4y3eg+n0JAkGqZ2DTFEg48
V3Ne6XDGXoyhBi3TuGxe6JAwtQU7eO+uE/IfWbk/Y4mxmdWtvBjS6De5MvBb0O6DukHnV/byYU9R
16X8u4WTZVWAdHBg4nnC2qZVohTi40v2jS7UlPUSLRJk50V5fJYl1zxwxGFon2bgFE2DIpKuBoqz
H9mjVDarPqns6saTSVXAnkUF+S9GhnGZZM5/9AF3L643r4QWhh9WeE+4mE9pu1THsrVJUm/wcVqX
60YAF1OvXNpNIghtaciClECeo7IphC3F9OFX6H3xV+g6EdBFmQdMJV+mS0DrZokA1nPujGISxFQX
Fg9YtZ679sIV2bmJf8W8uJM6aHzFqXGj8Uje7tvOS7kA7rNJFSa5Nxr2GfqLg0JhTbhlm7kNjoZI
CpuqPFt7tzCxZ2GKmPg0HjEcfRAMJKpCgT4HyYoPvWxnJlEGRR683YlxJz3XY9Su6x8hLlToJ/M2
HuJA632cd9I5+k8ba7Lp/ZCmGx0+5n/YRcrgVuuL497x2NPAbfSjnB3KbyrKvgqw8jOfopCLYdn9
JaaVtUs4HlW8dpQELipAA8lw74d1dlxreGFBjon4yX/hRXO8frBaxSZxTIIsF1aotp0ECK+fHsyP
TpJmnhLD+g6JSKkUrEDT8NCtJnPdJug/cU6gzgz/aPhmicEN3xtUUjfNlU79XP9vCVE+BIFIowNI
LixldEYZkrQsw/TbPCFStTywvO5AKaKOJZnasV8WDPooOhVD4l8cFx2iGjwxa2TIHqG+hjBeeuSp
Y7e6XSSuLEq1l2vkRSG+kfG5xz7gHW1LVh9xij3SOmYHKpyqPluHKbfmX/9o9fQdbIGw7bMRi+Vn
MZkSOFMkN5tTPwWyl+unU3qdKDF1FmbM4PCnyD6bc2scsi4uEEh/Yx4DmdAKelLCUyIpJG9zZ5zE
X/Rm+MvMpCR2Hzr6MlKlJwrojgc5Ki3hp6i6IV7wviCiLZFuHn5gwjPA8+uM6OGoUDleKMR6TUCL
U8YmsuDuTFv+g9oA+/jmWlfMrJwaVBLLjVn7zzYbFmQF7amB8+7UDHUD9F2yfigZMTxgvB8wU2tt
VawnWN1vlOO4WE35hkHV8FTy0eOTbtlpzWuqJ0S5EULpPPMaD/j4NMxrfnirJgy3hguy4uVKzPFg
vrbQC2DngGY6S6etxHMmYIwTx61aLHtrufCGSY6/ayAL93a3CMpYsC4uOFuyv6NFu1cNSkjzdvUH
49uCytgQVpCcbwpHn+CgQhUNzeK0FfPRgKJBEyXbMK2h8D9tRoQ/nQzvMPclJZVuU99oAuBnuq0C
fbn/2QD3yuotT9/qojEiXLxsH5lzLaW8zvK3EPHY64Ck08TDb8YNk4t6Pcu2bYHfdEUP5fbAYyfd
MRrne5K5eyxz0qjs1qVyg3aMY8INvXAaUjJfhSm9U+g9tfyE4kmamvtkOO5mchpdN73RCLhz06MD
jlCWNnhKS2LX2AKdiJBWR5R1GAUlcVZk9Jfn+isNXPM0nZGhAQGI1jnJ9vYJAb+9PrphS0MT9S/p
lluOggCPPV0+S17+TAW42PonpGhWf/egadpe1ZBS60vWGPqGAO8e2RcxXIQq8WOr6M8ehMpLD8Ug
fdkK4WpYmL1IlpF6ibF2ZWcuz3lFo6CaTNPDUI3AuK5qR8bj62GJ63WBFsYpBL7Y/J3dQhY7iXj+
peE4AqFmlY8JF5GJhEx6t/mE7RXpZMsweHNnaMEbpGkYpCmw6sGudUzCAOciy6ZGdXOLwPrgIUmQ
Vw8Hs0eS5I//EVgAraoyqOlV9DQ0E005ueBXBnKSSMsF7vZvBEU8A3Kk0pXVbRG9lmoBz3SJoLeS
SoPEB3KnoEZc8FOBblpOIWUydIbBYEdHLB4ow6WEDlYpUOFrSQcm+2sna33gicVMsbY02AHm2Ps+
q1tZSORgb6vXW384UfW4CsuQIBhY3mbkOgsB7dWQCosrKLxszgzxCSWq34eQ9UP/lQJfT+JuRkq/
e9H8+Z14xAL+qg/xIzVL3WvwD6jriZhOhYEoUMHd/YIy6nn0JSy5DQ9nJtcdn0pPkVCniTGaw05j
SSbc9v86eKsHdC4b6UFkj5p3WvuGeOlFdtnYznYy5s0ElZ7J23XbPdcv4AxNdGQ2doK89Jz7iVet
627wDu5oSGBb2J26hONHic4iJ0n9hfSJ0tJfJtbstWRy5ohr6Ww/bQFDZdxF/6bsgD5mUW5GgRRy
Z+N6zOOuTfxL+BOYlk2sL8wHGXWc2X8sy3/n1WM4EwcA4pfV51HwWWqFDUIvbEXGIjnAjnSbs50F
XlI/BbT0/Mh+sY9f/4Po+g1gE7fl9NIojdYjuNqooNLiHITBrNgCzp16J4gZgHF0V8FUYQpgHMft
W8xWsDbb5Sw+eNQtIcW+fPICqrLEyH7nEQ8LTxgwmEMxuvq0qD54Oj6z7KTCROQKWV+/PPz751vl
0rZcRWDTZpYDIJMfbB3iupYxevZGPetm6pipTCKgZOwZYJmZZnsewpwwh9QOfGfibKPjmIKCqeMi
+ngcz7rfK0JSxqMJY7iI+sPx+ztacL7y4gL2Ylc/q+fjsWhV29dRR36LdXPCjpU88G1xyWzgtq+I
5u58/T43DIzHkFMlGZZUTDjkJuaj69yxUk2BXd6LLYESrZzzApvOjG4yJvlRh6Ou5DRuXYj2x8DY
0gi1K8+2HiF1v1iRyzbgDVGjpp7E+KdJC3Ek49ZGG9TX5uVNphy6YJQJH4FxtY9FaMkxeDO7o949
pkypSNMr5SgJXDq9Jilqmej08KPSw1iz2n+D9iB3PUlVWjRmubq3iHyiCXJoag2gA9+RJw74YSG0
R2zr+N+RaxQcK69qVaJE6lvQVkXSslveWBjIwpLPlLmm5X7dUUmmwZJmVIAyxyxvDrysNLzoDZQl
zrsE2hA+rqKo2TM5EfRUwNqx7uXJvrwc/Gu1aZc1nnCYC/kkBlHH7oNmPwdEOwDPN/BDepal3ZkS
YakWDYPJapB0nepsOTe5Mq0sRsgVS3H7xzZJ2JHN7mJo6H1MWRfFSJ/jicE4R/+y06gxjDh3Fqgv
Ekja6jnyw7R1jVRDLh1D9IZ1yw6pg4dHcNfYqf8Trz0aGG1Uy332Lx+5wkwWrH3ThHeb7+p/hG+O
uwUhOCcalQ43M+H7edj0UQ883K/f8UMIJQXgT5aTPgCi6zjy2Av36un0QfxUD+mVWueJp/OlB56h
OkuRo1KFhm8mc7WdLP4xryxQI8sVrTDWon/n9INnTYmIQ0T75BCybHxtzZe+1ahqXOHC1SZMV3cV
sEVVut+a6lsl1QpMpz/lCKVqyH/0INUtv3sWtAnBzMYU7ESAo4GAXRWZqUWjJ3XygoTU0OcPW46b
2zvNHe/n+7NRWNsPn4Z3Jfyu375kaBfWBtd7Uq/vh7SS6+wrdG2AZX3Q5ddwyBO4+KOlytXyof3q
f5HsWB90VCUTiJrMs/9z8CH4SwQF7GzY6ow4NL1STgdz5ZlxJG0pr7eEif+SjzAqPu7ElS36iBUO
A+0B8id0oLlYo1vom5wTHwZCko8VVwaSiq3XvbV1QgKJha7FtuXha+G9IqHIUq4kGaT8wH23rG2V
mPatM3d1cJ73ZGw7nYlaAQ6HShpvaceSd5n8qnV0ZS+S2QDL+TdNnIiYPfqRIyLbC4EWQejyps6y
TP9MI814QWophhbqjRr/wGkrd4O2avMvvi3wOKN3u8mAqq4OOm/1i0iTtR8TxMdvdx0mGim4w8dr
LJ2oEneu1grve67Dczdog+8AoRKJlSgg0rngy/+pWndal/dc090N+aragjyPOEiHGLJXtOXf2rkm
LqGd00/BSHWSNI/6I9BIuDBzhk99mPzxsLucS135IX4O2TgdhijT1HkkSRxJKA3NgBMSQ+sGcCRo
BYpWg7N0BxxpvoiNav2aeqQHdmoxUhqJdP2MByVx44rgrf9NDUM7Y1Gq2gyycAM1hpMGJvB6ulEx
hhuPvcnmpQkT8WFHbNo1cAexvLwVVGjJZ+iNMm4RX1/tYfIj2WoQYTqGd854jF6NBQSS+P7IIKR5
upIe0dOPDVoxSNzEShPViWv6eop1oB7gQgfnFnPNmc/KRLE2B+lSmVGEwlnqiTNt9RYTdAj2+jpi
SaCGg23ECYkqCRQ6DCszQjIDqkaYpJq8zOqsYxu6L4cDM2liU/p+uyZPnWs10XMnzfeZwCUMQ4ny
TtStvbKer42SPUXGpC97pQ6ncBmDGLQXi94OEbmuEL6ISUp9AXfRSSK74CgdIwL4ZnZquB8jY5z4
LVFwDT/qHhXxe0o6stZBNFoMwgwYzy7Xsi479zCi9TXsLIcM0qLlQA1oNPKZIPGbHVTQ9rqu/znL
F1PAD9ZzMs0RH0PBfwOI26Y1j0xwYS752CKaQHm2HB9+w+ADP8FDX+qTSs0SAFfkwAW3ESYpcKH6
KFIofn9wsZLVs+V5GLwUD8vSGCE1/aFX//3rDMifCwBuciIhBrjQo/HtnUop6MAY1iaNfiy7E843
+81sy+np7Yi0JocxuU2TXEj1CdImoDsZ+SMNhO/A5QXn7Ba3rhPIrqR7cQGDyWLTzu4r348Fntei
7ldQmxl9sR5rhN28jIHqKVforxZCBxSs9N20QcE1HWd8qCoHZTf9Kq9nTxPEnHww4OrcJH2dQPwd
7ViO1m9y58dNX6U+Jwa9tSbkLTvAlFv+vXY0GkU+/mWz3P3vyaih5TW9+DJk+LdyKGB3F8Fktn8+
mt5JhswRGlP8Daz8rZ0Vu1s34BpHEYrv6Gq6j84vwukX51KnLn3az4h7u36aNZBHHsJ2YJVCf6OA
uGOER9Jd/7sRMmDdkXShcSmT+Wl+iP+7dgpXSJNHNndDs81YUs5Klu9rvbczMsA4wp4N+mY4NNts
ouNz7/bENwCtt7q0T9RgCwuakyvVmH7jAPV66Vfs91+OWhOiK43fTXXe8zn0I7xx2KNI7PlYLWKs
i8sT8F3cMxMVTMsPhDL7gOc3gqZ+PjP5tPWaUf01TyWBCcY87SUDuIk9cnSEYIzn0NyMZz5Mq0Tl
CSP7Aje27HNwErwAYAGZJkW+0FNea6eCuYNYmovqKScKCXZEj3HId4zzxvWsePot1f7Um9UubnG2
5Lo/dAUXFEMea5JoAdgvjTQWhzU/26OsN6WOviI9CX+/oX/oY6MSkExzEROv24YG7/R6jyNcG2jY
I9CWmwy0TMvuQQrarjvbDBCpO3D65HHx79JH1RKGTQCTvoGDZ9O5MGa+c9TJnXdwhDF6DJtGm3na
n2vJQDmn+1TQc+gNW7zahJbF2vNUJagHszKkhrXEoz277YCO6XLO11ZhTFwgIYxf2CW22yeTWPNQ
jiQcuq2H2eKDTH2wJoD8/7FJlvZi9UELJ9LCRhZS9nx+rCP77lSOXPkNdloSidm/mgD3RJi7KVb2
VL3E5srv2nif4HGUyD1ckxbwBH71EPAyhY/hDh2Grw8/SdEZnx0lHTOdNh8WmMrshhYMG/B9Tpmp
RltHlrSIrnlx4D2wG8V6t9FSBON18dkuFL+9PTlgKsfcqhe9Cg148M3hpaoWLA/Xzh5IIRKmPrl2
cMRFXuDxhraAuPgLpl5tl3uqoaskQ4rOe6rNuut0Mi9e3i1yMEbWvAepZMvdJvnb99QrscfgxIR+
P8SAcD+2Rd1ki3vMV3dkPHtPlQaH6Z6e7qEZBkhAKGPEx2WQpjcknj9APaJBU8h4N3QqJpf2h48Z
GkbhpxzZ2387UbzXg7qTS3QGIZOwK+4WRWdCRUEYVRySzghNtI+wyBuxmhOeT/ZnELAel/K6hCvk
kd9nxR4+NSGqgCgW5GAO7/tXgy0ol9CqmLbSR7RO0lexY3nN+7Cp13sxGQ5K25DheZ5dRbwbzC2Y
lT3K1q5e4KYVh3TnCUiRXTOs8ZY962QRj196ov2WXVv6LT/TCSHez5qiNI/IqYlNbBVqjCzNXOzK
FFGocPl2fWB1HB7LT1vBRIrWeGfICFKyVAh2Ugg8veCi6DDZ851pY6ZVXEj5MvyhXz+cESFfqLrO
dmSxcVONhDlfM2WFAbIPAtqziCsdCiyVkvoHqEME+0KxMC3Vvw4aO3EZ/+OSoexfxFjyvXfKZjXb
fsLeH4lBUoEg9kayE0LHMR4PtD6gbCQLB/oOh2igXlv3I0AjhVBIRzOf/wp4ZJ11aRadBYTz64cb
wSVcj+3ZRK4ReqxxBSs730Vt7Aib3yN9Y+Dh0MIsxuERRSM44Len9t5JcFWPLedi0kxOPHhwkXby
/0IBl4B5dPzMuCNAWFBRh8dKyjed45eqyBatG7WAmRo9qdqH63Ldwfu/j4Zu5672oNj1fBKF2VjU
BuAhnnfdUTB3B1VW42TY0K1g7eRipWRRXbayVpZhwsgJsxDVd6H0q/2MmmAFxIn3SDlH90wg+7Za
/0ro6lj6GSE64/9kMl3dWnz0C8HQ0S3Dmbdyvo/8i2VquQXIW7D5DLnsNzcdBJ5Kc3e4oII62u70
FTRiVtf66xu9MexfrRUMumhYQizpAZIEQMUy1DqzArPJiL20pI+NbioDcOaVzL2a2PGhh0fTw4rI
BRXgI7jWmj+o3wMyh7IsJvqw7iVC+HQIosw7zgULf9wNS2n1T9u2Gpj0zaChKSxUjzmcAxjEnd87
U6zWw/4b0yFQN0iu11dStqpn1NcUFK2bbKmo2ABt9IcgZNVX9ieOsnaJrIE8IWE/BY12UIh+5sL+
yjL2XnM7M08SKHrf/1aGCMEbifwoyOBVAsHcuEd3AKnTuZPSBWKQb50fidD3CfVtknqjmq3PK1hd
6WyfLcoCC/dzi0FHdiLd+1w1iaOG0t4N1MiRtbcrCOY3+cwhaNNI7fwQiskHaC2IM+xkuiiszNRb
kEWGbJ4sSDAuDxThA1RTTZx2z2GqH1uzRjiujBlk7sXdkPP79FxiuVptPBBHriQrrzowURL2szbJ
jp7IYdcUcVIDFufHwnwteRqGAitXYBd2XrX9/7wQH7WuC7a9jvyb87k64kBS9Lznb01tI3+GJc1G
C5qBYKsh+buvLgK3a0NOpHbeeeZ0l419Ns3MvNTAnTqkgn5cVtVo5mOKHqaC+sEEuxF6oq/oYtL3
kpvAJsKTlB+E+MSW3EAfmtT0EF6DkURcWgK/sSHT0Vqs68PeGMh3a0p05/S55sJ1+PZ+y+6cQndj
N1cwD+p1XzqbEYxKJ6/B8YsgoacLx0IErCchhTyFnJ5Bhq8QPMRf1QLoj4OnbKWoGhiXbgGwTjPV
Z6PpQs1DdWCfeO/uRFCllmoe5JqIrvZGz4ZqQwqrpYGV4a+m18KzaULa0yLsOifrisCPGokXkL4B
IOz/gnqCG7F554pOxotF/QbTmp37KYCTCgZG82Rx1PW9iNbhi93+6QqVfsXHNADRuEJOyy+q7ku8
ZU3KJAN7mz1f9qO06zOXZhVekwqS1KKY1HkUmbmBBsQWEbC6IhDRfZ3N+JNWYWnwJjZltlv8hd/E
QqsMu5VNnGS8VAv9HF9rRDpvYWBXvx7jCu0CxiRwM74eRzrq/H9psjrHEJHle2himyG5NE3v1dVV
9VEVt0mGwgdPU7JRc3s7Tq8I0NZqag5kluGuZBflsrToCdxVjFsKi1y1B/jkpaduG1XP5o6hXe4I
3in7TDUE6tLQN51AtihXBhRVnzwAJkgo9C3UCZg0zwNC+KxYZJSGsrAQNKys1Zlwm85g1pP4bcj3
kM25l8PGw5DEZ48iO41ggB4Jsd3gAN6BR2AeR4fqYxQ8G5wyqDX5Y+5hRg/MGKJ3iU12cYZHRj5O
JtcINQCarK6+yEuXN0qfJl5m1nOnZDUFnyH537sdPj1pp2RszyVEpPqTMje8cT68YQCqoS9BeSZl
75Nfx05nz+DBZYyKq47It/aiLYhX5bruJxj8bo5CYMt4gh72mTcHDkMlJawVAov8nMbLYXLjANxi
1LSFXg2/V2QQXleNCRVWwfJjldK4JPuv3+YkKwQelD5z71jppVaGcUZqAogJ67jpAfeNhYaZFoQS
kTLRWD146SExpEME8hluWtLKZ3ywWQ1fmR79agVNMcb2o+1eJkU0mY23V0xhDtB/iiARa7xnSMWG
Dru2385D6HIktxIPbyrrUKC/nDdyNST3YTSHlExIP9TdraINheM5PxBMPzpCIXuK3xGN9yqAedcY
pA60WeH/h8HICjh7K5+l6ysJcNZfMPVJWMz80T50QgeNuA1cMxttO3fU1Yl62GN4df96/tnKzjdS
6cpYTwlAGNxy1Vhdj8SnqReDN3BYi26+75ED8dT07m9mo6pDkHbuO7N057x9MRZP6foxR08J8ANx
AabDbe9eGbLbQPjDeH5uqsI4xeSL5dC7mnWYj5f0RpXmoKYTnZ6BwjvfRi+Tlz380fXQQuuCeNHP
ODPrDXS3hi+PDLU3pZeHx1KX8w3gxgsUlQlkQ/RlfuV3gB9BKwkZvc7+Mh6Zw6suvoUfcQ0PWjk5
+yDMuRF32+AgGFBlryeZNEIPlvvyZCjCVxdHLKpQY2oqY5S/nkVK/lmFpxHEJayetQDd0wqX1/uy
8fnSjftkBjVVEfv9W/rD69jMvgDz0MlVqNEehMJemKK2s2Rh9ov+95kJiZQYYN7h4IU5XpKi9XwP
Q1Rdkz3lV50vsNC2l8wgWUkr/hY1aY/YIf8s/Aosz/W3NNd83hHuuBtiyLAnWMpkv9XLuo1YYXi0
5obdsXwI1fb7Yiy9T97om422DHFt37o9ghnc5TYLQAT1l+IpCKwYgu2IyHMJFvyi4eug3JBc7OcA
7aSUUItFPYVrKJ64eSMD8sjG/5i2wSsC+uZFELL2HASOHYwQPiot5r0GeCcv0t49eBppmTTbndNe
2wBHA41wcSp/YYmGQpWeU4tCXdldvsZ5UN4D3nuPS7YJrzfcDnPsmWzSPdybg1alDdv1blOhiffp
TKYmh7HvFbOUGPfx+PceTG+2IPfciF977EdFim0lL9drwGjzutoGuVnvG4HqvS1FExDhtZKHtJ8r
vi916UplwQf4ixZAVwfAF1otU5z65kT5fKgITOtIA//MIuptlK1ZzDyEPh1Il5dqIc7hmx9RtzaU
Sz/2UjlEey63uAgiz0MSmmctZlAqCKk16SGZWpYx3qvASESmlwW1JinXZvg5bloXHPPwe0ZxKw36
RvP/Cy9GXL+xbvF27TAsytHq8DwzFnWARWXtQONAD05RBSjL03HSi6Y4Saw76FB1hjhy38zqeJdE
pNcqRN8tQy1lWF+x4zATsPL7JuIVdoaMVY/zOHkqmy45qoRknuNyPO43jO2uT0HlsDlQzRDW8j90
TTnaaXTdcJIdgZJJn4wmDEtv6WaP53PZ9KLg1Elw0XTc6X46PxwzWQTT8IGnQ8I+AWVyU1WSuTpa
ykbd6AceulrLKdi4uqJ3YbuQFo3YZyHLFyIrb0+mkNeryMoFPk+L6diKJiIpCGSTsLst43acRAuv
LZkxyM9lJM3/3j/pJ7hr8MwXBjX9dUYd+OKLSgxo1JExo2qhcOT0q9Ixz2gjm66R9pTCCh6fji5/
ads7osEdY7oELCQ/2btaBzT1AxCf1C5MeAtRykOABQgKhwHUv7SRJuFKB4hh6bBUturIxPE1Z9XC
I+NCXlb8IZ/ROHCupLGPfX0S+IWUJmV8P7OfF3LCromJZdlf/N+97mF6GbjGYwv+/IN5BIe+RPsL
tCRMoHyQHRX69pu+Cw5FW0fsFDSV/oQ5KMmjEt02jj5pS+yAieN96Y7VqG4qvVYC9LYQnKHhQBJ/
2WnwPGLJUyYRFqbqsB6pu9VTIyhC5X3/t17rvOA1j0LdKzb/zECu7xE8wFtYzgR3MNfx0kKJIgnx
3jS4RPmSN/1vr4rj9VSmFwv4N9zkWPVvQWsxgTlX3uAqYCu8QzHQUcN/PifE88+vLuZmfBc6jwLr
P9h9KDJYvBpxpUBEiPwPUr+p7jutOdv+O5M7nypqL9FDHp/5satSAMewWyAFROIm+Uq64fuDBmzh
iSK/IiU8QPfRJ9zpcc0H7fpj/pXT9yuzUEIsnGx+Eva6TR3qMleXoBGSVsWlohuANU96fsA9q1Lw
Yct2XQuF1Rm858t4/YmyqpkeVQWBlDKkC9Yb/U9mUJt7Hua5VjxBQCekrIiroO40r5FHz2pAujXZ
ZkoGmYP0IpyOVetKWHDl6MxectQ2RYLN661h+kg6R02dQKfNDOoyF5RVMI0BULrdiqYXnmhHZd8x
QlW3x0g2pBoevlxVL78jBPFhz6QjLLgoI2D32saGNxSfYIPbWmeIoPAv4Rn+r0XD24JP0rnQwhj3
7iG2OObBbtwvLpDSmngxp91Qf5kqSZdc7agxfYpqKpgLrmaaBExugcSpLdZTSBGmflVmWZIBWSYp
ZG46I2LscWr8Wd2QXVIDAIwaIyHcUkrDOUuBQfIP6eIumerjrO3tvG4M/KIfDH9AWOd8e2xCIblh
5x2TwgcDzDcSan4xBaWz2c02N6WLDduGfxWlHczzYsyEstuIL95XoZFN93HvW1llweIQdY4vCeIi
acoM3shqdCbGafKJDDCuIcbgrWjTJUW9juYxI5knUuXjvHwF5YjyfJzamlShyiq8cIYz7G9wfVXF
rI9w4YKlpo5pjTGTyQxANChrnfoRqcl1MTZ12JxJZ0U6cFHtYARM96WXFuB04MdePt5MyZ+IZuka
eN0DP68rs2XKxi5PG2CnnbEyF5uEx0XJsujcidTTaQyJXuv41HG9Vhcv3ugU1et+KyzgZc+wnDaG
Mv+nh74haAfwRjKJztZG8UgA7Hw2/QjFVZ2uZpLezzrdf2m01Ilcq4CZ4n/w0uMfZJAJgOvgIn6l
NfjILxxu7Y4hibVY4FN/RY5pwo8ZHhqrhwlG1O4D5FdMTDLWkDhZcePG+xzxHvaNKpOEMPrvKCaP
BN8wJbqZ9rZjnJGbm8EHpD7VOph0fdDroIoeOJjOGp1av/FWgTEBDwsd9KwzY81nVgvGv28HT7wP
5HLEGE4Lt0HsIMCLV9+14kQTPTMUf7vYoHh+k4YKSqY8LB14n3cQxL64sZP1LIPfw2zNtq8rAuha
KZItpyOzjx7rOf4qbxL4mc+hZk/KYjw9eTOxCwVvDKE8zM1d0sGohEww4nXTNfPScVRADjJiOgho
dxTDTLfSmsIuwGoF779GZ/BUZyO8ofjQz1rFKGBhjBoQQkvCRNpVrWx/VhMDBXv/QJWarOCKu5Ch
lJAkb7O7isxdHwwmlxQZqm0+QdM5FAz9523n4OGsooAEVPcXp4aEx6m8EJsHUkWtvs2wXmJ6AEfU
ZB0gXfA4YveA1IxFDM+iT8UCpr8GUkv91Zv08wc9Mz1V5nEx7xF8xDyc/MYeTZaJHNSIb3ElGNnV
pdOHaA6sYOZxTwjvTaBCc6c/jWobhnhAQp+KOTvSRdyqTMDIcbCSl30WwTrMI0dwyv8rsIdv1ABB
M98HGFSIC3Iqi1S3DE15JkIF0aDzT1T0nyKzK/AQoFJn8xvwPHSvZyBfJvHsRIuI3S9LuaIyVgXy
AAJ8ECZrubKwOJ4odX1q6Egs9Q/qinwkVcxrxt7R7NIBFRFN/EB2ON2svNCiFKuDRLO02qF8oZQH
gAvP6xPgZgxgwI0axxVzD+JooX6eTRXO5fu3fsApTIshz/uAF/p1ARm8ant+46JT+3Mx9KD2JxQx
sznhMfTwPfpcy9yiY+se+WvykSY8IHupSq+a4XD15QV4rmHp3YJz+ctaUhFgGzAyRsiLuBcmJHGr
Ke4GOphnKph+WWycYCBTaq7KzSwarHdRCkQI40qba/EJu4aWyiVFM3u5AoBOn/DJu+1TX64+VEfm
cl4TSQ6nSnBke6/4Jsd9FXX2GkY5RLZqpu6S6Jr5/BRHqpVEJv6gGhFnuPsNJWUa2jt/7rMrQSBU
qKC2TI1myVQu+aIrbo327X9E/AW7BgZeq0a0z6PJN/MFchPa/7+aSQc76FjQRYCLojKsMraNiN8P
6ZZU/tfGZn0vxLeBd7WKSODuWguTZ9LamYr8SuM+cFSLMFt0qA8p20A6UkuRUr5KD7BPvC5r+xC2
+5R1EJXW53j+980Qd8Bo9TmDI9eiFNl/ctgHGLnSI5uU+3t8UmgwthhCsiZJnz8DN0sJlH3rCGzH
er4oO7ke3PKIDjxgjaf0upVpd8HLEvY8ugUl2VjlZ7aqSuNx0r8tv3ya1dJ/3yJv7M6KiqmdI5ET
3OCWTxWAjzFHCTyVszE6l7Zwq3gYb+NMX7VJnbeCgz/NNsQtyhe+dyfVvwKPJHnRsvU2F4iCgRjM
w1JwYpGzh7Cv9BqfTE3+/D4v2zzMH3HjtYHfzHBcVzOZZrSk/Rro7il8+pe+yf3YqG+/EqWaB9aO
9dbuN2N1Q+fqZaFZc5SHkK4i8SoMxfZbmpDmVpeYPGEqohVvdnUd5cC+AarYjl7f1RP3D5t5JJ1l
n75TY5t1yVdGwIENNdX0NdMb8vih3rfRLsiz0tsEgUXux0lmGhvTh2M//SYG35rBXTtJqyDBOTJj
IgTgU7WQjvA3RZJ6YDb45bPl9PL/ZPvT8E33x/MeA+l2UcRROhA9yxqgXW9nkTNPTMZbNc1jvzUW
nL70D7ABPBmTurhCGpibwVFqkrZKiA81dTrivKzXe9dQlID4mxm7Ck1bSQZCWFrA4DBhsRJly0VV
us7eFcmyCeB0ei7Qg9MKWF7fXR88WpOmF01hzr1HM1wnquH3Se2N4DgRPMor5eRNiFDpiL6L8nUi
sXY0lOKuv868pR0nyYiuB0KqVrj6rClVPsIHFn2ReBnwNbpiCunHfKsG/rS19g8GV1nS+0nKHOLW
19ZJXKMsxSKQdB4qammSPWORTk51nasReiY2eyplOtWDHkF7/c+1FVEBnSnrUVha3VTv0WRG75xo
jr6igh+YAgD+pw6RNzYx2MzCCIMg6mTRruy1U60eWOJWLMCYs8Cu9ZyjcxfpxkY0D0qVzSuvXQcV
BAvQDv1S9pkRZZjaoNcaRRH/r4ddWM1EwlS02ZvuDNvLUROXVPDsX5TckyQiR+UmyP5vwfQ4o6ZZ
nFBlNnyNqDyR7uBDVyDaQTlEEi8RmR9a1PmK3RyGCN+iqSA+mjeeVYb7boULGYvyUCA2xTIKZY/c
scxUnddD4+JlNytLkVtS2mWHv7S1eY7brYBgXrBSn7LwPatL/s1oP/rEdSi6YZLWpOeBZaqlD3cp
EfwdaLbmVNidbhOEyTDi6cdL/CXtvbEQ0hmGXbYzta5oQ/XaOBTuUOhrWq5VYJmZDGPdHnnp28x4
zrxnCgEENCvPS+3TbeQ1XWqsatJlt1pk7VBFUkVL0DuZUUfUWPVzutVIeXFSdtWdGBoBs3lquLvh
R018lHib21h4Uw3QmQatc09aYZzPOzU5F5LYJ8ohB4R7Bb17tI85XnrNlpL59ZoRcZguWQJtjxvj
O7CI6c5UkZb5C0oTWi7hlfmJYW/RGvJgfUE9vDPLivKMOmN6jQvTytCTIUTQMWIEcXJWiaeDdSJr
32Ehr02ZBzMd6/YKdWeAEOs2o56hlKiwrKjJAa3m/orFyqLBSUOK+n70Cz5ChFABWa8JW/pox7Oj
HTApZDzkACQ3xN3O9b0pjTPR4zS9UgaMiQ8Ajxp/MK5g7536JQua1KddAjt4EoMsLnQxjmUgljrf
YU++XFPlXaMaCREqDM95upWuysV/D0AVuU+DNckwqSG4XbrZXR1cL8aA/2hK3duYgbchnBHJ1hq2
fbJv/kTsCqW38JGteWhShQBGjx2PAqHn0UMJAb1rpenozwSBhqWPc8oypjhB60OgUpr4ILPZF6rO
yYP2CaMNiL8lDP+5XzcF8gYGVrnAxa0MySdSuKvwS2xKG3nuAgV4pld/FFYLpgA/sx8Z+yYV6XhT
pgDPAT7/ydAxbXZOdQYJ/OAYGU9wmPIf8OIt2sL0pxrBNVjEohZiSZqc3neSHZ8agDeGr8z4UX+Q
JcVdbj1io9/C9JQALQD/2z9Xua1sk0bjj4f00erWHbAZKHua5FBgvNAOeGcnY4wQlggkxkVUFA/c
NIbKOQB1YJCUQhtF97fdt+9qhZZXGR1w0hqPpRgZxrZoiUUCC9f9NxiwxiC/U22bSzwLYOM9i9Ee
oQfnZOJG6Sa9DvI5f4OzDvehygIyOJxFaSL6jp7chGv67Vd6xz7jxAq3srBfYGu5cjGXiSpYiMMA
//Gwy00W1dZomf2iOGii4lObasnsfgYNqqD2GDdo8QJ/Gj0uCDo4K13624Ht6DLhaSbXRDQgnnEb
/OH85Kp/jiroJ4NGsqHHvqkYwJ6IKT6pnx9nw9IM2Swvl4WskaHV5xtAee7qKA3ViqhZhaB9ZMq8
H0MZkAWT7uHchI/n3jNKRNp7f2XO4WdbSsGydryHvgi5DDGa4+uU2UwRGV4fCbVzmfRyV++8F7Di
70I9kWoOLrdcHMuqpzToRQtdG+3J14pVqFY54nKwt0Mjls/KLqwkE5Zp+bF7hayLEYdQaIb3qa+G
8ykm/m2p82bKLHjSkibWkdwUgmqDjph8t4hXgMnmZ6vSvW1vu+9GuU68CWHuJcWGntc6klUYE6DC
tXlxJQbl6n4K0N4b3qpgZRaXjJEwo84OzWA2SecBct6s9ErHb8DeswkxVUdj3iyTIOi9POBani8N
M24OrYvA648F+ANfr6EJ38WwaSkQX7zex/R0s9oaOcBJU/9lqxuXczLg2gT0NlIZcM0I3J+48jwY
qavKp36b/JhmoR/dpc9a2TAEXyZwzLqXQbKGDXqz+zeVatR4Ywm53BBdxPXq+bpcx+v8xWZVjmHb
eBe+u3I6MSgi4yZ806f8kKG5RhZ+Dy3glJ7MFjn3CkItrmdnvOcfyrEGNf+oFz2u62q1SmsSAB5Q
CJ0uLSPWEDgyscEriQV3oKwV/yN6SFwVQH4pSen+Iz3xE7pLtteyudFOiLz/rUjdxT0DVRyPqnWq
lTiYuV7uLVFU2Ptpp/1+FzmvhXtNczI+tWsVwAU/970ASrLKOvIYcrc9KSvaLHrGU/nYtxG0W2BY
NzY/4f4PKT+v3EbkvdsayHSG/4gvL037wVyo+zkVEfyz8W9Yu5QsQ31I8q8wcl+aPO5RFvRN08ng
0D/8b+j3RMLv+xnhvQ5ZyZKJabztr4TwCtnsoyg/Ra7n11YFbvh/pQ42f6vBjJZ5in4V/fze91pK
DJml3HUdAZlMo2O5Uchto94MB0Zh9RKQUW0dDc9XN/dPCJkoSiBlZ64Y/rO97nXKC2maQ0Y8ixJK
rhY5GVyhGiT8QUsKlliBQDdXux+YO3z97Qa5CH1+1WkSH0a6Jg2acGGOyfUZ823N1AWaQeb+zhj+
AwxsBTtLAaxibfqJOR/YK5qckIASY+k4W6MkfVDvx8Fkkdgy1cvBmFNNVwhOR/Q7F1NNIY3QqGqW
7PMfjsAqAhuYz0WngHLXwJ95Jh/Vq4nnvPG+Z/S9CBu/BalIo0UGO1MJtH2pPOFqlZFcFGxbac2O
UMu7/or74uhgsxomB+hVTJSPYYiVVE1KGge8zMt2/7CGiP0kM/+bKiWgkgvSPE2KbWk0WY/gjMX7
XaqgTB6Wb9LZ+jAKa9kxMwS+ufA/2kWGqB444JvbGMn5R84OwaMVw2CbaZ8Rf4NmcoR+60MOtxfp
rGL4qNg2oKG8RrTRP/1N5L3lWo39ciS/2cNZFAmLwBFlu0Qq7xm08n3DS0uCHUwJ+HxaTil02whx
30CSNcmt4kYIZHQud2y7lviRRFmoMTJpSOUbGvFLYkp6uJ3B2stlQbthJOsony2qWtPwXSx407om
G5GEd6TtzCNkZw1LxERwmhqRe90FJT9Bi5yte6+CoVrh0bDIsEqgjZCxxCc5OADBVIX+uK6KnMzG
7u/IcyaiBRfoqED6/uNKoE3va/vlt/gKpiYgX9+0JSpBrVVJ4OoH+0dR1FLAqchc9pQS+um6Y4w9
Yp+lW0XUGeg3iDbmXBwPBDK9O/w1KLSCro+0JbEUu0Sje/bK8HZ6vgLUJfKFEXf/QeEfIGgIr/0J
+f8FnxE1UquL7ZDwyw3W3/oXUWiJRJzd5cHU2q2dZyC1SiYIWz4mpR2nZsB08//rc2ewZuY+f2uo
LEljL0zVyO1fHbefAS2EptneRoqDnUxZ8+n4KYKbYZjmmuZxa9jaGx2s13QNHsbi0S6JEHaB8abF
IJJDuu5xah5o7iFMVDbAYffc2Ee8tkw5QIUmGnaC6IApNcvcpBzKXTZghbMFWpY/YWhEMwACXz72
ZFXMLBCh6OXU8bFGAChem1FqejiJMHg5ujHVDaLFjIrFdGVnXEOHsKQdp4iZxRCvRjnLGMdIMyTV
H7gCI0SI16Dbn06jxhDozkA3NsIUQlgJsIFZTUi/RzpFYQXzYJqs6oApJvRpSOcPLX86iqnouLPa
AHqGC8TjKEUprmzP6gLueIxxIW5AZCFWEH+GcTHTENZlcrrs8DKwB3b9FQPuEk+i7OsdTZpBy6MQ
0s7DhEMv44yl0M6eFYwueUBVMRddMHOj3mY5hNaSIQ4f+AkLxpdZULRLk/QTkBjAlLj3+FJV4Nca
QFfzQErDIGrN8hBbGa9Ig8JN5W5CkFVdqxs9EIeh5R4FO825jMKtWkkVHsTkZefEB2VsuPV5wS5J
t3xvzPYTzgPKqq50JYO4w/9Y6pQ8JDep5vwiqATcwR3xUAlm4o1rjYVLTs7aGDRFFN2/GIFAZsVH
5JEFh4hit8tbon90JyWRP24Z/R5T6Wu6qHF8CHl+aNX9ZQpMK4YqNbmt7iiEfTGsOubkzs7LFhc+
HWADxvP10CPOIXvTi0dl6AZgrxNcMtAlG2lqwf3wJiC7Peudvxr6CQHVp8SrFRd1lspBb4o0BZxb
BCDKmbRi9fK53FFoTTRUfTsITsRNzNYl7ZcwVGcAAtrY16ENWTdPhtsBAwDAj3MmdEzUNYdC/NE7
C1As7x/2+Yqrh5rOYnOAvbYs5HkfSFHk4kHF32laJGbGqUcew6RP/oatUgBLtVBFzzKGsoDX0eGu
2MD2VOikT9ciDg4qqZ2LFVbV4MqGp2xnJkP+ng/Wt+R0OKpxmmt4RJZsvHtTJmd33cUGVA7ZwhC9
uz/pFTwxsLV/3KCTTONLCNJsfV6vK/UKQsFYTUlBEsO1uvYPrv0GfQgyb7pJ5WClqvAXqb9vaRCX
O+JXDDmNUtgW73h7Y4pAgK3otEvRIKyPGpyyCyeiz1tU6YGQHsldr6RxSjsi2nVDw1HiwhgYpu5w
qoqfmt2TqzCHxcckun5EFWGG1U+CMJP+cR1lT6Aa3S1mFeE8IZZKgdsl/3tpPrOrw6czlkKQNr3q
2w+10yjrDscW5ve1ip9TE+iqDOIw6LyfybM8EZWXJyOiDh3XYYQzPw1KUOGkzwCZr2useD0FF4ES
cNzx+jCjboJWcr/fG0QHwbzbQXqzv/z3t4ga8EDqDJAIpGTMQxXMeabsLhcrXr22BtO2JExbdM4h
3fW8wRKDgrQDAKOToJK5L+mCzmMlDpUb02xqRnsQ78fEOdyDt/xJkgW6/hSQbHp8orGXnyKAa6zj
Pr204xcg4T/4fIof168lPcXYdmYnJzeThXehSc4atdW1tIaE5uTXjggN+AkxnHI3LnAc46WjrLmL
UOmO81vWxBInYwTyUqpWGepoHy/e1x1i1Z4h1J5fRio8CNxWjciE+tcak6nSHF5iox4x/TOPQpxI
JhXZrEeGW2eO3DLx90b2N08q80QOOmuJADns/wZGLiSJsUhxogF8hCspX22aSBDW5zXQ1X9fK9GH
/1IWHlT77QXBhTNdalVVfAdrBcjqJwrZz1P5XhuXbVUv7Xnu2QIf6dM2Qwo2mbEf0WaTqiZRMjIC
un5wdf2featXkVVBhZomDjbiPqvsbta7XKFXo0jUJB3N+p0o30Bh2uldazOQlbagHsgBhqxfStzv
G6f2ic+c7kut0PDeYziW4s+KmwgBmcyv5UpOV7J2yxYuNAqoJCiKzB5tQbkLjWZOe4pxCohjYl3m
dUpx7vSBqymNpswiq3qxUNhiRC/ju/3S5tzBR0X9J1yqzk7lsJSh4myN+Iu/hAOfB4AHXhzP53ZD
80Oj2aMaYz4BuDxbd6JP40fRuqdynbjuAH7i2TW/sBEEAM+ncDJUmmo+ADNnD+cG23XlduG3aIL2
4+irNoFOhXuADhA6WrZGXD5X31g5q3ktCUkOpoggHaf31mFcFA7YnXHt2gVCrDadnAsw/7logg0S
jot/GtqqFkZRKg4mDi9qnCcXE7bHTzZOcUmdJuMNHbfh976nmK8Csf55Ct7MmxMY7fFgvXPPeLk4
8HLjjSSyeZTAApDrOhjN5xYtOHou+4skPLUjJrzHUGgSbnLcUITG3mSgkeMQu9VQreZr8mMA3PkK
rNu4NRnLA8tYuXnCYeed65iN4SYu5cESv9h0/uPsDc+5BoqR1TLXdy8wPe6PuZsgAs6y+v0knlxc
zLgHNIjGnIIZAY/sthTqpK3pdpOcSE3IIem3bgfrqjOR36RjgVEQ+Q3lKnz1F9M67HM1jOrpl/HK
vDKY2kKE+I2Q7X7o1q95r1OEi7vKY1D9YiTHqdDXsyuXlMNETI4AKJTeAynLaWIwuF8iHKDaEDxT
6fO677oZIKokjK4e2VHq5F6jJRrMeRjHPnMoWCFrewEui6QxwLjqLbOlPSQoCfkyep/0UckNn+xj
4Lesuju8kidlYeIDLGtmqFIUzS60zc1oWpwSRe1csICsxFiaKmfzgQWeRaeG50gc2pyxO1KmfR5o
XbGwxE7r7lwgedFGS6tdmHZElA16zbAxR4gAliHYtxJoWUHl+lHsrkl+REPTlpAZlTKj/sgBUs/+
jtnGCxY1l/hZTcbMdOp5GHZXGHveMLfAZg9ebA4I4nciOuWFlOnHOXsd3KB2w9WICWsP3lfP6De+
R3ZaMNE6gMmflNfAnWtqNIFz9NiVO9VEcjKZ36MK1EVyDgbNrLcj6qkKd9FyqbAWOSNNqAhs1NwL
UDcWsZBpYnJfla33WVfrtUzQkFLaPfLgPKJI8Xb9hxSgqdniZio50u+YwINlFHh+lC0BvlQ+QeQJ
fxQryU3AlRl+OuewdC4+1hcR848S+hxXWBQis6G4uWkyiNFpDDdZys8AzHzi34XFaijg+7tXPnTE
lNILK7z3m80ToiPqcFPc03ndlvB4K6YMohlCDIXZRGjFg8rp0QK78glgw1dVw+sB/Jzhv17xXRlT
8AcTEaeMQL+MjfkaiheZkd0ruLFctEjG+mnSCIm5Nbn5BKcSSkg3Nii8xOGHpdttPtRnQIDCswwk
MFUylWLsFIdvuVgf3rJxmFYehT+oTRjUFR78Vs0niSIEXwJhoY6q68p2j2HwArtiRKheIQ39Qa6B
5YimA+EK1/avSx1xwPVieLb8Wrnea3va/fOFPoH1BiKsx5pDj9Cod2TXf/oU5aQxhyUQFCNlPtxq
a5dt7hx75QJgSAXX0YGi6MuP5DukioCGR6ytVmEY5kKgOwsJrE6hbpRlhhLmpL1u/DmPvkHfc3Et
PhauqruJ+FsGsOT0UzocRtQqhj+bTh3BPVGWYlCybTkOUMmWOPWmwdEej5NW4X5Aeweh4DnG6/hi
QAQ1SCRiYj/aS0x+7zTHjFFC8wRmewE7rOZGX4SZeqPjJanFwFRkopP8q1s+7pqgNNN9eOWstdst
6UEQZyL5KKqgvTChm4mvz9DA2WuIZlr4UxbWw9aJF9kjxMTNdmg5t0LMTl4l0QuRUS0Q0kGhrnTf
Dt5/NbG4bgUJqwyuhUAr/PHkUxocDagqVDM37fgqF1h8d2Y/tWpm1rmDZLrCzYKYbMJOC0/XeOPk
yIhb1DIueQdKVx6rR/98/eQUYPaaUi+tl10hWGGceyWbbU0oLOh8witYrRRpsXJxin3wnT2Nu44Z
SoMYnrIRR2MtzAw7iEpd4huwbzELL6zwWNobfjN+TxLI1h5GgLOtXEHeJNgZpXqlYqH+jTHpNwFd
8VNdmsbB0NpuBV1kOrw2BcnMuKtszCBknLPXsCE5iiimcKP7aaV45c7mJRd/UzE7VtQUzWUyPrSu
omon5+f80LDjkkWI3rpxWhI86F6sZEAhCskg0IzaDlSp909cXMcmLfwV7ztkcknnCAkYxffnmuev
wtUcO7r20eDaSIfTd//vRKIArbJZBIERm/B9K+3cHONeGhi0I3+i6qgY88+wtefwX/cEdp4I4yul
hPohh+7vNhq/VqSXri116FaoKV//0Z2zJRd7A5KcPNiXnpB/XEJuii0/GOKUmJyfQHCecibNyxGt
UsWEoYRuRSK2MQyL7E1fYu1NQU9P2Czow+4ZwnvCMm8NsYua3JaLSu+FKPfAjbYgrByCmXDhTKKA
aPFC7SGc3Fl5/u1cbmSl13+0xQg2jWdOZ+jXdFYhz+gqZSPMPwgqr4ejDiPRqrPc0oBgSubtWrpM
WDRU6CVwELVpGPKgVbXijnF+MF9oA4rNgZnSnUi4xk/OpidQs9syKguhoVhljyjCszxhcf2/tLp8
Y18oFrVSVCjigLLYYU56tofJxo/Oym6wyne6gSwO/LJsN4EhedxA/30lytJTWki/A3EWefPlfRIh
VscbV/J6JkTx3bVtwvS97AdEKYGZ+QOtvjUS4uLwg02xovm8HDgOsvkRKl5U6W/+RA95xp+PDReu
I7HB2c1B8aKBErJihh+h2VPZY6/4eoxI06cI/2FTQQ0hB/vUNmE3QplITtzt/a1cG5CfxYmu2Wjn
oSjJjqZqUTxENJpNKrKWYT8fC+RIvkNa3n1i6p7OyWNZxWFWFdkHk9ipsw4Zr4MoA3BpB3QZDVgk
vGkkehSOJ62BdE4ildLWfhL+NsyENpdBKlmVgYd98DzH3KqlWyrb5OEDE/nHhMD8QkrCO6PqT+VY
YdbB6eyX/2ec7YBtMGwXL5nmg8Vu2H6Vq6mtHIRL+L7HnuYa97HKw1tpd874BoVPZd7fRp53cOUf
Fum9lBjzIKb8Oi1Fws6V/iRXsMXBiAL7e2lupRQpoWGNy9Ss3wupSBeHv3qTEo9xnamwJEgQh0mL
2pTjPRmfJeU0FyB1y0Z1JA9e2TxkRAja9XnxYwIBiWcV+Jn3fX6fhPd8r/AN+ZPOmhCN9pkop4dj
w3FhS9mM7mu8e9TmB7CAR8crow4RL8zlX/6szQ0QAypMSm/OMCer6Z/VFV/cNI6qFqlNCi+PocZj
RjTWIy2zmusR/8T2sYXKQJT4urys85lK+6+0X1IE0Yuqh40yHxrHtBgyktBqAsXp0FIJDzXZ64BP
AOMJhPj587LnnCxucDPZ3R+BE/zYmmvBQKRlhSrx3zhmUnZdmnNJWx/sjxZRiDEB2rjQYyRhCTc4
bsh9OH4fjFsviC0VOzNymdbsSaF/QC36owH13UF1n6tR9uL/4WwrLWlrDv6QuXaa/vIfe1hnevT1
3kINmLdARHNUPUrp8DiCL65Ux9tKCx1Qegjm8HX6NscB2jIWEfwNex+c/3ijcDBFa0V4feubiXX7
ar5xJaVVTHprb5XU7b1uWmTx95+oNZH8PuQ1dARJ+7qH4KJGtKGGRVgQqAuUiSjoJV2u8thvOcTG
JeM8Je8ARNmK4ELjQigQ/vSRRd5UQeSPEr2RSAPaTY1OyKXnc3mkDYKyoF6QjOk0/T2kf3eHFKqK
we+YWz0fNBA61Ri7+iSDjeoap0iLkgUWdZAmC2Lk7pYnKlzWbD7nGswxZNmA2fWF2RyS7x4W48DD
zvC3I1LaFKG2O/0oDXnrgSStnrxCc63LJUmpBC6qMZfV9OT4JD9jrlDFrqi77BenkTPkDJVjkTH8
dXLy4KKxZryXYQDq+G9F2HlhchR+IM7LJLoOPlOJhXD4VX4XS+T2bGBfIxX54T67jSwmKUnsX+ei
fMq+pFRczYj20RyM4azQmJHh3rJ1xPUsXgQIxMrrnuKNq9vkP+ykARcfbe8q4r0aro3qWuupsN6q
SgHnavnxX5z3KwqrRfwiKorURHZHytYKpGJ3/GuylO8jkPRHDJ2WiVzCHLWe9hZl3RS8amnTf8lr
L9WkNJcJdxAUfqHdGvHMuTNbzbBbo9ecrnFaSdUswbQOyVuiLTnO5IemRucV+wmVwEh8vTNwGutM
ZkKOYaXJvEvL2BoATq02lwZxhNK1nBXZol4V8XaNG0Tla0zzxRY/KhcoOvsA21Uh88vqZm4iGk3K
D+E2Hzx98Y42ZTSSeBb1Z1+Tvan0ouE8P7fjoHpo4BTFAPBG2B5R/ep4c2XgpQxmg7Bjcp7ZleF1
VQZSoyj9SFwzeodUuwS6zECGoEwqc/S292CcJnfXEfD3xR4OgyRrnT/wfwxxtZ1XYkxJ+8hTddE7
gBLzPO4Zb0ZHMcruI8eiYAOjMngkpIvuxh0l7b+YignynjshGVTTg4LL48q0OioNOZuBLs8eetC2
YQS7zli16uMeAZnUzfsGtxAUfV4rqBSdw8Anu1NutVQYM/GbMT7HNgAOuAZZRr4J8qEgb7YmoADs
STWhqMy+mq6OuzNzJqEzmrE1O87D0WZf59Yl8N2HKI6oerekO5FyJaagQYQu4tPXXBu4Mu8gQM4B
X1Ilv8UaY7WhkN39O4ZPk75oJEc0ZgdicIstH9qJXsNiOwSjcYSWVZ/fwDgzMMxuO6Fklnh37ivp
Gk0dW+7iPDriS0F49nfwKCv5cP4r61uSAvWWZIyqjXc+/cO3CJ9XVa82qyMzIUF4rtFURjMU78PC
29zE8pTciG5gTBx8ruxs4pwEPC2+Ta1nosKizucoGUG8SEaX5Yk4o023cO9vjGulC7yxb+HB/yur
EK7nC6NeyPH3vJHLLKZkBER3WwAjxGzHJH0niaiVHM9UvsSz6s8ovj93QhfIKz4+JWdHH95Qb6sV
DIuqwcoj4Ah8Q70KQ862u8n3Dvn3YpTDgzdPqcEIX06vsMdaobiYTpEi+v7NHU165IJKsYK+tAOO
h7TEbhK6iB/VVyYx10J7/ud5qQ99tBqMhe9UPQnXHnOBg248S8PNIbB1xmAaj3zG8nMuNhy1kG8b
sCvRKaXlLvTMQuZ5os4Az+k/x6hQwZhk2ecogXStjN8zJnPdeMdOZe4ApQ8BivYSL0khu5kQ/did
BCa+OCAxFzVqZm5c4/T00xguntPWMV8G1YUzrN9uVb+nX6YL0/6+xhLZMb+vwc4byaazgXPJi3+6
0oBZJO5thjZIrDhFCcumOka/cdHdWtTLfZPk90ptywCUuc+Jp4XZ7JxNB97XdH1lxLs9VPQ2bkAr
12SOy7JZVwUFKFMVvK03pZVAQVx7ayEi3MIXP7S3ymm+5JMW7pPMyBsA/MC3N5T/cHyuMakrjx4y
zk/J7hD2qTHSn9mlu1Xi3WFhmALhTSTuUpAGVbwj4BVrnzxzcpL89hMBY8ORazMwja5FHwT1wJMi
bVasWFKGnRe4IjkhTKF9JlqjE8ORboIDeEiVp5v2RcyvvKBMmBTlaVEKcvIRO6i2eEJNT6ARgxA8
euJOoMNHb8Rcm5209AUxTsENzp4m4cnaRQ2GkC3LJDG1svKQefYJ2P/8kvcUTOJJdVH3mG5RgHFy
MpCx5RTRUf/bdDR5foGyI04aIofdxCi4PEmUR7pvid+gswv8Z4TkPuvRleKAnUSIcLhGlbU8LptP
0zVBB3+0MACN206VrTl8+yBqRAXsEZN8p+Z23Pti1dGvbgfLGzREyvdxhaP3ZBDUNM86HUAsjKxi
eIXQiXxIlWfWnTEIxAFkox8ekv4awhsk5SbwarvI/oSrU1mAzIur9NcZ6kYB5oYeLNRAYCTf7Y9s
dSR+UvVszE6bireWR5XgSzyVEFaBNIuuu12qzUVa5n2S0KVkauEGTeSmRGzjBgqMgQ2sUK5eF8WP
J4cCyS+liSSa4ayOwZ+OXMUy+HUKPq2nbWUm1b1dl/gl84r54zOl/e7On2eyYUH8hmDsnhJ0eNC5
th6PUzXhhxm0JmOvsvKhodvoEHq3bzg8HhVokEoIecxxR8QPGKflzWSn0xeAc0h427kqQ+U4/Oie
SFAwR2gbcU+4uKiQr/F4mhCc9b6zkvGhxkoAye8+VZ3U0B8RI7USFQJmL3+jAIaMFmrIrDSMS87o
S4AwXAP915UDazGV9QOq15to9+DfP/59SB/+WRGQ1UBFCo3V3zUvvi7b5rOnKcrfQH7XyFCJkUPX
lbTQ9PFcjgjaUC0OlRAcoJngOy/kshh8YjKJ1rVJFK1iahEvo44zf6SwNGOJ+m1Wn/ryg83Hdo8v
HbB9eVSS8syJBYO+66oZgqB/sWmqPX9ok1z1NsgD9B3e3G2mjnYtGfHn6Rb2Uie/dTZUXhVImqSi
v77gw8P5eELylcH6AuZ6q3YP/cbvx/nF+IHW3wluUB2ovpc3p4sHYStwmVsYFGbyQaxOzoqw8Wde
YGanTJyTM0e6iJGbHt3JWCzQRXrKMcbUV1aF8lW6ADvI1yFRuIgP46iicUW4DvGD5p8XXS/auPwr
Uz4qR3BMFFs3XXSdg3rfOPaDHxHcMZjV/sVX4YKSyCnZaTLwTqlbE/SnkPVGIeIwrslZugCvjXn+
CeRpLyqAZZZChcTDbMcH2gZhGbYZWLWxmJYLDSF5DKMid3vv6MKfjfl87lxurI5lGUUfKn9KGRyv
AkiRhLCEJGpQwx1j+3QxW49NxGIPbaPNFVgQhvNIeyEtNpNDbWLeW3QIqf3ib4gd/oVylG5K7Qoo
bA96xAtD0odMTeFYVvPFQfVHyNn7kKVG0IAecN9eejnyQUgE5fY7rUMTSCrWvSSidCx/eg3mDM3m
iGaL8HalNBrHweHcwYxTf0tYjU2W8/ku9XL2J/qacVHzMOcSM6aAkRzXpyJbCz5YmckDV6aOdV6L
v+/BrL0wEfXu4cjzzVefZ+dB5mEggzhAwhTmOiNn5WhmXxJsmtdSFOe+tV2q6nbS9e9BtkL3Di9+
jY5FIyGGzKVpQAmYFWQaEiIDPS45H2v1sTw9W5lsc/sXzRklR+RkueoGWqRt2bX2U5Ksm9MQiMIn
m2Kopvgcv2KKAlTcbTaMov52mMNxZmpXXSdkcbvWBX0ubZC/MyJzQ5688KZag3t1CxtORJ77/QDd
wTzkO9b1FZFzt00dVrLuDOWzkU6r+uGc5HE6Ygmr58ekuR+nxPNnGTjCKtbfBlcA30GrJ5+qJOLR
uCJFkjOzj+G3UDRyIGd7g0fqwp+f7PbBjTQ/DTjLmNXhsDGp3ElZE0KZhDFCrlL/4srhScEjaFnD
ufMM/QdRlGwofPOLe66wNSbMeTHJzlVKoOzZ3n8kDMQQ1s3Ybz2sPN7wx5jDUPR009BhQrB79lY7
5MD/bIfHhw72pAS2lHzeCEedEuht5MdEGFXcg4rvzLgTjhEWScRQIoMp4Ph3WgKkIwx/bQNJaw9l
yP45YRdJcR6Lj5AJn3PmfNI3/K0h5V8tv4CukZvnS7muoBftqS1zy6Yl+tSyEfC66B1WtKUeZyVJ
YpkcO9S7GIDtge8mSNisu5aThPKdJXmrVLo/9uUO18wCnwUvH92Bo+L4xmFnwfa6nNPlPK+nYgzy
OTJJpyK4wSIWeS9/QnztBx1oV0hLYxjxnzCTwIGCUMq9ax0K3hXmcg/+PD4Vgazflm2+UpRoXP+M
ko6eSoMMuO5cBEbEnna39txNpyQcpxHhloJIV/s36mahzYMxbHk8LBILHPuvdRV9oNODgXVLDtyU
UmoDbN88PDgKQFMhgx6R4gLWrEQl2gYMiSMhxNUqILCqiAo9cXCNx46CBUUVYWReQdAanE1aZMXi
W0Hj2Jo61khG9gWuur904J1GuJ6VKXbQT4MSmkz71XFpp8Lg0p03PQ0LPURe06IeNzXbAkVhULV3
qmHzc5W4DlSef/EVNSdaJpFuNrZxI6EcH3sthLVwIwHr/Fn6SakFa2WbofavNU1m7THygQHLzJhu
NGV1sMUDIsO5ZhUS0yrKIAsgJaZZHoJGdNqig4kPasG8z8vmEyElawq55lsYrXZO1OBffgI+z2GT
SKVFxFM3YPqEh9xMJzpC0nfls3uqIOgXnH4XgtZuNQqk9g6/NHSf+J+ZgcOVl5Ahvq0xervcpFqr
f3MJ+1UKlVC4gAgirqrrdXteMNqiOoRgSiKWvp+U+vELe1+9pV7g7aFcbhJFDOGbdPRrzu+uCuwJ
btHxyJhmopdz6s0o+iprH+yRc7ijYGoSaKidnCHxnNX7DmkVD4mj4N+07BnQxse0iDBAuR9qzh6g
SbrWeKMVTcTSzFwXPLi7/xU7598GsWqEZNVYk20UBEoAmQhEuKcgZiomOQOh4MV4N3AcVA6vqdZs
Te1BrW6rwB08UVbZ1jzJv6c46v7dfS9YXgBrAnoVT14SJqnndUs2aCQBYTqX2Os8ocFBOnoK0Y+7
+lJ6BtVuJ91KT36hKfkTl82bJOFJvmQAcI67wdsczqiuzCUveSofFGqcY/KW5c6joPH2HBAh/s5V
3Tz8y0Grbte7u0EcUf5+zWpiC7nxGd2Gj8LuUD+csjZON1PeLDyZoNRiK+Dt9fHMA4jlkfALeDJH
KANFrSgoCWeCMyYGcsPXztTUDm5bkEBIA+coIG4GuMmFmfA7+m3JqaqlMM+9H0MIA5Sidr8yb2Hy
+0qIAHj3BaSqOEh7irdsB2XEEj6WeMJ/Pz6n9+BvDwDKJlde01RKW/WxNNtjV9KjVe1EB1/oodIp
6OuBZGjw6ZzpY5i3MKWPjPnWnckZmf0gPMIlvl1gPlPjuXoeH6DUF7tiqvhqnAaVuwGww0rXRmzQ
aqBBjj/YgpwtSFNnercq6e7qtohY9MxHjtQ8IDLWghh0IaVdxRDt/SbkxI3/0w1J4Lkpk1n8QWip
mkCnd1kW3VCGpGGilP5oSkNZ6ReOWliJ70tlqaObhnQCDDc6PSrUjuGh1HA/2h7WpNloPa32rLZY
CKahJKBQpA3rvQGMtzmakrFtCHEqllYSZDuNrlM2RbOIEA3EhmA3n8laWz8Sg4d6aMfelkeiFeLI
RaZyJH8Tz7R/IQZJUojA3NPdXynwePl9uAZbwQGtC81g1b3eR0JWeKHo8gYHejZ7cpWfRdpUxL2v
Ze67hW/iaryImvSD7GqpRinv2o5qN2rG29kdSQEGBJpjtDcnauziFVpzoWLN0NCjLraqAQJ0EkJ2
wKIqP6PK6JKPdGETo3Z5mb7FfU5BHv8ytQunbcblRa5v09dcX1NV/9YmDwqNN6XMNqc3RpbX42ct
D1W4DFddDr4NSDBpo2cwpkNT7Bd2W5zjwPzoS2+YsPQ3UMcFggAVqDMZ1qQtIBLRf5g6xZi9spzf
qTKiBUWcBkgUY5zvLXgt4kCaQzN8YxyH+0/9/tDpj6j3HmUbQpWh1t04AnATX7txEsE8T3J+8ct7
QGuXu60kwB2DzmV6YFVOP4LTEVGVU2hz3QB1Ardk+Q3OsruB/JhYIooXuSzLgnz/m00LO2mcquIu
KmP9g/KSy0kL2gm+YFaIe/exMlqwqg5o2a7oGfoU0tv7wiHKnoWYvr1MiaT7nqAt1LY4UbchXa2R
suX8umIl1eww7e3oA13Cn9tzGkFXaMblNP3bTj69lx/pW+Ntuzknh8bpJFhOHMLT+uiYf452hoWx
xTuJX0eLuoqIL9mkhHKcSb7q8MK7p2JeR8/qDeneKav7X7PLABbEooPrztPB6q2AJhu3tjJtZTZA
I8yGpraCfapM5Ykm2av/2335ujMV9M5J2r3Y53y+dcyELAwscTloJUNrx5JmGrq7xgGAuIwBoKdv
sO93omeC0rXi3k6Bu5EjxrW4CwAMD/mzDFKAbFgbHx3Bt1FxV/UJGTuRe3p7XKERwJZYrK6IEKO/
iXcSfn678P9cvYudDRdopQYSNweivbEyDwRFzN6AlrRrlD6ebmX8YsRRVgdIJCo6iADidsOcv/LL
3st6DV9oH1RE+jHtVcRQ7RNFzWslDKfPiXPnA1Mg/xkUIzibnWkYuGo//dM35eX+xEkev6BRsSBk
A6hApAEaVURVxJJ8LDwEWYM+xDyZ0Bcr8vWkQzgUme9j/63ADpMYUgC3LpoiOKFyfQyvpawq+ipu
z2wLtG+6jPtI8gWkKJwvGizu93ylt47qmV4Tdlk8/pR0uhMLVUf2Froh2zrA0LxRyn0dpnalykdz
3pTdxpOzFuwo4Ayrj5i/qYJhkC/XhGubSgv665Mh4XCjT4j5BSDToKMYNMl2RteX7+Z6cGEhatf5
+qElYHf5a0VKApRQLeXgimuAtVtToi2j+Qbr+eRFn9xdJzqZNdmoHHWPXkRYexFHKQYdi0h/jgBZ
uXKuv2yoDK3KMcHayO6TLVY2VCHVd5YvAMktu1qmTNkhTm1ld9Wkt/Nar0av2f8BwkyuDzT34inb
IzS+XMOBomAcg8HrejjryV//aeVDgs9QXYpDf/lowQn/6BITmCXDRy81L/ajA3FbkmJi4itUN+Uz
GwFu6LfGREFhdl8vKKTj6EcQ6tQM9121cQMWe4JxqD2L+bhz2hbmAtFF29+evtHyhXpXd33zmSHy
2bpsBuD6IMxkOLdYPGxW9YK0JVjKxOr2rm3aMbGyVHgOOeMXZ+Z/v+DqsKl5rudpfK5s3SWpOMMU
Ag7ci7CIMHlmiRUcXT7Zd/Qpeo8bxCRyfi8Fg0yCIjJgflSO4eX0/kd6p9fAfRBCXOnvqx0dp0GN
fm3PRiGbf9otoPnjpRl46VUGlF/V5XqSNhHE4ByJUX+ziefUs80nVp1Q21KmB1U/5AqqcY5CpAPq
ivgF45uSiTkkYJ4oSb2PZhycTsYqstsycjqxrw6qnxLgK5PKbIVc1eJB9ZZ6ElUbCPE+ERBhBON2
2futQK+Ebey62XIce/vNwhj4QDD8jEoueg7QpL7VHuSZ4NLTWY741rCY2FQb+C6rxJAzjSge5np7
pWhlnnqxYPUWRbJZvHubTLP11kcrZttRUdCWV6I1sFmwwZh1GWshNmTiM4F7BTv+wUx0hK4vZa9k
Lg7GkoOZn3hLjfmBdzMcFk2wjtkVO2Kke5otVGi5y7TnQKFme3Jx+ZAQ5I2dbe74mLnXrHvPXOGC
0AN8GhEDVD0aHmzNwej+Bg/f5Pi7IOdsc4mx4UPrnDM3nVCcXotDimJ6a++muoSI9Vv/zk1O+4YZ
zEs1xBScoSvEFH4mK9iCrXdzmhy0g3SAvXQe4IJ5P1j5sXkF5mCp6UNoF+KvAtpjLatOHTV06yop
yKRfz0lGf9qstxM7hQO2yu6b4sUNDaaZ49LalGoIirWhMx2dWT/jpTcXk5wrFBEP7foOOAKUfBpT
tRB+HPnK/oaPG3CBLE6ZLnggF8d+ZGUQxEjNjOyWBGWBYRU8wd8lwdsfUTB7TrGqSdEVM+UkxEuH
MvFytjGgBQiM/TaKlFOJTxku3HUOCaORp2GC900LLHdFN7N0RoUZ4ZFOQPd/0FWJVxpt3+Tl3DcX
pees86pA1vic7WcdthnIXKZnhyZ0MibQ+pYJ4UVRT/lIm9yzJ9j2EuolldFk89al1hmyHLr+xt9n
YTnoW9zoBurtq1YyvDCD3mbcXn5hcFG9t+bIvYQjWwN7s5MNuye60A//8gni0DdFcPT0kETynGIw
i/ghd3HXONMyadx6Gz7/baI8KKyqnaJ0qgE8Eu1g44SEZU4JPTxCX9+4UaYZbMxo/PRxM/3H/HQX
jXCT4+RDBJvCCx3dXnWSEnFvYcZ7f2W6Feo5YUf8WPoyWsHtjQmP2A7naPv0l3Lq8NFoMwLZ9O+7
DD4w7TL9l0oUO3l5WnYUBrRqD/PGjgctT+dZmaNbjvESt24UYsS5vHex4D+A6I1I/B1J0sIz+gHa
E3YQtdlMQbt+IRMPd4+Ct80bjeJip0jRwGUFsLWoxAQm997BbY4/++74AD4oedwz5trdxNR1Qapi
LAo0TChpKpxWExv2aikobEQ1dkWus1Tvo/W03nTnAo8h+qVBXXdkHH7yr4fBfF/2gzTlvvB4Gn34
bV0OISal/4YhwAhreBorTidoOVb6dj4E0BFmyTU/kBRDrkCLBYbOp/iQ/filBcMLubSvL+qSFTME
j4AlQnUUW9XB88GvB6b7zxBriXpMGigafMe1KZmblDImWFOCWvLT6GNJluPmcQ7TOXlFbo815mi7
zYcDoHXf3FcK4obzB+qGxgOsMqKT/4dT921f/HH3kQ5e16ohhZQ+5hH30iQpYhviTz2KFclI5kX5
WXLZARbOpPq/Uyw94WFmlDgWXhFb0a22SRohUMZUg/n/zZNYpj7siXouc0AR7YMD/wonhNJN6vsr
CMY/9Ut1MShcJStgu56KiQi95CjPOU0gPNI0w11RETjunP/hUqI2SQAkS1BrcuA6mUHPsfKy/0/u
OtOS33KSH9Z0owNIw9mVDziUH7nCkY4DYuZ2PEpQ+1w+Hi/Y4lPYFvghoX5TDiKBSdOUCwZFSFI4
Ss/8CJZpdcePRjHGTmfMBY5ERxOQ1pUYnlvg2ia8srZmu5l7UymvD3VExrMqgtK1KmR2DQvSNkWh
dEqGid0ajY0Rpg2MtvYYLEgYd5ALslO5cf7EtblT7Y4zMsTknxfRiOrvNlTQ7yKKWm1Trh4YippW
/dmQp9SZrv+szqNb3actf4mfHbcajC0CUpu5U0KQHjVjYoEe8Gt388t90bFIy/yxcxSO5/0FKrnC
t5m8tYLv4AnLfi74FS3kklkEbVrzNK91n21H45UDd24B0qBaSliEPQ1+mJnCamKeB0vPSCIctUZF
8ddFFvvTeiUd1hv3/9GVgZahCEaCyv2Di05PkbB1Lh1MFmnTfPvBe0+7PqsYXo9pr8yetOAobVxy
fLx4r3xc7mGyUzbVcbQhHq+dZaL8vSycdWsjmpm+qu9dkI+MIXc/gdinoiEG58w32M/wIE3VCoRv
qQDVAuWAeP5Xv2AyLKV+z5wKxiUIcbdm+cmYmesCfi2MdZdhpyxrwEDGMKXxvPbyJiOY1gSafRQH
N8hN5GUy7o0elqqS966UOEDcE1D3SeVgTkawP2ZbKfqt4U56iGW8EwZIfFuk4FGV2d0eQx66hVhu
uycM7QHZIrahYh1PHVx/mFGRS4uA3xLNQPydSHWYZrV1N4x9VA8Hpgkbub4SGXnds/8UkcsKG4F3
+Z6/TFdd8FB88rDcI46KIzuFI7oSbNJsKajwaA1x9hna1EBt579dFf+7xExjx0WbH0L4LaJJhzZ/
Se/JRokPMjqd0hvRH5gTftQU2J6brDtgvtn5LGdvTCytLOIVZyexx67Nx/OkhT7QF95smQ5AwnY6
UqL6+PKHXZ4kJa4eMl1qwHjk22eIWhsAcR/obdmfLeKWW8oAMDGxnWY9Rvp18sivpzJHrP8+J6Dx
NRQGCxSS8XS06tNnYjkQNhITJ9IEZNijUXEWIpcEwvjQq2CFmz4b/Hi1PLuki8+y4Ta3mCDPfhuq
4VQUeRIXcAVIjDyYnyFH/NTyzFcMKB6XA85h+rXjGr58KJ7Gi6ZNZJr1g+NlUTLoPpwZF5XjET01
CE8MlFrgioJuL9psL1VvysJ4VAzjNOnqce91g/66s/ZScEExHCGatceR/Jl0Vk9pcZOtqjObwp0/
uWG9hNrh9XvENsvT6/fxtbD2hycCSGtQNM1Om9zy09NhV7YYEuNXLSYu+HGCj+c2MbBKzkEaGc5k
iJ/LmsqmV/ZmOHz/RkhoTUYpdboh00pOXr3oR/b6y2INvvC1DV5uily0UjF1YWiiR3EYfozOPzPf
9FTNgIQF/zzwAoQusObVrbd0scIjumf6gaVOfaySTDklKfZ5rFpDbvxrLLaMQ5vi9wlcsDSgeoHz
IwyrbkefdbdrAlgNejDZiiV7QuPzZUWQrujUKLYkkyrn2J6W/ofNBlWAASaLCi5YZ4hf+qVKmoq8
2bWgXInNmSR7STXlgPLgmzPBgnqdqsFbWFDa9Ni2lJl61WDpHF7uvLbvUEn/UTrMSDzamWYldTzF
WcQAYllMmysElLXuk9xFtbHQx88rsswHCxr2LJQ6Xm4RY5Vnic94wzwhikiumj9n1B32Rs361lqk
gHo36c2zRMhGAKa2PbxD0HtpOs6VLXL8klWsq0W1NLGGKSmWONnsC3NLuwY177pStn2qJ4eilJnB
YayRIoKcPdbPQ29tQSVxV7yAZ8dubXBDXfB9lsBp12tEgK+lyMOL7HJ9xB9B0wF1N6G8oXwwvBRI
iT3wWezdPVgG7ZBeOymp3Dk47PxNS4AKQP/y90xziMJHBkBFJU06m64tPyRjXAcd0/kbcpexSqy7
MDMQfkioUIEffQFBnLBvKrkyYAJV3QSfpDsDXLmXWqA0cmdJP+FX+jz7H1w3z96Ox0FHXkws7qLs
lxTrE7OInYimneqpO/Ti9ChzPqOehawMfmrLkkVQUPPvzpH/78hDp4FzDzNWqBSlulvcbX0XqQ7O
21LaIumiutXkvUYQvzGwh5YnCE1l2yO1/r7g3HkpaIIZUoZm+YeCVeCZwhvn0ileuAX1ifcH58Mr
wqgwPDxdBi+oBWHlvem8CZRxGNJceht32PdI/4Uj0Q3v5qDnaahbZr4UrAyeAyVYNma+OUYmLwyX
jKtvJYwQ35nIMD3Qyj3xLmuwWG37+vF6lfKAPlIgJe4HUisSD+tiAR6QaAOF4HpFFWt1GIyuvq35
wupVgGaxA2DG1UQFh3gmcTyYRk+lWuIVGkfeB+0gs5Pjnvgy2xnrBmalDvFWuLrAZV2LQkut4ePV
UFBK52wQ1VTfXGo+L9vG6mP97eeFaBpsnhgDZR+PYa8fO9mL1uVZ5fPgGshGcU3Kv8LIbASQV7YI
Z49Tk7NQUxxXkVUp+CoSlTEu34DbqdsKvCfOiOVws00K1g1xB5JkjpWwdged2DUKg7igYUXchLNs
Fcn+MJpOlU2ROvbIggbLZdRH7RpdJGXGlgnjmK3tao97vrrqMVKXMzQ2kys0iOzUUWzhfXtoWTX6
2NDxbAXQ1g9QWLMIrHl8Hx1+89rLg98FjErGdPt5vnTBIiq8kH8buRRzPt/PrJfbA6+KIODuGzUV
utqsWnKTT5xSdM1PY9S9y44kRTgXiFH5UvMc+QfI39NWO3pHbW8hTe4DUDe8YVTnfgbL4xrNq2zR
sH0Mgu4acaUF+08MPG2pztwR5V4YJZHv/wBbDMXHbp3uWulIlRaSaarO1D6BSxfYUQddQpWIFrDe
qMZdEENYCHreuCeq81s8rfw/MK6Wb/ZRPLRvFqBtO1I9P6HrXOaxhEML/Uiw5G4ClvmqKPgZOAh6
Lra0uEiAFsDuQiT1KazdSS1MGhXtql+Rn4uLswkqjGl6nWdoatcbX1C41NUoPXQvX0H5CbJy5/xy
h9YyhIOLyKzkKiLo5sqWyOIujboAiFcEQxLiJHcMc1YqxHZq4zC/C6zClJIg+eA7dMB2bjOFyBTQ
N6R+NHxQhOaERTly6Qa9S72dlv4UymO8vdO807lyfCWhO2a7WV0cfD/atrohONqPkKPmmZcwECl+
+AhDTF+BRLe49RvCVVhEYtwo8HLawC3Nqkgb2adpLnDK6DnYRxTal3YqS3ta1WuysZDyNajuxd1o
qefggXp1RBPfA6XZrZAWD3cTPcScokzUsi6M5OA7pfv8Ufp00CrfLqiggAYFuSwkYYo7hGME9qBQ
0M+IJyQRgrmis/D6pCaJ6M6eKtKB3Al9hXvWpQLvG8HRZnrtwDIDggOGwcpcsiFqlQzMbyPePNAJ
1q7XhllJT46NbYFH1IO8eslTsbgiT3ZStShmr/Ce86y6b05X7d1Z7bAl48mRPeWtWmG/IX0eijs8
xOnQygKFeQXSoAxYKRju8YNcDDrdcRy/NJTWkxU5xZQAjDKECCBTm940xY8pkMPsIyhVWdP7I/CP
5Y15HtlVcv9XP5l3fFIhi6KpHnvBRcDR0JxRu9BGoP2UVKcrmTVlyN7kY9yG7yKXabBCRKtjHFmQ
eyL22WCIMxOYr99BXc457TgFAVpMFFQeY3676i49fYhobqo9z/XD+Iz6JDegLTbT84xFS6YuKrFt
ULOjUDaX5zW9k4kfWDBd29vnmoZtHSUjyLgRUd163wzTsNYp5MS2widQPjwR+92zhV8CAE4vo/XF
TFq/C/kmc/eBgepGE90kc7Ube/BnvhHOqiyM5N0DEFLdZDUPBPrsJ1784DNs225fOM/w4WV6bO7k
1B2cmx9UKTCEGJfNdRxOO+Wh4vrGpEAE/fFiUHSkByO2cFkMyMx9eX0v7UguEAebqepmSl8FTCXu
sTYdklPHRw5I4NUliA4CMFtPx8wzkAQifCTW77AtbQLiJSKQP2jkG5GbsV5g4+RkYkPdXl0I7oHT
kCuJJbilPmL4ca/upX+YDrxNjh3jlKfBKJTlcadm1Sa+sWEM/uh0bimLNklJYInjy8uZcjF09hKk
rLWezsO60B0zlApAW5SmL7qEgf1KftgReP7SfZeMLX0bzKf5nafcoLK3R6z8JX2349OQyFfd9INi
ke/7RsCoYufiwXZadWYx9DWVhF/WogjK70zVZiH1fWdbtDwCROLmXVsBKZvIcXAA7FkZCsDdXxKn
Nv/HgjzJwTPS6N+JUvlYtw+mW+aEmqHVPYzH70IDgyjXJlGlhOSZkx7ablBdEsNreuu99vQ86tTu
vx2p9rXraFECRGCUXFUklbmnWxXgoek8Y6NTamIxpZckUjCE5FN6NHjd5VBrRsjCggc69oJ9J/AX
5JmpPfF1RofwrpblEZu76J0zCtZE4tN5ywml0MTV4KcvDSGTgrdZjw7QOJC3IorVPCpSwWnwhJEn
P5L9Z0qxayO+311DjkcWI7OiBEkmODSiJKFQnHmJO4ueeyjxMwQKyZOaVCzdBdR+oiIdlMmfBHji
lZLDzxxUkgl8sUS6YTKhC5VPWfFTH+HssgjKK2bUDiwqkUedsw1WwVvQJC6XWqvxF2uTPteetqNL
3fk14kr/rRACeCjBZuIVQO6GMooOCPHncILmPKaPHSCePn/0FacEgQUXkmvD5AVcBJyxopzZbqXD
j15U1o1vaS5DF6fw/NXvxAvbhzqRX2Mia9KvxPWDPLwdDAkWuRa+rs+brg4dlY6V/Agh+5kz/iOR
QO0oyaKZfPYnFULMMvt1QJJtmdFLJg1u42eZme++sFU2rdhJoplUOQ8QcmGZ9ANhFAseUY/l3kpa
xNA3rBrxZW1qUNMScFR9vCL99ut6MjudLloVjpkMzTaklHmUwwA5KDxgm00QZF7h7bGSA5DnZILQ
ewrnARtB138dtTBAbVoYhF5suR6rnvXvLY/pTBiYHnmtA4nTSIcKkTMVn8eqvFolHydgCoQy3Vcb
ujcBmg6Ge4mokPJAtfF5FWE54yhPNB1Fu51alUmTwxH4uV0bGdA4xJC1UbvcimXlP6ix72OdefCV
ZA0kX40NXXCIc7BjDX2MYwb5/cEVcWTOckbHrsHaXr+DT9pMWjxZqJHvr7vYgYcwOZFXea7P+3EH
1Y9tBctGIqKlGltck0JX0PK+w37XaLLgu3shBcJayD/YFmet/qaV3dUpNPtr8nC6PKzAtTyDKh52
8CjiMF9MPdu40n6CgO8qe+fy07kqkVY6+NWDkgD4Bh0IXCa8N99jm6dCrE8mqPTq4q5vmQM8eaLd
hdcW4v1OdxNVvuePDBvSAbLDYiUj6WNRXPnXFJ7fbptgIs3RId5BYgn4OafQOkv4LTeM74xMvcQv
8qXu+2PIk2YusDmKYYZcIlrp5E6aUN58VbkVzdj1zAvsXcngZL/dm43bvADPew4kD1xkRv+jKXHV
GmuZCWGfUCWG07zzuKYlZiIsvu1TiLwHfYG1qXdck1xOYBbWpq7+83xYehFJNGQ4xxnOMqx9d3CU
JQbyFt+nib0xBXVr1NgWPzw/3HmRvJoBpuqVCooRREroBzqOI0EfZLyyp07sGjtng53yuIz7gP9E
H1R+R8ENRkwfkMbCebhGc3MdsoIQmWCaz1GsTlryZvLkmJkjHbWfKVlbUpHK2KeaLgfcKXtMqVm8
WWydnZ3+Cr8p9KyT9LfafoIfv1PTBusMPuyT2KBDW3cD4yna0OE0HiSa3AKh0h4UpjTjcDbZcqAT
JY8xBZl0C5+AzDLkGh81bPsw0zjPxYiw2esrXOPnNmoFktZfUA3kPfTLlg/dsMCbJtW0e+LTlGUL
svD5O7G226TLJdwTFrKJXdURiPCtUmiRpV2YfpCUZ/LkErctXR67spGxNZ9ecZgibpsL3nGza24f
R1B1zH34VbIaLDNtDh6v+YWE0VCyqqpnQl+ZsxRqtbu1zPCe1hMnYv+ExmyArCCnFyQvMYF5AX8W
jtQ79jR5TpzSd491/bJhcRg+9G+D3JqeguFwvKMUVrIfA9HelavsEOyiOWRBF38aVl+EnVERK9Ue
+iketTtq/lUM0tIrZ5K74zlvqRJIIytdc7TwUMSz7KnEAt7FhVvIBv6W6KL6+GAI+ztmKKesyzUq
2ZHPBH4fRxw9aPhn72fxhkc1w1ZDl6FHPzNIEoUj35BwNrSLG7Sv/M1M+y6iRQkW6hkpJFAz96xD
L3UEb/Z1jl3KwACY88Ps6GsAby8rN+YIEwerz867rXe3weyLuME6bW6NkHHTQah7o48KJzFLs+4U
EnasUcp1ZfIu7eI/+gYuCsgZw6dstZaWkGdwtLh6781yEKQAWGWDdP8+C09LfPzhBxUXB+svjjqr
pjCI4HtM1TQtM9qNVj6dzOx/pYzY4w74akx3wMKZ5IhdkX+4+CmbdXv94i6GzkRV59qmq+aQRALg
Vd62HKovMzT/cfdYOVJjcpa8YtTn8XheOz4M8Lnt7FxBIUSKSPWzVLLOerXyl9R676g2w68Mmyu4
mp4JnjSroZ+Rao1+tEqU4MA7QgCnTcTc3q83xjd5jFtdLW8AuzuFVJnUaYMKQ6IdPxd0gkOkiz9L
aYYB3U0T5vQ/JE40hYRO1JHYVH8J0bxSLBGMaF4bUbTN83W+YobBOMto3PK8jgz6RgVDRedb5OZ/
BfLaQf+2W/ZlXHPR+LzcOeWddL8hJR41KGOrDSmofGLB7ZkFF/TpAV7CZdEM21tYEbI/Vu8PbED1
ZZ3SwOSspgwMbQFWyG1Vk2kzMdt9ZKPGWh5sqOHcQAk4jt9cEzGI5jsv1Dqt9hGnWAjKI9MN65f+
73c/FUQax4NZPCY37r8+DVMdb0K4CSh1Db9HQQSZw62hfe6cj9oWkzlYAFRmb5/psnl05ZH+g0Gc
jYuZUZHEGti/63FH01s+C+lZUk6BkN66kTQYVxmVqnDKDA7uqkITBSni0xFlcPE/hTPgRzulQxjj
O13ofcX7bJw4F6YWRf66T7mNUeDFjFOkI8elk0yPVRwcnyHVvc4EFd4oHKyY1V9Qqt1VbsUFBPPk
HrIz8AUgr1VVX5nuWCTwS6EzYjtlw2G1A5D2FZnbZHHipse2mhWbK+glNFrALC9ElQikKIbLG1tj
iKTPjiwNcuTeLwq6V6OLWOydCAZKZ1rOqKO1ugg4MezsmnxXFQ1EOgqV25CCATKgujhRdT15b4+V
Xl+gC3HpJlkpB8WaGXVGL9q2VX8blGmraKg3YNU+u+cy9aV41IEXu8OUoY9pVnMdRgUVOxY1FexM
aTqDfJIuGjZNcrBfTV8zv2+toE34PvD9YisGbKfRXdRibuTguwAo2vpGyQIi4ZfLZwiqyM7PkxAE
G3ELlX7eDyYMHRGBRonyClqAJnUBLfOjEB/AoQhAMQp7TwQE+KBfo9MsxRPONdu7I+NFJA2fpCgS
OZMR3mlBaC9VeiX8BwamivWByw9nnTibfgwtU/FdMfzkCwQHPc9darTSonBRpq3uWxcs06Djz5pX
n8hLciT/tYSWJ1Z9W5CHxQ5CisAWfKJDCni5YaR/wgdyM9y0CJNjRop3kXgXmYWhTqavhQJtBohp
0N2NGniK/cAeL/jqCaGHRDMhdYkNkvGzExme47isaEPa9Fhlnrty6Q8qfhnbVYcZYQkyc7XfH/l5
/zEGTNzxgzBSYL6VpBWXJmx/uySkOLPa2au8hh+y6dGVOmcP1FFxO3NvCRDTHXwt76qs86GpgFLY
J+Vm2SkzNjuEjHiFstFJ8LsxACz/vlQ0q80pnA8Rmm3xUEmADibpGv+ZVM+43Lxo/DTf1iGNOLX3
BeTe50hSXUy5+eyLaor19k9twHQKdzHh3esfRoo094ounXH6mcdlKZpt7krAlxeaRCvkQn2zRonj
TIFJSTmvPeXSpNUHRq/FC79VYiuhU8hKkR/qgaYAbTPwibHA17GmQHc/9ukvbXMqq8SeLGenRtjB
LfVqOGrf0ZIPPhcVxt5/ZvFSpHY5vOIRzF2fBrcnE+2ni+FKOuh5v4nAXQ6lVIsolXaVnbKReppV
jS+leT3cHqHdb1Z8xz2d4N5qqFtaTf1akU/x/AOllYWb8RdYfsRpvpz30zdceqI9vhrboEeN88BP
k2VF69jX9q1l7/ZsvCH2TteCfS0VcJL1IgPxNZkCFECuvBNpSah1WjSaHhRn8ho3TNial6nkiUHc
Sq+LBTrRqr653n32aqw4R9BLdOHXiim29iKAqQ316JstsfVjssHOTNewiAyYoDf8aLk6HSjmJZmz
yUZddIshnBPfiEKnYUQNNpEOP3WwgEI8ea/Fgvp/JWlXMH1awuDXM6uNMmZh14TRisRZsEJyPgdT
AtH3dk1AF1GfyUotVr24Tg8uLgnxywMcPiNmFJeKi2LdusI4XUx1JeiUVPVVZB9PDJ+fvlDi4XXg
PJTRVK+Js3r2fN3Pyb0g5JfuMOouUp/MyWLAN7N6SbOsd84mpYMQq9VEH52hNNJkTzVL2Tm/8RSp
jt412E2PAPDQZpyE1dDkCiBnZs9HCKanKaiziplFBDciHLIofsmzidTIZzkgqtrslO4l+3wg11Ay
5ZsapqgiRSlklv+5KNyB6av9yX3ShDBaHt94odXYorQkm5SeCJtmDhhyNQty3p9t3xfwB3k3VstM
0uUjWMF6IapQyU5A9/je+U4D8HAJX6HSFUYKbmclJcjKS18NcCE6nejbC/qX8pkmqFCLof2g8qLG
tqe3bnfNQRPlE08T2uLI1juRlVMM2yYbwL7HV9NzyldpPRe780N+CL2WtiOklRxeVo92TThSLsnP
e55gzKzMa+NBX4uON2lLXEtkGT5mSW6kH34pne15qZn4p8HtoVEuJprTBdHIr13/LDrcEfmSyDE0
FXYUCRu/s5e7McawZCorMlrXiuvR1q15Hpiz28EaJmL1Mbc/YwqYIw56FIaMGMNIxfdFARNg2QTV
1MFdT+J31Kiuc8iAiWym0kn/7UAaaRP2pBhFZd8EJpfdR6JjdIsdCFwDhzqH5bneGNRadwB/eC6w
EV+I80uRXFMVvWaYlngtz53Bms0tsMGzbxZBawPBSwMYjWz6FZuKQryYAwl0+N9MbhXwkPk81iXY
TEMJd3RIueSZRcB/3Au2phGM1a/iN0BO0BFKmobbZsK9uv5w3Pb2KSQ+RG1MOKFzo8KZPEs/hQjS
UqV8L90cCKujg3LmgG/Bb3Fk5PszrW9ANdoV6jZuA4xhgpLUwlZd1716QWnRnQ5/pOkTYnIhA+Wj
jvDc5hk6Khc9jN+FqJP9poV1b3C39p4xQxjwcdgzO8bH1yEwDftDcbZ470l0lZb/DiaGXOHjWIJH
4i1UbQISfgetdzISj/gEBqgg0t4Oxksh+xQaalRsEr7wMRjMtb8fGiumxKX0/gPBfglTheMsaKDs
FxFpGA/5Jk0Oa+EKdql1+1BRD6Nx3B8paD+0FviXoLNIldZOGJqQcIWkmihsXpWI5vZjgzNNIhNL
rCTFyRJvOpw+l9q2VYR5pX5hQZZk8E9mH2fEVqoDpJoUGY2qwCs7cJblErfgD4/qcoitCFSplMxk
1NIE8T41eYwdjK66LnIow7SxRBpjsK66jNntnuuqQTvZ/7yF/6V4PdDPcLwePpiycMozYFmnQywC
rFVyLztRgkm81H7SfeIEv6Wl0MwtKUWw4mXjO7mdS1qSJc3iLqxleKok0X7PmJU6lF61UEA55v35
kT1SEwRtKON4SlYM6O+NFBWEXuNCqtJmZ+CCDHCr2y3dPbf8V+rulT3gvR1mf2X8Gd2C27ojc15X
O/cZJy4ASQrpD4Pj80fSuuo0I0z2DwRhCrgM89pl8wk377YiSedvRTlKSHnGujaYnd4ncg5rrUW3
7JIOqeWbZ+a7Ij7nC6mnYtU6qrGx7nk9AKOEX/1GN94tA3G4HJ5/hRhkqx8fX/KGmT/Cg0+3NYE6
0fvoi8XbofqSuNRG0VW3oi4aZNcAQQX7xoK/qddEE/1BpNmye12VCXfbH7+QG5ITxSP/C7+SA6cw
TsQiOvu3Z8Mvk1UuzuN87ao7VLQPCpKNpIxBZcjDCpu8MGmzKy4Ptsi0PpjVOQikqnWvC0jSsuX3
nvNk7SngL6tKY90Qf92RzxqVgkLv1To25+K0WzjMNaYx4aibPMReGN2Q2gQcWb9ozKj31Zn3Dbwi
Wcjo/hw28allth9DdpEHvDK2Bzr71z7GQsBPM3qMHp43QxfzYON2jZQAA8ePDXe7plXAEJvRKTTk
XQuKvkMHQtg5rLTEfULFJtC3Do3mgvmBcI7i/n+J5GWIzrnhpJk+anCTssobi1G4WLMyQv+X5sJu
mzD0XXYlJCPaHXUnZnwezCquLy17UCe65B3+aSDegbpV5Z3S2igLnWJbOSi53JosjiNH6rYISDTG
CLbNgZ40WOniVUjMYZQScjlqdqAuh9JLU/RZqbm3i+3W9Sryr/1fy6flO2EkrcZwFamDNohvnnKe
/FekvkOTD5dsyFM0hq5HLrk56tq1D24HTcdeUXkHabVCehnRG5L+uRQKARRLbeHGcL7aP/5LvJr6
pK5hjbhXgiz9J/b1aOamr970zC182RSFaPrBLKi6g8X0sc3H8cv+hXKaOUDEYwAVBSapwM7JJ5o1
AXaZUIHSXxX63AbnqbREzp4819RzZM0h/TqhFLLDgxRpYdbh2TRsAlPzpMexkgoPep3Fd9XzkDdA
33pUTy+HcFepWqOPfJLDnkrlCavALOYiqSW/dhiwr/s96XDxG6Pv/tCbMkUMSgfKO2GE2dMsFGNR
TQ5/xIv/nBmSF/gicCheV4BnlFdd3bQqbBHP2NPIM9FAXudGKtOmQdxRHcY/5MOLAUzL85IUJqj8
s9MhLv2rwwnx0tt8k74bAfR2/ps/NDau3pjqCHpWkCXhrjyuBYz52f7yAU+FIRdlX2fVU8fVDijQ
8efUACasIkXRfNmaYyQzBvJo3goNgPsKl062otHDKYVJ1iSJVRTps1LDYxfeZQOyypkXoOeckSz8
htGizFaDFd26EsCo8aYkKZp5AxVbRtTnN9x0PXumQ4ScLmP3CEtUB86f92+weLHHX9WiNZ4RJMFE
8OuBK860LeOo3kDfr17Uy/JMT9gaBxB6xnUh3sfTJab2IaAXxUHm8m7wglUNy5xqHrJKlqEuEiuZ
tKh1QfmH5CxnISWdGSsUJkpRjRsyz/0oGG0rcvZGPsr2+0tiw0lBN8nLWjQxJiOOuD3LMMEFdO4a
xGc/aRVG7chPTsOaMYuPn5K6X9pfrPlJtCGw8FIv2P1EfWV+iUB0fWvV88Efs+9JrAF7lsvcnmUW
/78Sk8h4+mo6jArNoa2ta34DpFfT6/ZRZmFqXy2Tt2IrPahI7Ce5bVEVZAfBDCGLHRKFRMpehkgX
HDBAB7TIA3zef42MnNTefvktt59xpDTe6reRmyZ0SZK42BPXezSCpchCEGVaGQLlgYP8hgTHH2Vp
PP/gxUxEYPL7LOBwWKv0UqfZmU3dPyypu3RhZ+BYza6WFW2GRTOUiSp8VEN17qw4EAP4ixLwj2Tm
hv+ICysNupm4VpCDnfilQ2RjKAp0cWE/U/cgkF3sfJIm9Lhx8chw4ldVuwGIuc8b9hIGoui2Nbcz
VB59TzdI1JzpLHDtlJX7x3rhDmAL/YXxAJ+unYa6zztZn8SYv13Ky82/DutEhNMSzwx/NKoh0BBR
pfMvfp/2UdvVXQrNf//Tf79D+5VwKYqhhmT+wyCLGSuWAMS4KZaoQK4ETr030i5b6wcpmJMj+0pZ
YP0Zm3Nn/ZlnNW+XznVWWLva7Co1cpUiHOcK0W7wDDZ15N0ZxUqlcjDZuRfWfr8GdX/qTJuwsJVn
Z7oPO+JUcRozWAEe9jKON7XwXUG2aPblO+CRQZF/mXUOvDwkzuvbVaH2tEsZa5kenss53t78JnXR
ZiSVkWXwoX0QUSgSbswvjho6IkwheM7VGk9AEmuY28p+5DT9BHz1mMT4KkASQ/BxGRF0u5QNpzaT
QxG7wNW2HOXVNxvFCaYUxriGa6I4JjlZK+bYu2KRRZUdczTjfq8hnrQRj2I1PpFB8nKNsry0JMYr
t5EiapF4XRAigRqTnrFDISgRy7CC85UnrXfDyvzXMt7V5IK80jIINOI2d8mwoxI5x3Lpn4w2l+L6
UnfKLqV5IgXQqkw0Td7fF9Yzh15q88yFtIlKq5OHqVL66qzIYYNWHD/e6R5YIDmIsjgeJMnCf9CU
kXFXHxOcB2eoG2D1sUBY5sM2ELoLhKNoGCiPGAsrK5a70eiAmKsR0t9bx/5qViIO3KKAOZ0ndaTX
lR+a0r1M8vD3dKP1svvnV9x8F9hVOX486FEbzzFUjwMN+Do3rf/N4yIhEvmLQtB7T/oygMeHruin
NufYUbCYDT1cTmvkB01kbD+5c1BfxiqxxRrJTaWUHY/2vKyaLT0STYApBO+cOM3qq/+oVNf96f3Q
Z+0zYeX6XcwqUsbUH7FP8IaCBmYaDS51zeRC9jsRULQ+rGdJFz6rEwMVM/nJI9A0uqTSBRrlwjWd
QrCwlXmZnkEQR6RzB7R3WPFAKx+1dl2ylQmevXU1yXfJLH6V3I4rocNfIUfvwt7OonMd/W0dHQ6e
Rj79CZ36ZchrWNbux89Rh4JHFipmXXBgLuK4ejItE+Shpp4Nx4pFlzcRCIRVlMcNdl1DCd0PEYYp
E5LKXce+jNkZXnrp6tTWsvGTOlQnU/a51t6YGnG06XXUgqWjBAUN9lt1arAzLy0v1LTx3ffOlmc6
nLHwonyBR4upV0o8brFcam+6zQcEWDzVPHb4DGtpOksi9ab7OcF6MATc9UzvWe1fFveQTnH4AXXw
M/XmrMw7/rf7L5pYHxR8VIRPeSwrbt2cwVNbHNhf3mTinQJlaMfq0p0KGtVYlZ4x2dudkXqY+Jjp
zdGha1W2yBux/uV/KN/xydZS7rximunQS4WASeL9lGNLpRP4p5Q2TUOyglt21IonDUVLHAlT0YrS
aAMFHlHcwRIIVa1bdVdVmhZUL1kBSAzCgmQdjomOFU5GHMfNTUua45o3svsXcHUAgqdxxuSkSz3b
tq7g0uEJCQwg8oUmUGwM8MhsmZHZ07kEQ05214CGRxktdKUtjvKvXGahn70L3Ka7EHSYxFivfVR3
BMvn1a4qyyXHHQglxNnyp0DUPqqihE8W3jz7E9SNL07hN91+UBcZIkJPTSguplLy8/OTga2IruZ7
0u4baO1e8+iA99KJyMx2nJDEX6dF9Ny3s8dcZmL++Teo/r0kV+eSXUNbw9y7diwiT+FBPjwu0khI
kgGDlo3OSs7U09pr6SZuzyqeTGXeihGzZbkgoQKPR5YDET0TWV/MLn3YbifMex3arleyS8UDFfTw
4v/SeYeKW8inaMfI+V4pqs8LALGpzDt7mae1qryEXl6cKMO/+aw5sx8sNmAARxCrs0eeCBYQmSCq
UH7yFKkA2B15UdD4BRwyDVsXUVYei99OlhViwXBVKOw+6JT2zXMg6H1dfUyv7r6aNv3Hkj0teC0f
QMTKBn1R9vhZCAQwle6K3b2EXJchIMal93eOSVvoZoo1achS7AjrrBLs84ctIG2nFIoiQEPZjJep
vTgvetDya5S+L5P7tzskC1ug/q50K9LGfWboXrZoffrV+taQ5t5nJ5Oe+4iN2oC9sGLE76AMMiGc
HTRPaBxC2FyYAT+zvvScKGSMQSopQkA5luLrreaA86RcPKVtEHZm8I+YVzBAEEjDBXHV7ikJRx0Q
NLRCEVi6qeFe6+E6ESD2OWJrbFtHlNlDu6KN8mvNSVBWzbQMiivK9pHR5yq2FB9SapzOhxuonjag
Ga7uN4PenwZz/2pfLU5gnxLIGTrPXVPSymoiuuAaqffs+A8wwh+vvXG2es5On4yoYd3xbtprzCwy
2v0a4f2i7HXv6HQbs+eqkbI7k7/okxiN3W6ArNQ5YoH3Jk9PtwPEuc9vPwQ0QNlJE7X5d/yzCHTI
PXrgpmCV680vp2ycR8txLnu52Ccl3cgMZYjrmwF8ldAq6/zs6DRbJs4bFW/UkhP+ctkKfBcGdTwn
qlDUeS8MxCsLYKUgiO6kpyutazQQXmNVKtmEG7CWXJmxDgCdX8drorJvg0notQcoN0oh9ND+hArJ
jCTpwE26gvfRyHEEUyLbcaKGczb38EC4nx+gUpFKRqtWVRhymKgjk3j5vAWjycuHpQP0WqQWGUvF
UyoBeuPv3i8VZgFxn/vj2QokaxcDt6M+cSBquJdX89lzB64ScEtS8kFJCSg9IxkPBOM2rLLyvHSW
hf633bn83rc61eIHPFrXh8BjJj4RGyJ7TUr03XAPrVGRkgeMBPhaNEsH9uDcRTUMOv97Hs2oK8Lf
n5cAxNtqCli3QqCjT7U5sFaMxznZCr+X4DRyKwGEjg1q7WOsUO60yzdTXSTPKcsYMmbBsSoa+lvL
KNr8gsS0PMz6ZUbnwuc0mSeifvdM7L0xF4LbVlS3hIjsCfON7eHJO8w2AoyxEX+Jr00rwY3DRlN/
lUF6+IA65l8M/vPnwnHx71smKqQGTafxH24yPHEDMOgwMYr7mENfmr9txyFNOynJU+o4W1a87c/6
GOKPWrlCiApkwtwkSpba+A/se+QYqyj9xgirOEG2HETUqpwVFA4sjpGRcIMOLYoTDfrW5lvoSXkS
USFb/LIdpGo3yg3GsrfSzZ/z52Nj+MR3BFR3eNdC7H37MKf+twr+t1jY6scRfBU8kBJsWzbv9Ar7
9NeUJmllAyavufOuO0H/mXdOUeZnQm7DesdkOtycT5mbzIyTt5wdx87yvSUJZcZT7LfsOhPQqbUS
qjAUvpjBR2DGwm2Y/lZ0k7/wNE3e8JQE2tLEOFdg/A0okYugY7eJ7kzVTmgORETotnvvJB2tYMrG
M2odzsxxta3dLxPW5ORM5UvCBTWqDC26XAqwOsvca3mKjPTAEZ0XSKoeECC1WFSwMapTP6JScTas
P9mUJs8XMteGc8covbeO7/DA15xOiEKxFZBHEtj4I+F01ubB76JoFkpfqX63VE6He7EUGipJuYKC
w0AIvqUkfvjLQams44KUD8JliM+pjQy1BhjRebPjQLiEQNlR1+VknwlHz2GDV8H9xKq967b+cQfY
MUEOMpUNtCeZmk5ns1adgHbg+zEvSp65tZZ/jq+vuTatFzWlqZGvNQ6qtXn7QHvgieufR1RAQfnn
dHz8iqWKTcB7RjpezuRRq+c9u6nO9Pr4Tn+EErp8g0SK1b2ajOwdDSjpmip83r3TgA9C9bNxw1t1
/JHqT4YL7vHRQJO0RnuMvDvTeKobqI7OYm3JFxBsZz7JwCyx7IHeJsIdKJs1l9/qSXFtMvR5dxZS
l6rM9ZOtskhm4N4w4B7IZg1ELk+DBJgfKvSOwFfWLN8hKiDcK54Yaz2Kx3mEIdtyUP7G8PXNKYgo
Nd8tohNfXbfE4OXMpPykPqUweKfqwV+suCHmMe+UAVRHxzUeP3luwv36ky717ZdRW1ExyZNCt7vp
SRB41zu/Er5wEf2EL3zyCSL8lPg3yWhsljrvDodzkbYDlc2NWRcM+OJAOPbvBSOCHT84r+AL0rtt
+R1iCNYHlim6DbkFHbZ2OfQlCM9TQzlQAIYCUuqoY4V8P9sMr6vYNDizoSUO8+U76hrGQF/D7SaX
NyUvMabiHaQ6HFe9EItPGS/0aokd2Zgh2bQ1iECIEH1UcO+zcN9dViR6uiaqiEo6XogRPDoiefkl
pJjldwN0K08Bxi7ynzcAHuZEalJFRIwW78OEBFFly+UTcZtkmOMm/6AXe5blHA4TkO3VmQXUsEHO
t2Au+0nUaP1JsiaMIfWP2Jr/g+5lhxNN70biC7/9z5QZ1xMjQl1uNN/zlnMCT8qGc/EE3F1/CZes
HEHAAO6V1FDLs3Aly0X78s+yz/rh5j9afoGSJAAz3MAV6ajp8kFAVKLg0KMFVAQpNl0YMLsFd6Xt
gqEkHql5We/1bzMjNk86IxOIuhrM6I/74u7fA9Au60CZu0wIiYjEIcElkSOFwEF2BG6ZZ2+P4qMW
CTrOdgxFvghMbce+X7hlm/B5VqCLpbx8kgA607GicvRm3iAgND9lGqye6aHcKMzQEAGI8YW1tHdr
ILFhovLa/E06yeWe0fGUhrBOYWGhA5AvQ082phOH3RVarK0YADMZJ7brWCPNigEcjtaaJ7iw1zix
fob3LPpFMXWo+Gawv5JmXULx5E6xcRk7If4C7/64mJKUJSDTRjCarU/hjN8CGrUoevW/1oc1Og4R
UURyTWUKCCOcL0kEe2VZptfTJfgJv7NGjTXOGZTZSY3DIZej4q4eEH1C96/emPUvp49n6xtxcjJd
PVdM2H3akjTUt9YH0CByvd5F5Lzu2l4XRRDhl08QCzOWik8lT/4WiHV1zVBKzJoMiT7L/C6PQJNd
vRnGmkTnZKT83hPgTygXYyhb50xcbviW2AdiDeATl+H7a6+TfaxuJW+wEDLoVzF2SclNiB6s+1iv
3Qo4xpozqK99K/Z55QvwIatEF/3lYyMf5IG6ad3Fp2xl+E2KMUNstka8jeeszmIubL+Lnzu/Kwh7
nzaDfdBXcMRBhAIW3/0slpg6mcl8TbE1wFTIqTBTAzX5HH8qGCwTrJyK94sDJbsWO/t3l484l5ak
YFJPhAGS+6PtDt/8PipyFC+JudKwJ11XsBcBO80OFF1qolTPxkcF1q3M9UbQG+UXG1h53QqXDS48
ZfHOKsVHvavdxk+oG2udrZBlzB9M85WULpRk94vM9sy/DFZKx2TRRodZwztGQycpizuZWekTr8+i
tQEJnAGBMsXCmA/h1KWM9d8AprltLIzH09EiYIzRf/9BP1VxFKtk2knqcNSjz7jwW15rqIobPC8k
pYRFP1DpRg74cP3O8pTQo+3Gm0TE5dok/hPygn898eiGkFpEHy2Tov+oUgv+/SYgGmWxq+XlXhB9
AVSo30RVmH29U12elEVBK6NhozEStEtduZzDHHSC6A3fn9UctleR/JO7N/ixRKTDukuVCJBRODyZ
QRnI381fvp7H8aBGwclWnJVzIZfTDAH+evKgSpQ4eL8WuCcVwlnr5+YvYx7IGp2Ht9Rw8skeUalU
lyXLf6+Zr/mXB68kLRvXY94p6dYtq0KkWDyeE0ReuqksYipszexC7NBrYNCg8ZSPcz3W3kGOoNct
w6I8dR+dbS73X72ACZRY90Win163qeYNNWc5nrRitA1suvZ4adyqERsLPMEN2gFiASPukZQ2CLDZ
MjQ7t0naF6OXnBkEmfIZYQvpu7spjming6OkzJoAR2KlHzJX6Qt9JUkNjHvPPutPV/8nsLezemDL
ACWH/84acEhCGhlY3IvJb7VW2TdiWPlU7lwUyKSzl9PJe9Mh2QL1BaUPeZ1pfg2O7+ioTDjb2Ooq
rDlAtKrcAvhVi3XOFCmZbNJPdj4EkqW1EvZQ2HljZw1L6eXGEkhMYptIPc+PDtSn9GWregtZm00o
gb0BNoceLnci1VXXMes0O4PMBh88nKBBmT00V2YiYqKxRMI9rqyGIO5EkWuHQfxOWX/0z5K3oMFl
rbOOQswn7q1FZeZCWeix0BUrhvpFiKJIYohG3mjRZyohfmyI3bviM5rV69eoJ29YPVkrmtFAwGe+
Ni/Oturufpgi+4MSpAT2lY4SAU13fvItx/kH2BDNXzfnZ05O+Rs9IRUivgvnPTBBdY7R99eB/Nea
kumtGMAm5iaFPVBuPIqEQxuqLm5kCCI5/ozj+TUd7SNy826dse7qcxvV5HkvS9KXzmE+kvhmeV9Y
IWko12dnkdGyhio9VnndhcARbzZ9jWMsvDt+lrTrAxlaL975iymJ69D7EqCNrBJGm6LyyJH7wDg8
3a0XyXestKFhAaD6slVQqFYlCsodAOgi1DjAoq+OzUwpJDA7s+eZLXpK6S1pqOiR8+iY4kaLukqI
MwSi4WPFeefAOInjbQxmecoLAXU9a2QnkUHxs8JIbBoze7LWU8BMPZXuJ824R07VoOAS8Bt46LgZ
pttRLlnsCkjBzGJbQelwWzTjNeVm65cNAyFHKjau/bcQmxcvikUvX4Z4gbVNsd0v2MPn0whPNgav
o9rBuj+8g2ewZbiG63OKL/5aBdpkaQrNjbrSz8MAOSpegnbClL4xn2meyKvW2YToY3J1igoP5L2y
ja6U/o5CF1f+0ClXwnZ4TuTLnUMk3Lq2KqDcxCvuSM9vD+0vfPJZQFNIkiIFgW2koG08Ymd72q+X
NMZilteBL6tEmbYznCy8TLwb3ReXTYm/ivLs1gk4wItVBcXrbePfTi4vqc76vCgcfXdkx9hu7AC1
5TwjCLzLicoE8MuIH2OEGt5i20weP0VkFL4jd0Ly/L5c0ZtcgH5MuchLJkipxwg1tXQC6NC+JSg4
WB31gAJn5tEJJ//x5Y5kgSfgZ4Nq7biu2fbFaXMT0RUysksq3gt9Yq3fzO0SsceDZaWhBPLmyoxF
ivCuXcjzEdqCxGO/GoTGaT2AyCHSC+R9vGMWWJ6MsiBSONyv49WQLQROM+wDOa0tbaIgsG6SyhNh
j1PYL3MChjHKNqbWshZ1cuGOTtjjg4ffFn0spsWpOwoPWslO4Gte4Ge8QgXd6A+QRzB7pEILyeSo
lBHVUc9+1ZmmyAhLJPXRF1Pt/Dcjio3/zHP1vqItkuI+8CI+u+mkjQ4H36o2/Yxr7fvcbUzlpD2W
Zc1qrbUsOxtkusk4wLy+QCAJCGOCMW8i8Q5CAmE2S41pC6He+fmVL0EDEZc0LKt7sfffsP735WVu
aNKWXOZ6lCciQpqPSk0vcw7vcNUzJIw5yM7s9ozUstiNDrZztA372LgztqIQ7yIsoUNSVYWz00My
KFR00PiP17gWQCIFkagloFDKEVkUCG1fKe+fQfGL/vPJSgimQgGMZfGr27kI3zfSlPiG8EjJQODP
0svFL0BCqjE1jGzChEo3Pv4zrsLZ07EC/Pij2qMEbgOD2LwP6pw2LE9Y2NPkvvLOTV3M0jRnKE7X
jpGlLiB8/S09BIf7ECdHxsZFrSFOZ8xxkXvwxvNtsZ7atoMlVsW1hULhM+iRJooPLdkcm+JsUB0r
JC6KDOL4w5i9JGMHNMJEY1XI37mRW8Q8KxKloz76j3CV4tpSgI+kuKOFYmD+TJD2Qs4a8VSpeUZl
lnMYuMVJplJx/W5Xhy0cFmQkrZPTzXTUioluWnBwGCluCi4pRFvbjlJxoKI6WPLBZVbMX8XgBOhe
w7WSP8CSpkg669yzPiZs6PHufw7RSaq2a7TTorIBvUy+VC0AirMtRRrrQiRU7ql7XYlAVURLXWLu
cVxFNHNFG3kUvT2M6vt5hHtEVaqHaDB2+ziBAqwtdr6KoVeXJH1tdVGwlu+SXVcxiigilV5YmbSf
NC/rkdF0P+NFJvyor7zQaUg64jauYR8JHNI9G/1HxRyrw1ZXtYsLEIRvsXukd93CptQebLKve476
7n/FwdwHkhPeEp69msdnbX2CAHlIsB/xP1Bpu0z8cxLAHwufjaSYhVDzbsOv9zqopvjZ+zXJDPJr
69fHDljl6dbMwRIRNUZynv2TjmLSXApV9KrBzY20xZjgrkcG80fpSDzZpaoA45YTr7S1OI73Vprh
RgzFANRYKkIpF/eZSd2T1P8EHQ9jGLjxISOkgvpNGKcUkRxvWRpV6GhSsb87ky4Hk88NFdLzLlzR
jJ+vxe7bzs2aYxvVK94pGmxi/xXkq9CXT8XGtxXp/N84K82vXUNwQc45semzA3cNynqPc27JryNv
56XVhLTO7G4lxq4SJIRuCy/2BxURtBPU7cIv+i3lSo6NplThusK/T0dfySbizGZO3fHweIp51bnr
ZydvNW8aN92LKqb/IEuAff5dTTS++C0e9j5MmETckmDvtvPeGQjnPcEN5Xtk/v7FZ0KaC4XgGVxm
dkHTCm0VoW6H4TNf41amgOAt9Tgo7YxJk1XKtGRhwihqkQLjEGLItPROqxAkjape+huvrhkpkBan
xAUg62mambXy+a9fySVaRA3nPHgApZXG8391RwB/hpGSrts8kQqYxx7k4BjSDvufEkkK3okQDsY0
zSrr+VCxNhSw1Tdlk48evhXMgxQY5d3shGv5+KyM9omT7DzVYC7bJixx+OeuZrD89FU1L7JFuMuj
mifVJMuz2YRchO5VrpnGDtXdLnDQpMZS5j48Q+fMIS2RJ3p64pdU7NPH5FYQZQpHTmG6xl9Fe6+E
X0DOxXdI69S3oeoectN0XzTEbu1PPNwsNA0xVT6s6Z6dWg/w3XQ9pFNZ9XJtW7xwkOwD3/+d8uh+
nhlHUoJPTKkTnwxCuk+WDSJrp0ENECj9w+HIPMh4nZu3jEoe8hChpgX/zIb1A6mO9TYM35MzI/4/
eW78IWOCvMLdyGQUbCKnJmoUJrrQ0CU7A+t2u+Llq3rFFOF84YIkYqXwzIA59PHMd80s/vDS7ZCH
I9OPxvnPGwym+Xg/UTMFziFbY6ZpYmPa61Xv2FBDm0PP+kOHvXotbj55/BIKrxw2TQDoHZbARt28
v4SrDhg1KovSHfkCrAHTd0PwVJlAk0TlAa9YvYShsVosPTAjV13ETRiPdqWz8gRV+rPFGYM38+RP
DpZHijVmM7zLmgBHkIZHbean7pEpN2ARnhMWdvltFE/ntncoS8Moo3B5xROv/9GM6AbaX2MZoGl2
2LpCoUrkKTgzA5cmtJWcZ7WR7Ypj5tcdUGn37kPP2BeBBbwxoLpVnRTsOdPY3QgMkBdCHNObhLzt
E+RnigDW2DvHfktwm6GQAXdo71mJbIw2uysbc+pjrYWje88mlAAv1NSZ2jPVM9UBaDk+/QKAwVwd
FjEQ9zCiNmm/Qzh31pgiK2iymOKKYV8teNZv5KqYcsaEtOngjVIBa5irhZ16bGRoIc8ynP0cp1V9
6rP+g7n4GJBQNmJFw10+dbmNpa3SSXjuTQnJKXSJBMhar7g1RtteSSo2jqQmC3b8lDIfTEBFnKvP
jvV/lmC3iZczLYYtZ1mPSu9QQXcKHXwszNuY4zmhihuvFTjtN71WN5qfmKO8CSy9/vSSWTYhi8rV
ru+3p7wIJOF86aX2xSuJEDxRr2hvyGJEyuy90rYQ3tm1SCa2pmDN0YzG6qFeFV38+M4GboY4cvg/
Fhbi6v+IRbnRfYRx9jEoB7jC9yaYqjTdMPgHDsEkvveIBHmx+kodPMhp+63u2cC8xvu0L8EJ6dDd
gZXVZ9SKDH7d1ykqgxKYeoAuNQetlP7TZJT5eYymrqJBtdJjM7lfWCuMsWkKRzVSRP74NBr06jEQ
ocSl9CL83zkK1sKtUFtHbAiCisbqsgedNjsgteTW8tJjmOKZQM7cBRsA5NTuAolj0gyyDGHwo8Qz
4Z87cJ300idSalBGap0aduMWiClXa3uzN0+N0pjNAHyFoVT4+CdbxCNh5rJFIytafoom4hMmUlXc
tjZVEz69rNHgo3hKTNWvQ51XUoQG4pB36HO0hoq02u3y2AL+eGhYrlLsefHoU3JEAd3EMN4esKY+
ASTt8oln3tR1bi0Jw81GxM+RO1qsN/9aTW0l/5WGk1fnQfn3C8DX9QFZaOTROq9yjS3/KTKlhZO4
9bO3e2IQQvzKysCo1Wnfv/YoymK9mzpsz/qVFsT3y6IQRzpJ7mnBQbOFZk+2HlS2E8C2HsNWGSsp
7DCVl90F5riqiDTtfkpd0syCmxOzaVv8AqxTBV6ciHi6xymqXwe+B/ntTgtnA3OV5SBiB39w1YSL
Vkl2KoMkGYeELEUJkmNpAs0yGE4z11FQrCeVN7cqObAN/cdizVpejszhObtqM4cBnAtCG74tHyJT
GQYVvIH/dxbhJ2kZ69uKd+Bn+ufDuPj/96CFIHXUfs6XeO/G9JHk87kn2AovGT6ts86ctRpYl3Pl
w2Ft9Y/5gEHARYczxpNVXMp84vi7mqcNwHTIVrBmQbzgBmRpeLPuDkYQeqi/HOcNdWeYRfEv2pPI
Pi3zkbRyRQ87z2rXkYrYCiWmwcFbBeXSMPYFKFxewA+uwembk7k+rdybFvY+RmQtzR+/DRIywlCO
HS+7Kg5VlfdDZfwdiysWP8ahvyDWTxWhqN60GQy92YzvRwlMjue9m3JsFk35j1OVq4D/dYQIEW3f
cAwxLl/+JqhoCKjr2lvw6Y6pt8N/ZyLOtWb+pqGgTMHD4+EDWLOU5TPTlE7beilTF4RqMmb6iDpW
U+Fzfc0tUxlXMr/2N0EobzGWAER9s5oT/kQn5Nn1JH2yhwmSP8Z6zkcljo6O+uW5UAnXEHXky9qe
WSMFCOXEpRxm2Za0wAvlxU75SGaof2ljjGftI0744qP/bHS+IS6Ur6wUXSvos50te+a9l78eluvo
4vC5/wF4PSfqL37Qhu50AA0fB1T2/bBHGorR/pn/IZi73UEh030KGAPJHLbJ6yPZ4RaCpAVPaUZt
KVrDBlBwOftsrbdbS2qPxUq6hSejYBfkOnnfmBepyVuD4WUhsYifQswL9CzgNutdpZPQi/G5QoC7
uFf0TjR6N41Qx2jmVDRRyJnc59RMYIi7XeyPWg6wz0DScjEXm5XVkyagIDK+yGNVBWrShI3yRwVr
TF3sy+nozT/zKn8NeFJY35HjJ58yAaiTxWt/UptRQsJwejLqS8hngMIXlFNxgiFR4bt2AfBVFg3r
8boQRVndVFrn5s5v4dZgATtAYT9RM0hjC3u5+CHMN2+5lYD6Io6MRrxe6NXQ/Y09QGTToeHvPd4A
JsCIHmEA6kR4TjCnzXqaFszRBHlhCeem8Ixsk2moXI+au9s0VwRVkHbsodT93XYLDF647pAFeaOw
jqbN7Q8w3HtNVOz2jiN4H/4we/27jnxx7vab1yfhETMGrABLgahw2geNWsL/dC01dRQyhwbPxF75
8BObfA8LOi72/jjzm2OeWRLjSF9LFsslZFpmlvcfTWI712lfOdTl5qY0izvLc0XLLUpe84Ufqzl4
Hrood7PhE3/pZ0FzOc5w4/w6fC+XycwrH3lC+c8XLWT0hmdusOv5Bc7WQ/S/Wt7ZIJXK1Je7NwkY
MIKrgrUCNktUwOqEvgCOlPG/BZh2mi9G+czSsJn/IikV5SqGAZMF4DwVq1iTTZAKDzV0OGVeERcR
abSX9J66ShCRU6Vy6n5Bk+TohtQ3VtEBXK29l7zVDbwMKxE9B/MiFuYYbLiVc84X2BNlFmd74QFf
EPDZiF9l5gn/dwKzHMx4gSzUlsQ5m13v6TaZSbhk93l+teP3DfC+HxZz0CnLp0UkcqbWhE0IGJ0z
NnWQXd2ZjJgBxvxSEwI40afzGbbvfi7mE8gJJZy929pYkv5aFqvVLdSQV9cS518QzaJFbAKd5HOu
WjvfM44SuGmHKtmDqFOj2vd2bQBoWBSLP/UL0PZ7ySGv9qtBcaB6+IN9wXLMMBs6xT4kfsyiIdyo
BincrFw15BqiZMoKGWdBsEXxJDFTaZae1nIxkOyOzaNRe5TccU9qTJqH8CL8L0XRlKqh1gAtUYgf
ZD5f79A/zgTJRUT+TurgXfT8q5pfHqUfBc96NtPAuW0EIsJQaqgybFmI44TtLPkWi6zwZl5xCjGu
JmXUwEoo5GushkU0irs3yzhGd8bRQ4z3AsVJ86NkiTVXtmVkAIeexVM9DeZ0ksz4oeJZHbwdnskD
QQMl8N5BHssM2wWlIZ3wLlVoLycVuG9TT9A1NmWAkUB37fB65uVD8Od71HemrSPnLGBexggb3/YT
UocOC9zhR3kRVt8khxrHLoWwyy0Xbeqxtm1I23nvsxrf9Lk9UiU2htBlmCayVo5wrajqvNA3JmfB
2Vfgn3nE/cN3/66V8M2DQ4fCATbM05P1PW3gbKc8w/dEVO/LV596piCsNkK0Cjxg9VdY+ldqW0wD
ksyniZ/t9gtNLCamw1fmRvMbyfpX7i2AkuAjxOOgo9s0MjpMHgneRm6uXVFEez991y3bKwxS47rd
trbefA8yl4zMeOw8WoZDsQFeKX6S5vQ/i1ZyzwCSxw2oYy9H/hkGlxQyVKD8gfFHvMCdZm8smYiq
/ZYt9cTsnBComqVj2jLAZCBbcX+R0ZDvePkfX4Si5kd2ZJOezrcXonO9+sg9O1UGOVBnH38Phtxn
7aJh6XY9/vm+q3A5fdMWpirxAYwHfVrXT+AwA0vSqRjR8t5rn+gvf5VcXw8GXnYjpapV12IUxgEN
23B3MnK1+xp9SQbEe5ViCXKekqyVqwZ3oOSZA5+fmZagLoZBJeEsAwMdQMFTG1mq1EL6lznEFtJ3
GOHVpEnn8YYk4bHrdKvKbdjGJYXUo0r8G4tf62mEZ54OwRdMohaBhOwy1HHNP3QTfrIKzAJUzMAJ
5qARp1j1Wahf1m0kLkkVEAh829yJ88gJMriL3zI+lDc2+khfAbXZF4IZsAPJoQysllFV893UZBXR
dH311Aad4mG6uBdttFcpHhCuiMQjQ+eXzILM0FmVNs1MtqgQElzLCgQfnWPqKPRL/gDnWRxNcrFm
igut6j8/KXAi9JoAe+pNrUYOJTwWNgxz3TZi6UReycQm2QZb7ThA1dgukOxKj/0j/YljT1D6/beq
mwZjucDqJrZjX09LvQYFjDSABwk5yoJ7roa3iA9naHXKCSWd8UMlqbvO/6VpAUtYozzsbO4sfzFW
A02Jx3/sK1dbwXYpHGPRVVWr3piV8oSR58U3ZCUuqI7hsGAxopliE5wMXxA1rxUgaEX5MV2Bp/bk
Q2v1D/5kXNxLRz9mds32/yOytUh484Q9NxyvPVFJKvyhqh8zqSlF+xMkysVXo4PwTrqWObNaC7tq
YvQykyOYPlHC+I+NjMo1p1yE6LYOon9WPFUGQ/JHOg9qZ9GMLzU2PxYIgGdUmuLYV5FVINblNphj
pgiq9DaR02Ase3t+2i1BJLBWW3q5ZRApOetQUB7MTqUlNJCEVQOMbcTo5DNR7DL9+5q1+si4valb
D+mFvfCEhwMXm2J/R6+9sqbkEDTvedioZ1zpVjcDjzB5FSRAIUAZqT9nHsGvnaGNwX5j/nNSlkx8
R1KFkqdfUmx1ZYuiGtoA5ukS+eHLpNE73wrRMxk5Ng0frrfENDi2kOmRk4EZFhsNPuOeKyoGvcPT
JMDkqOCvNGQu+wVgHWMKASDBI4luUCPmdeg6Zr2xbZM6Wr1cWFDqSB99MTJ93O/0ZobCIb4FEJMe
5U3axN69QNjcqSHyoj0J1fAnpWky38DVkk7vb/If18QPhy5goqCa5fce0dZIAaAV5lxyGEGWR7fF
orEzCVKIv+iwz8O6O+ZXzAZh3qBk5G86F+8mawOD3gfv1ZhtdYSHon8KQuGIbLFjogfe/41Y5Eb4
ixDfsDqPFPUsPe/6gk8SP6Fo/4MNEh0gAYnBI5brvApZ4i1y35hs0bR567c+o6LWBJyzHAF5Sja1
i2OFG1o9jlTDG6IZNh2f4TpAN7rIqKJesCCDK69bLMRq4MQTKYSSje7rmLfy2fTi0ePKO43CgWAK
otrcMxBa/3sA9F41FHBT6yXNhruhIKi1MR4RMmeD+9FGZdC0Cc0y8rackou+FyXXUgPeUFW77af4
5seNrKaePKs2TSnlj4IufZX0GQO9GjW57GVJ9QQ1Y8qOvWE26GcOcgKKP177ezVYbhXfDV/aMHXI
APnH9GyFcT5hajmZinngrDzniMLFJQAT1lzYSSJ1r30oZqYPCG6Ki560RFOl0nN/QARzhh0y0tqT
AbRQzZHKuBb83BiGOeFlHuVk8fk79DrRG/Dhw9qN8fg4L2n1CHC3M7NyGvWLyzmG5YE3ed5MskGA
4BYv2oXbyUquMKDWDKyVs8X7ZSbWmleauG80kax2JZ4xPWIjQSqKdrzye3xn95wL4cCPodr5i3Po
aJlaEnKm/Ta18WnS8YtfO9A+/W3FOiBWUKI08p1B9qcxAlYPWsjWB0E1Abx6RzjCB9eXphK8Uy8d
namUME1JRqH8xO2iFiMevhrdKVigQlyiK2qo3mOXhxGVPqpe7r/CRwXPKeZIHzF3sIK9zhddAL3X
BXA1dDFzQA5lQia0HctD0ROO5k6dmZIIgJNlqsBWddmEcVYhOYTWw/chS/vogM8i9kR+FgRyFC6u
MF6WeeDk9DXmJgvGgTETTKTZJlHQch1nqgXQKcOEnE4lcW9DdVAPDChcy9RoMGZFldv/XVQqWdxh
OlVy9sYDNtp5qEeoOPGfj19mKfsKXHVFqfUPQI7b1lenyEFTIub3zupccXM/PNmJdf3McG1xemIV
BRDRt/G7NBJDQrRJQBcIFrsi9N5jQNbHAupfNdBz4o+6ZecR/+w+JwYE3rgXSDf12xrXSp3WSgYV
uAsVVx45s3dtAe/1tJOePtbVs+omTk52KjXTDQru/xw5CFidjm+I5QZaJfHQ2Bdopz+ejXoH9nez
pKPotu+esozXisb8SrrkKfrKNjuUN3O6Nj24t33Oc464VSxItw3UVk0da73p5Rx045El9hOkq+x1
ST0/COy10myS8U24e4QhUAzr5F0eULzhVeB79uLb5SmdGlur0Bj0aW3frsBNyxkVhMWLF2BLB8ae
EBatZ0Hy2ztLHl5qT4BcohtZtIoepLYd/eFjv+WbAn2zgHKsLdSJayFnwMcY4rQD3BF22GB4nRRL
7mO14um4XRzf0z9zLmNPVRHx6yCLKB+pcpYAqT5ApZmcLbpIQ8zCHeevQVgY8QUOXMKgAFnmNHZt
t+q2s9yFi/tVVRZCVyWK/FGg6IMW3Anza0VBm3f7jLy/8rrjWv+HpMbN/ZQ3wf2IPl2/WDOPwhqr
k6OukvxPtiKZzdFB8eHPVqcB9aBqlG2dTD9wDUwygEP2hqccouv3mkTq98MjXTGb+n1Qx7W0z0H3
IqilgfH8TH1RD5g9nB717zH34QajrKcm17eMaRT3/FF7se5+S2t2u9UYbk17mU5jv/zBRR+si5lL
jXrYaAt7oR0cu2wtfW6ADT4S21l0qlMDZD7QkbecMYGAVBmsGQRL0ZRZXlZL15mM4kc5YhrgtFun
W38qZ1IfcVm2Em5pu7UD4/PLiBHbvcYCHRZVbsjJWnrhTczXRsYzW+mSWpaFsskPEzVAoQxMCkX7
4Jr/D7w68CdYttcb1mgxdhYMhTF6wj8ALvM7GM22SGh0NO+3UmBsW8LPN7ObkIQ+v1LISu3xrdCG
d6eXNq49X4zbnqn5cr9CDTJUJsU48TFgdyqF5cCFiDjBiT/i4Vt3lPO2zVYviMZpObe+pB+h55dE
+v9b/phPsXwc3VQ615Xsn2comciL4ZvTzI4Vv7vqnmOGgBtdRSz/0GMoaoI6Hxrq8WHmnUyWBTWy
OnT1RlFf/zPbGmbb9RwpUNPDxJ16TFM8RLIk8vP6qm9ZH36Qi2CuSJ0A/tv+mV58Vfwa9qAzUixg
6U9wc211ifG4tb63OzPi1XYSTVDpdqrmC6UOgojnS8jX2i24Kx1ey1gOweqhWXa4VJhrQLJS6InX
TC8dAzg1x4sBAMyXIbXe2FGhn3B+8/GTZWBKjnplqgH9Px6+ni4GiMQ1q9UnMbbrSvIKUd8ABg46
PzB6dR9cOlDQ8QKh80XEkDkoIIR3lpIOtsx4v3pZnyizaAEaBzG4+TH+R/mQi1/KNXuqIgp8qv6A
AHeNGyIO59nX2rWEkqUbxVkSfstnt21OWkY1CExgPrSFKARLdW/NBpvrwv1j+wUzrx9k+lssyI3s
mkDUjKUf1SGvaBszKtUE4XOwmMbBoE3RC8PQdTG+OKUQT9y+YDb9rb/OQeSo7ePCLw3tj8VQd5+r
Ks/n0DFnm4vQit4PEGoh4nsHBt1rlQDvQtKNn8Al1KlHac9Arw/XCSgSlm2St27H2qXKAQvo64Iz
0IlTPk2FqBZ9dvACdRO+eUzzMeznu/rj45vtS/lHh/D8JYxUFggvtwPgcY+3RwoRD7kympeFOQz/
VLc4yUc8Da0a6eJ35mHAnsPlFwfDLtcuX2DE1FdLPLh9A75V9N7xFzIqV7QnMxxc9KUTEnx0P+Fu
XJXOAXlsBBfzHU1C1omj9VhtR7aSNj1qOtL3V+ShWTrV7CTDqkjr3FdfgBo1LxnwnaXEKIc0soXo
0uEnR32GNaSgP9ObA+t1+Pyj67gIak+HsArt0eqkrcig24S0JolTQ3d1Wvgx0ORDiLo57yu/FRap
ZsTojuAbd59S/k9bGKsP99oqPet6vWbIgnCKmVqUtjVWnikE6U3o1xLw1BJCzv+Vg0+HTIvtgTzC
X04N3lJOmWUXH1Im/SR56JofujH/4uDjLtlQcrPWFuDP89RCA+18MapTiW2UJzVh8f/9nqAUJUkd
4/HTa3XX5UBMT8zwfbYjORDZSjb7k1QOh7mizpQBd833rdcHLtlU7jDGoK6NZTkc9eHJRGHczlzn
9WW/I1M1/uSTVfkf2vsNiyrY35oSUCv5dNByQ/HxdxScTZwtTBRclTMpDvn/JjC5HTL2vLNM+mz+
rw6VBDdBEfwZY/pSpo+ailycjYOE3dy83rXmJxQ6vG2n16LrEE42e7qA5ozqVzh0vSlrxAjLIBlr
F3SWYwyr83xaU9/ImsrQwhqqIV+45sCSQAclf+f5OB46WUIubAcox55/qR7buqRg/DT/kBH6FtfX
jQDlLrDZIty75Z6sdLlyfqoWkDRrKFYnYQc4mr+/KRslYig0gKHXRjS8w7HAeBhgydH/IVhWMvau
im2goTtJnJ1MEZaAgvYJWwcaCqdVdYimaocGeBc9DS8LtHa0gwn6ChqDj2+w78pYyZsFhzqKMH+k
ftNojC9Es4BYT4tEbz+TH2t/nSZQWXHNppiStX5V94AyW8pqLcgi6Yfu4yWbxwShftGiP4BN/dhM
P2z9Hx289ZdawBQL5uEz3ttHZ5bU8kLd/mO5p+Rm7U/a+G6t2GSDCzFR61eD+BaIL3p+7W4R8etQ
MbdaaQaYI9NBIoMHJ2VzuTO2l+QZMYcIw3/80kysKx3yKRbkcxOf9gBybeNN5SJUZerMWZbbzK+z
vRl7TPmr89fffBdgtOS2TAOW/tHMptLRSIcVUk23z4BShEXzxKJA5xSp8pPodi9Df6jDsdWqJXYr
1sVRBfbK9WNnE+xxatA7bCcJ9bK9PBMLfAKM25dmT3NffY+j3s2XTVQC9e4PHLiLKooYdJZb+r7H
EI7JGLa342Vlsm7S4LtbmQ9bprX5t6LoBNt/3tFm3Bcxvdn02IlrbufmqBNWgoUN4Ql7NRm1Qf2j
+gJg1OwKhcpkrpfFTXDVrHRpWfDUgsS6Eu4kaIo4COCUac4cCFkNO9NlzmWoH69ypm0QCsvxYk3U
sdM243PRyj7+HJPBNzhnk0YlahdB3f2CqHYO9dKL/XD5QIyO/5ZoGAT85pyBYt2mUx+NZeELf4jj
wDjbA3w3cQJg6GkxgMMQE+WKza5d9zz3AiiC178QjQQwh6YcpRCt2RfzbTI4ezQM4Z1qw2USSWZX
IW7Iz/evDQRGwQxeujS/PATzdBOx+IMA6erWPONyG3eBPOANxWQMJ6w7zYBWeQQHV81I7TC4kL6x
tI0o06ur5+19kQRvubxtUixv3BU9NVj6ilX4u76zDcyHZUQOfWTd1KQkLrXuo8joZun+fFF22C9r
Sz8J9V8wv1xDavp1g8k9hPQvOIIjWLUk98L4RvmqHaOaXK6urT0UuUds9P66Cyi3ym8n471XUB4H
OPM7kqV9hFqG78hUnImgynRHoiuMSvypQstdjniBUSp/XsTtI0i1hFuJVkPz7F8JqfyJRiDQbmG5
W8eOOo/JfMkAQhKjz5mSHBtK4aQby1+3UJOHVq9Pj41Ts4Eh7oHPzwfNJ5h9+z5ODDcrb0lFR2nB
bRE1XNW5kETBTUWD1chewg+kQCTEDCY82s51gdoVZVtR0oj2+ra0uH6+UmwoKK7Zfvh9C7PZKeiP
tKEdgJ2h1+n7Ggdusbo73iLjWq1JmJ3CYK0gzgVmsvp/2KrBsX3xAk+PUX4fVmn/nCWqFrHkXR2s
PEZIRdgu6RZw0LvzbHsvv7vHCP9iI2L9dx80OVawmDlzIcqgusffgOPU8WEvSOtv5zYVdxdNG+Jo
NAOjfNMRk966NNpFLEjqDfGby+DS5m9HyctdyEl1P/t+m2T6eOvR/buJH3BNmokSajUjK70R/z/I
FObj+9mrnTJ1XWvk6aQ8ld915wHo4aB3voz+d21t00InUzAmMEVPxichcY9E36Pc0eOFtlUMKVp2
rTZT3DrBxqNNQPVMVnIt83kKSsQs4HYfm9fmd7h0nnDiGwVtlh7GD3JI7uUsf4xNtMpi0N6q6PXw
yu++BHhZCBN0pfmmb8kTiAJmrWLwxk+yXj5HHWMQMsRz9IdwJYyYQs7QPPwAO6iCc0ec5MnLZDrk
atTeypNafr1+swyJGqxlkRRUDTXiMpSWH4hB/JfnApGaxdkNCHySkuZkPghONzTe9hElzKEIHESm
XLQ4CA+zPK02z3Uw4noUaabKzrl5BwT9aCyNXMxNW3OiseDRq801O3nJs1w4RqNl0bGBmeA/tGFG
4wgAUiM95Kbt7PZheO+nuO5ZwaNv2nz9BbqFVNSJ+veoG5I9eXDkS3ADz64Pn9gFeq5xP03vRIYM
YLy3KzXOyfkQSHjKGv9bd4L1fekBtEHGAJWA9y+sOS21VkgU1Kh793nks14bgzu0sff2YuuetTz9
VGHZ4xNeuWJD8p6ZIlXPTSgQPws7LKn3rwomDXbgPHoQuyZC0MlmXqPf+tvIbSBkdrnLDMFnYJF7
7cl2d6GRRGTJeVNy6JaYzEJevIW1JqOXQ27OdbQBgWm3zXKAJJX6BP4T8R6gUliKkioHj9Exk4E5
UrcRgcVq6K16gNQp6lj1QxfA+C8BxOr0dDTEWs7yY02SnrK7ALm9lqoTkEN9DqGv60c4dvBlF4Bu
b2GPAfSwbfLNjloovunvO9UaV+6hDNr7W5jsFGQNdO15yrZNI2LLdEHeMDPMC4Xzc6rUeS9qFRwv
5xKZoYCaKNA7pCW+LCQ7A3FScjT4W3YpORpFOt6tFPqOR/EwcHxzLMPYV4dIod5QAjd49iVK+X4c
WSjMpWNmtTpbq0K/VPId5f8UbcI/uGsaSqgNTZbQMHSgzXmlCsckUhCIPqSR5wBK13TCGP/UUNFB
aoJw5U5DSyoN7Gzkp2xh3kvQ/lwdSeWT+mnhRv3JPVGLLDe6IiwcPSdfLjvHF069Y66N6MH9QwIZ
Qc3djVLGLfaMnPea2KJHEnES/gXnO0N9oh+iOXCa6sZ32Ot0+30prMimXAbchQ1+u6gr2rQiNylC
9wQHg2KqzhZIKnZzAnTV/FO+0HtXswlwsR+v09g+ZKyttIok4jqEwh/Y9R5zpnTRldcA10vdbE7O
iW0n/8PJl5r1CRUxWdi8rQaFJ+ui4r63Nu2l7wNwbGEAQ6NfMqZkqonEoNomfleuxJpyILQk022w
AsLi5ml8gm0tHLRSDzgiLoB+7KRpVNTV6loHITcCJGFIosxmxJAInj8bydtnkjF34h0M4ABc5aBz
Wut2lT47m8acVNivCPEktLpYuxopTT+rTIK7W6NjQ+kPsjGn+FTH1cwMES9a/5rT8LUteraql7+u
iQBXULeA/WL263aFtEqfA5d9RqXGUlMkf83WQNuA+RvkrWTt0mKgcQdqFzZTb0OjiEOuztG8pnoo
UWzYVkcMV09o4pfEGjWEpl720gIW+n/4AVAQNVTdvZx/BL97/0HrhlbOvRun3Ja6UUNkqiVF6Z+f
i54osX0vQexs5nAjug0zVWxw/c842eHzsEbuNAwwTtwxXdk5H7cZfkR5G0XFvseIFnBPU1dD1Dj+
Sr2JBF7s7PFAefjSFD4M3kUgsbBpa1v4V/t1w2mqYQs8S1HjyurA3aeB1CFnDfr41D+JAgxpHt1N
t8M/oNSvJYVRfbYuZM+6ElUR6AObeZ/vt4u7HUEc0iQmZzency60DhMvvhQeDVE0eJodml+9pIbs
JQTEitK5wfGbClf9op5+8MzaNkYRHTRvZJ2IwlgQw/X3x5x0uC60clIIyFor0D2lTcBqn0/IFhOS
orYKuiu2XWwQwg6e3Ccix7jR5tHHevXPU0UX7rHQGtqL4ifHJua/ArMRMSOgizLIS22nFDoAdfUh
OTbgt6YcIix/LXUk6mlLTyCqKR3zy3Gy+Z1FpgMYJhl6PCee4C7qr8rDjxBs/BMQa/ZYtnXVSdMF
29HmovcQmHB2vD6/MzybrR4PLcq/2hOskZYY94KOZSOiwjv7MHo1IDiAd8+tToFWD1OJvkErB2oO
jdkQSVdIsSs02rL2nzKBjcoyfIHw2BhEPM4f8+MdUxiRR/v6IMxnmvlCBz/qDNCnycuvqfcti1rC
tTmUIRocf3AUDtREMgDz7YPYLKc1Mo5f9iTNYX7YB6tTY4NG7cN+u5dIe3tdJv42Vd/JSvj+0MSK
mwPZpU2zXfw1ONh3+CqQEGhNZNXFhSrKz86QQIUMJyN2jGRvw7tgpYpjarmaaS8fNjMVTVCd+hft
191rzU2lVGmavAJkrPphFQOT3Z88/+tmnxO+/iN8fzDxGN16YsG1cOX82lrTglgxK2DlI81Hy2lH
11dbXBauEpVVEf0n1SxPCFYFyBZZE8vAs2ZTzKEZZ+/rK9l1m/92X7e77RdJYkvcgthi2cp68E10
/QnhS3A1nXag/dHj+pOpGYdr6rX3afz3xDI+LAGu8TKnu6/K1zJxzrt8mjRcRaYW8zu00AfeHpIs
EDMvfCOLmOVOQRo55nyXG7uFo76av0zzNXmSHvx8l75CNq95ab9eM8oW4zIzuP7L3f/eYno4uVGg
ThPYvYsVEe42BGRq1AIGJLTYMjj5cKMX7WByt5B0zAllICBwA9E5PpYN+4Oo97kjaNE6Tz23+2sM
iYAOdD4NnNglVCmuAXpGGroZ6KMiW1HC5yP7olbX3xiUasQT0LuihUEE/ppRpW2mGxL5PKHRNN+U
Z5GWyufi9fgG07wLaF1ImGuLZZTxFBSWsX3BiHHT+07Aco96CoTbfuRJj/qRBYSTGk6dI0t4vmXO
oYhzQh2Yx9oeK0AvmSQDUiAFrfJt16GadmvvasZImJO4ESI5swoKcc4OieyB4qcH8dBMBjbJcJQx
hCLK02LYHcv/nbQVj3Hj0MieN9Na+Oqcc9NObI06jKkaGRKMMnb5Y+2g65SroWIM22vmXTOu/ORq
zXz8yr4jzsMYOXbPOel9Nu5RsgyYQJwvJ6it2EJCLeBxxiF7rLo8BZe1RsvfFY++J/CMSXCwnKPd
LGTMwIGVgC1N5LPsz7TQrhjwNfo2fVchyzYl0fSzt8YFqlpa1OdNznAzrHZp1Ai8VDHefbD9+Krr
3UpMnSAz6j89AOTuLUT59GN7gbOHtTeVieCrKeFS80079WVw5T71Ukhhzw69qy/CavtAQMUofmKq
6WMSmTff+2+jW6o9m24CwwUuxY40O55w0Yv6/H47dm6xATHtrKcK3OyuPXw8UFCAREykoV2EYw/b
tU5xUZQZkJDRbX73hmsQ50fBm7SKUCzSQYs/BmN7o7ypuDa2WA5/a9Y8l2zheBMTAZQ48R6xKOkX
DR/wjEeFxTu8qHf/liXVTBD/OY0oig9FWi7kw/Q3WA6QV0f3fPuUyGOJ8R7DX6qWjF9Dwc72nSE4
enGP3KOzmU1rJFBmQnTJexu24czD0mlBNl0dRGpWjMS6csQ7d0dOB5p+ed3VghnlFaKhDve4OXas
ed3c5HwiNHSAo8klNqy5zsMTukwNPOmWsNDuQYo9ie2+IOcENJBxqaz2lFBH8agWhgIfcx9GSFd4
F5z4xpccng4kviEB4XKSYINvNHkpSoHSjib3/qJssbu5vmBJJqqcXn78VBDgUQ1+lidfvaWMybea
c9CvMTvSftcieyQdp+JLK6ihdZpMKqOkx2PIKYUTXBWQyns21kAPoaQvvD2c1BkJ3Q/uYZ7HZNj/
30yLlFlXDp4u/SnGK/0YNkRwM86mhRF0VmVB7bMU/q83f/WiNms+mzrp8TeRqbIKzCHznflDXPjQ
n20a/gPtklRISJUZn6NPmxrXTGMIqt9nsGI54Ck86dVjfdhywBkAp/NvKW1M1KTvKC1WXiPCOeQk
4uR5vOS235KMqARfcBHN9bRqht8vuLYK8RMNMOuVAYtHniNMEoO4sIG1+B9vHgPcj8FYbhZSe3PK
MNUJzsKQAKdAQmZLoJ9cSSv6wWXJRYtXRrrNCwz8nQSjke9YlG6d+e0Cbe/YzafTcby/VxjGtiE3
a/FVYid2YunriG2l8ndmxECxXXHGgpuBnWdjGjrNpMlvTjIKP4jEclRmzH2eWYSRYJKXN0xKeGGE
F1psemwJbCAXPIDw9S85QP7GHUATq+uzdqZ2SawbVCZGaD1tgPfVmvBSSo1oWgo3Q+ibUJD99o/N
qplgkTLlKJmGCOnyFdPdNXj4ClEHmpgn0inmt7+y40dwWVProB+JVqwmIO+Lms7VB1kXL01/dm6B
2z4NURdYEIOVKXgfJpO/F1RU4TtGWBRAz3CZdZNxebPGQlrHCGHUb4rjB5RLDLfva8QVrYBoFSJn
DVHtI30m0x+a3UTQ4kcfh8HeF3Ow1bmyIBveECdXw1LgtZlIquWJp8zK9eH+U//X2C21QRYMIgv5
p2d20f/bphknYdmlHLYQvE3iqNKQeb2jqhyXYxUCdxC2CmAqZ/lA9FMlpTTL16uwShacQoCWN57I
MyVUaFb6E5TRET6pm27nhF0vhIfBK2fpeVpRq/YEZzuBo4w2aYcHwajigN+LATizq4Axp9xWrc8h
LmMqbVaCpmHh8gzilI2PocimqmnjUnzRZ4PGzKW3uklTUnhNot4fekJofuzyor49Jc2/UUXqj7Yh
qq0NaV8NQElS6ZygJMGw3SIfwpjsOcRIVX1ikrjMoZ7uJo4a+2xEv1eqKdL1xmqZKTnIjwOWuZwZ
3tHP7eP4n89uMIDpoAgQrxz1SEIwHY90nRHk+bGaRTAk/9g47QbrifWWrRqZWKErdsRUPRohwztI
PwObx7+yPR00YjzCrASjqKDGwDtXeVeyMKGy/XV3XvXK9OflcvFYoTQVvMz8Xn0cSLcwzi6VYBt/
Q3NRR30zylh3tdM2UdHr9G5uE0A/DEwE6NeUzcsjQlYcBh8B3XTT5lvhDFak1NO10gU0Hc5nzZnv
Efj3ItrE4KUjLtvbwcO2DZkSUIw4MGI1fepRNG7ZD8NGVEi1QLBiNNl+xPvev752P1PhVIRijR26
u8vD7htA2rQsV4JkDbscACo/7x1D9dbQyiubSLbc0KQ7vvDNJZNscpiPjb7TuzTJUP/4OPjk+TrU
49KnhvbAvVvSvm0LfpRnO3Gmudqhcp2QnKt45SrLCMWq/peaI6PBrsouyPuo2mIKrFNW5kuoHLry
if2raJuhYx3xyJ3iLYr0bH/SMcrI5wUJpWL6XszYyMt+J8htpEG+TAC0UGGA4CUo6+de3+Wz41kx
/T83bylpISe/z09hHB0ZAsJNNM/xxNLrUmZyzXtV8G2YXo+l8XsKPEPlR3vDr1Y5U828OJKgJ/4B
XX8Equk/UHxgromgLD6vgIRl2r/gbb0FYzdiVecKJEnnWw1C8pHDNSdkG7AqUnMPnkwEmVpven21
/NAMYqJ9QrXvo6P2vYj5x8I0xCjZZ7fQx09k974UNgZcXsQipk89gX86KRR0zAZ8jkd8l/ov4eby
fK/Jnen/BPmtHynKPgRKEpVO4OYVNJLTOAQ87kAtLlS8Wnqpie1n+r9zf1fi50zZshKAVPoUrbb/
MspZf4FoCuXRWcivZrAjEvrGEfx87pKu1HtxoRD41dWCnV+flGA3p7Pyae/l+OSbfq1jf4em2m+x
BV5tb7e0yGSS7BWuOR3WFRJbLJuy3SMu/yDL5FB4rCiLG98pitVE/UgbSwqB29JrmUT0P87bfxB4
RvPw/s9JcRFVilrEmree0wWvLf6VIbZ0unsU+xhOBfH2TGA5BjWJRsSuh2mN+On5Koq0e8q+Wt/d
XIKQeMYnRqCEgQKmam+l6ougMZbGHQXPML1FvXUj/kvtL4EHZvAWiNUn00CQFu+115oL+4proilY
piP9R0tbcA6oUgvyMUnQuRAyKwUUwPSMBECusm6aWWLqGa9LZRsnYU4wo4zf0sJZcI/ODLSmZzZi
oTSh5gbJeW4NjLs1OYVHaJtfpcYplmPsHVvTIEsyY/yYbouRbFes6g/xTWXVa0vtQMpql/rKCVbc
Wmmy/F1vuPurmDuYrq6jqydYdPizQQ5RXKD86pInf0MufcBf1G5fv+tFgO0fVxVeyHt/6NCs38BF
kjOD58pB4MjBnJVLAEs3aM9d2PVLoHHnuDZq/gocITJI9ccdbF1EKkmdpqJb4rRLoErTRJNQ6q5r
yhXtZtb0wEf4wPeJ1gEAuEfIwdLlbNsrh1/tGZOUaXv6e6iNvzNASiTYEFTZfvG8631TzYOuwMZ/
mJ/dv9tNRcBEHd1pchkB7R6yumHTNQg5NLmVxqIpgcEwf3dWATEgWPgkGX3bWly17x6tP2Aud3Gz
UaMHAGOgSS2YX0z1d1hYc5wFK5D1XBSdh/31Eu/t7gGtUcNYOc7zSRDVR4dFZ3GgtXmRSdTJP0yc
ayrmvJ06lO1sKh7R9mcaUQLybsTmCaid7eFidlwDgja8ZE9s1sVpAipfgebXtF1S7WW7aYEB76qa
m4C33+eFo8L2nQc3AIE5V6ZAjOk20HJzX9E0J8wzP3K8ELDPEtET5eEFh20k9OwpgWF/nqIyEOwS
WGcOAxBSd8RUD50ZL/rwt9t+KXvFo+CQU/CdA/jWF/lKH0cW2lhk1XxhVbSOyRHuJxr8W7QBSKMY
vBNaNOVsKerkzFUJJ6Q/9JjG/hhIZTN46j/wuanybFAeqoiBvJBTF/8w9CdcvmiM9TLPz+6+q/wW
kklZ8JAVWenJC0R4wcaPzdqndzowxhqwfr8JAMdeAfksE42/P97bAOOeUxPkh6BqWhg4XB+4cdeg
SBwxBn0ll3T07XdGpCLYQY/ABuOb1JXVENw8lnwInq8bB4jH+46/fkeIgj4yhxLXDDFwrqGDilJ0
iyp3MDYJeS2rA99XNonGmjEE2C46j/XIgIe8/NzS2Im/Zjw0iWDbhwp6+sGtEt8gUD0ZRPXvT3Zp
Bzi2p/oOO6eo028hQiTInnetO2ieQx0yg/kpXyGjLjyEwKvPhV5iDwEMXdkhSYWmbHKVoKnOLc6A
DnmI85/HMjq/bLx0WGyF8Mx11H0omiX+Gtc1rSfarW/xYQmJKPWfPqR5f/Mw3p3cNDEzCQaTAsnB
Ve5WDQZL9ttJUXh8MzsphnihUD/pABefB1O64+ct++AeyRbgAocLfa8yOmxD8unnxo4CaD4pWgRu
5YaalbIOuTBrKyzyx9vE//9TXS52s7R6WzXNjrCl3PPmNUbvfsn+W+2FzwF7j9KNoE2TGfPAGAle
jYdsDgK/SoeOPMiO3vWlme/+WrcvmusGFMVmLOtF83UzpbiljyKyz+KC4q62kKJHObKH48y7xaxp
Bqp8zuv5EMoQ8bmO6rbs6xdFzbvYlAZE9zfYIdDZWa+goBL6MufqEkHcsgmfBCcF11ig6/eAhKoS
T76/vaTvMpusFQp6Sgdkdmsmzb799Iwc27PCrGe1/6mXglr/AuotJM/0vccrY5hNIwmgQvWfwwFG
7U/poEhZSYAvgcpNEbcAzBoZJrKbrVhCTB1FTI+ab4NEaOw4yO+k5zkp0vXFNrpr08sGIS6vw8wW
Nbs0wb8n2P/e/hG2Ll4+askG8sOLejMSAyJPU0q3+qQzaUv69MywRwm4HWSNYxSyOS4X9qIXfI+1
7nQN5tbahi79dtgHFgQK6L5ei5oXMQ8yAS4WCSsXvuqrmBrPRU+PK1cd9jxJGGO+lA+vmCfbEUJP
uj+nrchSXB/vRcxbGVVcxGjyz9pmVlAOevGUN8Sb4H6K8l+hRnpkpwlachYtglegfEAZy6SUzHKg
6g9A1VitBpB33IsOhz3G0QfWdJzdzClL5qPguia6atLft8+mVDA7T7VnxxohTDbp29pQpCy+2xrT
NA4DC2qn8bYyWmMQnWHUdZ1bJbvNTHSmSh7gCXZMJn71lrWKXOLrencT4CoE3Oy6ypJB3QmjnMFN
oVfUAzmFwFlzDc/rYBrfi2vQPMWkCC4HpmWz0XmI4IzN+heu6PwRN6+V27sXLLocKcfb8qctpIew
gFfMi9jh3NgBKW/fHzQsHMDJYWEIV37+YPkJMysDDrIKY/5lV5F16bTypHwCrWVqnzSZ4RpPRS4p
HFWn6RIOLBIjSzKq6xfEzGqGAZ3bVm1Er+TIDAQv44ItSTF+IuCh7IMx0LF8i/QZ+gVPW9oH3e8x
Q4bDua8UuUNDQ9bn1Rpa6v0Mpx8kpUNJGrqDZ3R4T57vgVP2CReDWtx25LwlB87VNoyga3BM9H0g
CAtDLBHCCnKKoQBj/wP5VyUHBh/4Iq1HVMXh+E/dTwm4ntU+cgdY64onjVXoz7R42VQ4rBTjpkMf
rRSOLOL3lxA19dLv5u60NnB8z0lCVp5PTmSSr7BJxD6/JlXT4Eo2zcruyZk8778czZ4gPTwz79fj
0xn2PQN7irMUXzEY1BYzdI/lLEiQRjZmwR9IGOcbEamX5NTcDGVGjEAaU8J8i2YQ1rOUVa2JjMND
pjDsjI0FUmUbX/IjRP+vRpJTWqqzjvW3dzFdS1u+8aQMeWPcWSmoqg9t4XTv4IHey+L8X18XmDUi
HnMQmqmbbbrhFgh3TBkPvQW5rfNgj76UpClEJHRv+naLWp/lJeWljdopcxfswSCTM3EvE7v4hX1L
QNBSQtL2BNwWexvunspUyJTGkBLLswkcae10vNA4uuJig1aqyqTWqqC1iDJ9vHs6KLozzHo+epdT
QkC1bN+l+v5+T3ZO+JwpDs8r45ZfUcPeBlKoHwaTDRiYF8G1H55j34v8GD2Qw3q3/xBfeZLWMxA3
DhKDMpW54Rs/9/zTvEnplnXfRDO3t5eZjXccy/B/nIaBIB7hQuPL6dkJGLQ94+ph3qjnDoPND41A
eOu+oX1bIBeFd8EXfbrCiuWFXeKnhMVgq9ZN/bTKnRyt0OYyucp9cBGxLIyuM1nNmVZDu/2znGrU
wDoMMI27B4B8ZUTkEKw+gJrRebz0WPdeNBjvBZc1/hfuW3NLyL9388zX94lwvXMK8MIuTjGS1y8R
/5FshocLxN5zPPhrHVUkdwUSDczm92C0WwYnYf1O5K0isC2tuLMXei2qeBveXvKTjWfx1HLs8Ybd
ErD1fy5tGaFzoBTFcGBHkyGskolmbc79Ys7wESMet9e1bNy/SB4dRKaI7k9GylLLAVsk6s2uR5ZK
dt+Wr8vlg4pJD72rsJ8GkdN575Y5k9GJHSpcL2gCFm3u5lR8RfSbB3tmWYTt4IUbVzKinHpU4w8G
Vpg+QzuEkxB2CyrbkaVOuGLzLzTqhmoR5BK1/JH4ZIF3KhCzJ7e+vcePL6C3C2W1DPQSSPLXUv0A
rIY6Jec2ftuMYajME6X2/fBdGqVVBLTbh3S5WO9+aYtkxDs5Nxia9VZfBtEVb85QLVMDyLHwG296
gBoSUk2vk7DzoCj5E3eI/vFqZ/7zXIuXi2fSzt0qV2NP4va13Vc/yw1PEW2o9g1f/8Rv3dzsUiO3
PJSuWgUEZ8Q0gK0hQjpieKgDQKXGfw8RYpG3CRZXexcixyq3JdpzRnhOihXSwB5wh+HwpwIMMOUZ
yKjBIGxuedkOupQWVFeZ6AV6pME55SlzuqeVr6ULl8JfHtHEL3UOLIORNH9+S7VUi+oBe+/RdDhP
0qRbSeIDkBL17r2FEiyN/eTPnqCDAZ8kaPqZKXAXgp6rEN0m0IYfNMLy8m6BCu/jj3K2EWFhU/b9
uCMJk4w4nVztIyVIRLVz5buhC+G0daYYws4+BHmpZbtMvKekFknVysnpUwYN6aYTLXtqx1xcJKFs
A38BTqRJSW4a4FRO8VqHef74BAaQcxYzDqkem4rtPQkg9VYK+6AHibyDg9R/YvFxSomDgo8mHIsE
IsAfbNWK8Podyejcf1qctDT8ETgvscbTGag4pRVCOfhkd+E5/hsXMQOVAZRzJfvuJ39sr7OfEJsv
vcaGiHzpaQmW/hhxEbUJz9BjRohEKFEXFQWchz6/sITgIye3e9Fgl9w+Y7M++y8qsx+pe2K2Cvoc
GgJcKb2BrX0lmufdwJrDZp4BxIFxy1Svm7UAPNZPpqzDx9PIq9i+O9yem6SCqDdytlmaYAU1V0uG
Ojrz8OxSpLW7gTI5mLmXRL9fvBHZLHTGVLCmd6AxHTsasW9Q+iiGo6AIcC2PZW/a7IFVNIjC07Bo
THZeeMrTbPiHbNMM1Y3+DgxnLmWS7ASmoGPhNwZ9mSWYbFlSb8dYiyetMzbVvqS45H3s/KkfXwZP
xYQAsNzyqJVhHpGcubGhYODB2wjihDls9P7VJ9Fu5XNsC2w3Pi0kgoDUutt5CxqOZKzWwl1AIiTh
fi4FpDc0laegmzh5e4UQT4IMrsGKLPx5cmENVhlMy+CH7YzIw9H7W2RFXBF4T0OyAwwrbpagmogv
K/oUoTx9zP3hxdxuCTtEPNhyTUy4MSr2fYiqJvGbQ6iGqssLe+Oj9j4vY3Bot+ZYLt9/0UYzIukS
AmQOWsuzn8qnsWJnvgq4d6zMastHBGSM0z/8kpgTM9smBYlrXdx0hohwWGPnM+BYcL9OiuWkHiR7
+8wUJc4v5vNlRQy7xvDU7Qns5bpJQIVU+/QY5Yke5F+m6mvTB/QgpxBNZ5p07zvjsQzeHWZ3a2g4
t4tGc72DdOBtyRdkdLBIjqq19BvF7ydkDhsLLcu0lEfzgkxCurndJrzroDN9lOK4wx1b8qZy+ABE
1n4tsqx3JgINq2a2pNeacwsQ8LaNep28jHZx9udwS5QIDwG5M8ZVA9YwbUlrPh/HZoWSSmjI4DE4
khX83fzFuVM9OUANPE+v08EAewsHepWvMFBRz5gvBe0k9p0hHLotiQZRX+10wOMYEPCybLvseUex
r9R1If9uwC+P2/ZRSSGHgnVxRzWJvt9+DWO5WtvW8/HnQuWAzZKR+nZy+k3vVhaJktiqiMrOWuDh
DnMeTY38sLGc1yIRvvC4R0c+dTqguBkhuq0PxxVARRITSXm8t9ZLmVH5FalrVjJqIlw0eQkEvqUT
LiFM70a6qPHh09tHngZLEG2g91iIQQOPqf9xC9L4s1ERtSqnrnm3O1/2/G8qIoTJd7Qn0TX30Oqr
9X/jaIr/9tm1gTrsgoJrkddf5CuVTLzi7xmx47ejII+j+KGXqvlnMk01ar+H7RhmzLql5wtMZh/A
BlFYPIXbzzkYWrKylegzHYHtlWZ+aVkdOkOnEQjE6srPAbV3nNXjhqV7JKUTpiTAIQdaiO30TxIq
a9Sf11WK0JeM5MxaA2aIcjShIn+ZkO6YLHwvVodE+awDSDIkBASXPu/0/q9izzjMlr6kcOK/znYu
xTf7dqKgj5/ZENWxHDih5B7qf8ZpYaF9usSIH8kqjOERJUJ+uyNjwmEaG9+DWDDPos1idcwU1Mcq
vnZGHxZIALujfrOmuNO/N4K+eSptv5lDc6+1IX4FYuDaFPDtXPCfUzim/rxu5qExIDeHlQmtaN0V
4JUsRbjuRFbFVtou73TO5GID1qquDBNxQItywV2mPMaUcKJOUxYQ8flg0zHFIahe1f1b/00PKXOZ
dSewgTj7F1BHUdDKGBIPVIU8U3FQx8GcM64Aqbq9gdNkpeo78N5wFSbN9BhHtA+GqNjrWGUY7gSI
51TERTsM9xw55SKDK+myISIZ0WQCbGromTbgpe62BFOPwcEYiEMI5S32CDg+3useckiBy+uzOZyA
cBF1vM3BJ8iGBAHxXUiF0MiKH4E8LiSgA+wAeIKJVPY7+/JQLNQTe7L17sby5/LcpXRAKTGjNvn+
j5hSHaJ0RKGqfj7zA1bvLwj2elTwUk5MrXaidkpwY8wDnFr4rJFFKzjq9eIvz9f7UXULB7k4oFXM
sZ2EVTjl2FprBlqwrHChbuCA9Mh0uQL7RXOHjK5hDbxqTektNr79ue0bQ9B4cBE03bsLGNbJk26Z
6PQL9ZL0D+4XFR9CPEZCptuNgudvNpAIBLnRvrJ4iV6ejFtXbC4ox18XFoqzLCENRSgZcDeumbDz
cArlYo8kFax9lewvNUSO9z1gJLzhCR9JZvxap9R/60beCQwYU6BpHQ/6m/M8LEhmmxhdKjMG+/AL
WFmbPsFEafIV+sOxcdRB9EksaSwPNh8RKbnxMtV/XZsvR5Ay6ZuZV0+g8zwN4X9IX1ylCbzNOAJe
F9xJfQaHkUQ+AlbDkJbbzmjT9PnLFo/EO1wty5qp+zsJbq9gTt/VFe52LpBB9Qx8imLNYhwl2p2G
snCmpAHeKirVeAEy0qXDE4PABndKSvxUVHgGyEnzchN/uXm7WC7fBx/1suPyFQAtASMMFBN4XSue
RhimdMCvilFmE8A/t1/jvDQIOqbuXLZJ6Pgvb9OFJtvUjOGlsHO8Hh/IjMjcB/yNSllN6+GFf9ka
AImMEj5sLWDNmIMyeOzArAo1e6+J+H72T00WoZ8fwm7S2Bi5zZBvF9YubY/1HJhTv3ekrvdiLVu3
F1zJalQcz7Ab2q1PKLkgPGRpsu9Z/aajD1OFIYVwg6jB0CQCdqCtI/6oD01vUTQTc/Pm/qA9RODf
CplB7164XqVDeZhkGbC/bFNkOq7ip3LclMCLkDxg2rqiBxicVzPtt//Dv/zQfDNO29r206qdypFq
I7WWbPc0VBpVrA4IdrkXRezEqKGommPUiVw0YshSNHgkNRuGdgaH8fnI+/Dun90QulqVT1Hsa2qv
iwdWNetOl2xIkN9NaIxxV+e2TX+v0WJztfLqtlRZgp//qtCyreMb3mcQ0KFrOAtnVWZ5tc6Lox1J
JqNDjasSSfPvKlxGrIePf5O1NJo9/97gFGD3vNIPSvLAofbUchXnI3Ip7y4lpqItpIG5JmlUODQ3
y7N4QxNrDpveJZwP/dZdV68L5105y05M3iX6/3IzOWp8EUHOjRCy4GOa7fuLZdpa/QAe3hIeMokL
nc7QAGiSoG+ECjcwTvWU0ZWG+2Z55jWoi2euw8NLFVuriF9p35SE/SRhNhTlCF5poFWJS6C6zvj7
+hFSMCmQckZy6GlmzW1BlrPrpPro4sHDyktnR0RLYSZ7bOPcPksQFHm1FkNuzhqxnMYKgLa7NFdV
AFTosmbKvoTTUWtsbu2Bbnh2HpmJUlixqnkQBEYZOzAH8YEavMbRLfoEd+plnY82Ne4y4OCcLbTg
bMI0Jvuazl66QgfVU9co1Z3i4FG0YPpVgjpCpYRjuyQKe+6s36iP8KHmvEbTXcsoVt+qf49q7gch
wALpvTf9ltdXGSL5SIsWgr3SI0SZ3YeDhlMTZDp2W9iatraMUYOSMCfObcK0vhr4a8KaR0Cia9AR
UGVUCiAAKNtDZDDHIDWaqR6WIkXtLLSwRYRE9UTGwJXGAnTD6RuNLiAPZVoggMaxU+F/HRwFsOb+
MG1f2wGWOZMCxb8VsUmcjlVzSqFQhJ8eoNn9BLawD+3TMFNsnGvm8kHSCQ1NgfyxGf4Y2fqXcG+P
jwSelxh4Hns0ktllo7TEyIA2x6Vshc9qCusvdOgQLplkZK2itvlhRZAyL/KSZa5LiShYvDC5gM5s
C3j7eHivnhz61IK/hp67BvE/rWFLMsDL46bvxmk/kh/oxSlos4BziNEMXPGH27PKVaIRX63HeR0R
cU7NIBnyNTmTg/JW4TpU63wLF/N+cGLuTf6zDdritFJAJQeaMqLQGkgvc3wH77tTjJmuvYmCCKZe
T8VgA43f7ANQ4tXGtT1GRAd1IeGnE+b7vPDm3xrKqBXu6r2Na1x15FiI3sYXYcBTN4F2E+q92cdA
QSJmlIHDK9U+nVDBlMWmimcatf/hChTT9b1Tuxu4XVODTmNhsegIYn2XGSXH110qqxGxORP+Htj0
HlNJZth6yszbs6hWqgI5PhyV07+h50L/kIL7TZXCdIUdOgNk2SlxQxM7vMDOxkHIU2pP75848Owb
nK2KOC+NQ97/Ru+5hn/etPiCauhho0se9eIQlsCtfGCtEDxUCaQKoCQeOmLtKOMHxbyG5iQOrXK7
GkcPnbvrLUPQolep68gOSfYJCHnbb5ijEKrgxheSh7JZYUz33ZssvneCaclX7qehIWJXaIZ2h3V/
eTJNA79vPuPvqnolUgbe8ZobuMPVfqR4F2LZsiYDoo6/fofwzSmvaCILnGZ2pHx8rmwheZTNJraB
Lj8ROrqcOkcGCPqy52i0poWMXNO1iwUoejBFHEw+qRLLKArIGT/bZTiAIJf8xJYWh59dsqBiXa4H
wfz/b8L6NKu/wtepKXWPa/PviOV3C5BGH/OiMa03JGMPdTV5mmC5Osepf8s0NmAgjImnc5tYh3lZ
wLyjzPMS87n1Cns0yXQt5otTc2CaVQyxuTYVnFCZZZl0ZzDdipCl6wF/vgxpff7QfYa6qSAC10LR
NQ/IMarD6XxmV1LMc/dJl+8qxia2NAOqYX12ULMtytUVdA1afY6cqACDyKpUlNmaFgCuJrHIt5CE
mwLCFcesMJZeDXBqiLhF6aotE5Ntezroky/uU8/RZqsrW9SI/wGznKGggOn7SJIXgwQ7b1cM6PZZ
+N3sxynCQc9xqJ6IIXZPS2pTe9RRv3kF17O9KDchkmfsahi0tfBKbTFLQwcRG/M8dakh37nhjBsB
6U7h3gRSXp/jOt3ifzfmJJP0O/AFD9cbcb6AqukEcTmmGkwDPPBRbfBRWHau2lFG7YKsFNbEu9De
abENtEXrmxa3eywrItjOsX8knXnkzlqAadUtnZOts+wHy9986FyMPryTPdhgE5Ph0cfw/ZnMHMnh
ewx0dD3qA+zSyiJputWamNmhz6ThXvPaVUbIGl0vgVksRCZaWpWeJLoVAu07gzBmb/acYHrK7SSh
SaQtj5D1wbdvBJz0ydNDWXXtPUJIGT9M2BNCLw1BaMLyDTsTJf4rBmImGpzW/DKRvFxUmDiznL5z
qE6DabXE8StwCqyqz7JMOUv3/rWz+DZ4qP0iOBMfqwGFeONKk4VHaW2eYeMGq097H28GkoIDKm8Q
N9zA2t1U/V84OkwFCqX+prxJaKb1gAGNk+RGIHUnTW5FEniuYb3aM60eXdqWKLAooXs7IskL8R/H
rgForFmxMCbI+Re0FMveo++Nw/E1x8LZJfkyn4KQAPVkmtopZ1s8ePM0o9ANNxAjv+jW2cU8HRbC
tRI71rZVp2FFANW1IHfqia5z2PlnUlu0TEU7xNo3UsdAW2rosjeGkUQ4B/X7CoZWq4tTC69DcSjd
NUJxt7SAfUOSAKQOmD/utog3xm4+0Przk3WIqDU8C8ef3D62yewsYIE/Ng33qr6EwXpDP111Sszx
cLCdwqgC6zWGi3Jxwt5pMIvZ0rVXfnoJGZzFdgN7RjMMXMKjQrBaevp/IGiI/KIBZk3ZDExlWY4e
AmsVwqtBwzT0fn6KDivAXevCQHT6MZNrkNHhRyMyEl3gx2S/gex7nmMFWtwcfhrzK0I/5u8gAxMj
9N5+IWC7UfCYLkL78QQvPFTdcGISPIfcqXEU4xoX1Ui5vy1XVUcQx3XswYgm8EBgd7eOVCJGQ34d
nezvGH6rcsG2EJP5PixJOkNJTPQ1l/Mclgr/3mlVNLDhskwJa6NtdmL/d9eEHxTm+yYE81tha/AK
XtGPd0+KZhCz37qXYnowWiP+xJOKNdR5L/z5u3920aB4KQxb31e3LVuTnWEgDgEtPfyc7oNo3kvv
EJTUtv+crhZ1WlJw/lwy0wB2FGqtT5Tb8Hu8pVluZF2UlDTfdjEyhAM/aXvsR0prkk7jDs9fGJKq
7OvkF3yRX1dBKiVt/+jiChIlALjdUp1OWWeY50xYcDV7BzAnH23TB831JIJ2tQDNNSfOc8A+HvX8
xzuvLXkSZBQjQxso8onNWDAHPX76FnZQK+tqF/Qu5b2TL1Q1q2yl4YG5kbazZc1CI60AmfP0ys+F
MKdETuT6AklLsFYVf9MHnC4+tCsAOYegO1ZVVH+T7lXD4PjG8+Y27ARvZUA0odBLXFBX1YJtY9La
ejFSUqbMQgIRyvBYw6uDd/gEOk+ccwM9NYo5Hls0bb3stDbOKJ9+/mc1NcMyQYSrrk4QLpGBlWez
FFMgu0ggnmNxDLYQ8d8Ed08Jb8JPH1BXyh107UoRB6uV40xlWFrfrvoN2tCDKMY9uUWLgGzU1P+H
ApiW8p2RjM+61QLHA9JEVdpflXYXNfxG6krCtbkTEOsNFEY9nqC+uBGg976Kgs149GqCAEFIpKYO
UbseP7xJBxvpgAkKpT7qqQDCNoVm8Th6311i62oKHbmqAzzmPPYmSgfGV+uH2fdJJAf8zSpscxF8
XSFWPS7FAOgmL8TWBlvUbE+7dx4M7NeKU+RQV4B2Rjm5fPbMgO5VZ4byL9p5RZkP1CN0F0QkPa0Q
BEaNwWxbbJ6wp1SvDKRk8fMwMbwfQpKec4kha/azTLH4kU3RSryY/3D1SnUH23qOBSP4YAaU6qT6
uSzP+Ecl5Npdt4Z8TCoamxt0EvciBDJ/hJi6ULi1dxxbVbryW/c4HrEIqhTCw+7A0c0Gf/oZhCMK
IHVcUuSdebpBM8WiazHhNIGyjxuW9/gExkpK6XtwUfJqRewO0JdfsfS95HmI758vY+rwfrJOsiAR
FfI+N+tpJFHiPGslQ/VGwmADPABVSmK7vTsmZi+DF7lGCXkS7PZdJVKgiD5BOvdxZ/OBZdsmwmY6
K6fYjm0jF68sEu5W7rkL1v4ML6ycl5X3oIhppFAfeE854D18W3h4Q2vyw5P7Bq5IO22aio7pw2qT
oiKj48c8oykR2gdDleTwJUcxHmtYe+gpP8/AWVMjxXHpFLMQocd4x52eLf1kzhrGTkGSiC6XVH61
yETEA6ODyjMwlDgt1/FUd1xAugb8GQNIzU3HN2yBToxEJb1mA9p6fyBaCFaWHlJg61OIZHyj/wxW
Z5BlAbklzmLHgG/6W1Jd9uOth05HMw1VBD2AwRr5StUVpI62nSvNaaTY8oSevaKrl6pktZIbCjiS
GL6A8cXJiFPZuc4VwfiAb+aBlp04ACSIHxpOV6/V/8xJK/hVVd10a3eVT7awhO2bCDgsMQKPS536
OfRdYIZTxDfVZx15aT6yOt7CIIZckzv2krxZpBYHOAMc+A90IU+lKWC3nr5K4BZOC9Kx8lD08J7d
/31A94roaDsAzD3ha5fa8bSjemLNUS7NwAKkolheFTfHlgyvrG5EQ6JQg4t4tGmedpbTPf2u0GwH
SVFnZ0Koqs6c87PT6GFbxWBr+BjTl9tivhZCAi5Kgpir45iNZmqvGaHjkHDwJ2O0GqDISJN/dhiR
rXuXyc/sNhTlEaC4z8c6byZhRKrS+g5IjAXB3oQZikWwba0xl2q/GVXs2x9u1jiUPq/zIRyrmMlv
0KC5p9AtXEtfLC0AQY5ZWZY29BO69p9VgC3k6T5j9OPLtX9b8mntQ7myAts3klb32G0FxOCIC+vw
1akTf9TlUZG4y3TzTwm/j4StEhuXG1Tgv2WBGQwnsVUxWEQ5O2QK817l/f4I6maJYKlGQVvgi1P4
1dNztCTtE+9KbhepIlF+TV5VDRhyMDyiqOWFPFTF5j15r49dlvH0ra96F+iXZU2SJwmH6jfkoyRn
DRUdoWmEVQ6QVOrbfqXnswiKGRLsIyEgStydRB11itsh7Trf8g6o9JeNTOLiqZHXVSylywLOGn4X
dsu8hbxTaM4q6eCokSMt60gru83P9k7tF1HvMXeMRHgCbpKnl/mUxw0CRnW0D71jaWxv2ZqzxwWF
yg/qHgL8xTyhWQr+3A+WXI903/rBut3MEJro6LtTQGNnbzHJ0CuQ/aOip0Dh0g2+sgg72A120rOx
nMPzqNhrf87EBN7SyWNagx5OHq7AfZq+6rWYHd/aVUhDLe0dbDSaH/dekrr+SBPM+jwhSJfb5hjL
AqfsYzH8GN93uA8HsVTrbDJsNlzkhbYvcj/ppxOd+ztlvBBr/51mHZ3SutbCVFp+ErPezrBKRXlN
DHwT8lmo71Hz1NiLS7O/dchD1SiOJuICgx/fUPP66DUrEtrmkG4hMLxD7o56o4pXPrjdfrf/t8wS
/oTZ0x8/O9b5vTnvn0dmPZ/PeOhhcSa7wz6oQoJq7w6U6gZTHUrVqj0+uQQr++Y4gx3HoNLkkpg5
TFFRZHdI/DWgLUnWdrY9g0IFFwQlRDFDuqsvARKjeT/INecfZYumED72cDekll0WxNse5BuMx2sf
dGqO56QBaK4FZvxK7bfCenhmbCD/+ijn6W45h91Z/CMPD/E0ZhWN0OqME/pDJmiH2RZOz/GvF0rh
FuCt6tCI3hFIdjV5sIMw8LGizmJByDWXdhtO4vgW1zM4Gh06IhvO8i1qyz/utRkF6wC8ICpNTpBV
Kv/HrcfJMJdARjH4baZk0xJJSFt/onMZvrc4/zp9wF8Ds0nEiRudz9OMeGPDJ1Kib9umfdE7QKPd
ltNf3zp9PoagvXDe5Sdm3uIv62e6bS4nSDQuXdOgDZMWc2fhSCE3t0BOur2ZRAaN10ii1+fkMe+g
6foR+vFQpgfVeSfUXXV7qubN9Mu72J5RI3h7ra/nIbeo+G+M41oN4MIelMWGoED8ou/IKHXANbg/
mQyfFyN5klhj5CLGxYLYf+2olgPF0n+BY7KQfZuZISw2tq4Qw5vfcRgbLz9Xk+FWIO5yJ+4Fcyca
Eqq3KPA6EfYHdH2GaSLoJhqihJ8n42bA+Sj0SOp11F7e6XoEo8H4PEz/JRfXizjmOHM8S+UT857Q
zUp8UN0H+94SvPj3f6v/GhgtoPpW11zRHndQvGKkCzYKb/hHKgbqVyXU3yrKvQKmrvfwQhnjTPni
75QOm3ioKhMYcY1Pj1ycYrWQzeBuj5y05cB6HNTYnJz9lgnmUAbXt7uh6nTjih4p03yURUFtQozV
eZVi5WPcjS0meAweFGRyGUXsgSJKG2PDYZn2WmPFIzanYco5Q4i2lMIHgL3gPDS/vbC6s0wb7QNH
7xAItCu0JHMLlsUrpKAmK0ieYjIYF4ptYyKKXmGVqwEtZAIu1kj31Bo54fsPmKQbipcKhX6iRVHd
2LT6qoJ3Gt0P1N6Q26M8sSSLIGH3PGGJg9L4ycQPsL9niwHYeI/sOg9b1U9GIf3L99XhdaJygNzN
dh6fRuiDUXtnzc4VaAsixfn48Ge7Exdl/BTKaB0IK8mVq8bsM5muKJKFk6P84T/1N3Sk/cLBbwJE
LrU+5YjiuPBTQ5rEtz1EV26pGnjE/PhVtcm/YQdc6ojfAbpknRgzhF2lv+r9Ykl07TxrsLufwrrg
aXAOki3Y4zzefxYFYyEqIu/vQ5jYUqSpDpjm5mpHRtigrd4JjRe/Z6JtXYSPARRuWD/9pxcX2SsF
H51mxFZ7V9UQYtJ/c06u8lkM5Yj3l1MFfT4BICjqGOf1XPi4jc0pJS7hLf0er+Bf0P/hZIJ6mkCq
5IUe7wjB75p8GsQ4LJvGeTx8ZnllWvQ5w4cy4S9XFrj+4Kl0UOHB9Tr/8FTJMyZHk+RYQaqxxPJq
pVnEiE9bqEmCE5TK9sK28YZH77GKCv40Lxwr1xwkDxd3eAWSEEezYP3/uHfjze5rRTXvtr4wC1hO
s2xZ8khxKgo+MWgDEsDs277XikJdC2jxbwL0QaCJSO2UkmXKq9R8+W3rR/A/F+qnENPfLAqBxcb8
qaf6mQKM2kGYvfN1QHXF9+aNgAbzTQQJ8hhdVxoeSUISCFQrvWMjqunZKUE2i0R0YlW80diEtH+F
nevUy+jY/rGw7GgWlVrKFHnRWF1nE2uqAcNIhN83prKS7ya8xbcK5e+eTWTgkP8MdtkmKAWCHVCX
HpmK8DoWgGlsWP6M6dzUqACH0LEuXSlI2YSXskZzGZrrXuGOXjtsbYklhH1lheWOud799TA53ftf
qmzag8AShARWlQ1V9wXCYg3/HYuL071WNw9H3sl9mD7URUPPI+UxZwjpwpCtBv74gFqPEzZCwdGz
SQdcIsRUsek5wkOhIZcTIkEQAj+h+qC1kQCmHk6R79zbRqUleYLZpbayOr4xwoSlorsffYWF2GFw
qZtbL5T1E5E31aVa11odFJdS5paxT2ZQtMrdkwh3f07W4goP1swLnlXlNeT/VUHR45hnA+kHLabq
8evV+R00VFZERLcrUoFiKWJC5hZ95yhilunlMZGeIlSQXfJZ1ylEZp6g598ZPvEd7WyxRFEw/kN7
iE9BwVeuM5ScjJ6z3yAe0eKPF2bMhsbxPIro2pVC7VLf/jAg6oZd+NBonf1FOH+mlOykbALN8bM3
05EdaFpJKnE5D9/y4dRMRPPdZ4MQ5af0dqKpR4CsAT+kxGMzM6b4Jqs/2JpllLvpQA7veKvl+IXJ
DlPPaA7CPS6O0FNCgEaCv1Ox98k7L35SUQRcgjZu04OwMm+0k7cNa+6nvVLzl1xrj/Ut026+Dl4L
fsygBswJfzET+mcihGp9KS2kvYomenAfHMmWysPyj0JryAn1CmEKbwkx1QYo0ckqlDZsoNc5wX4m
goqfhdTpOlq7Jniy07NZiqo6VrmMOj8b1rYOlMmeicqJWaiGs35HVO/g3s+LPuZxUBN6ITpGuqHg
Jd7+4DMUf62p2M3c+qUTJYyimp9mQOUsfC6Jv4AxYxZRRdtyeYJAmid0TrpjtdEn/4WK7zoEUMgW
vDtCSM/hgfkp7oEgxF7n1KfSpz5lJqd2n7/kpa2PXEwOHgd8jEb5ZqLV4WVzS4f8bknz5EHSyt/Y
tiwvVrgbyIlpdpEWzY5fGfCNwyNG/x4ivHAjjlTrXTNxSacCW4svw4HniCQx8SYTb1Vv2Ktbb1AX
TEabOW18CNyxjb6vcGav7Eici480jOGMimTDLelXyIIR+wRU7ks6qYKSbXMv+6zoalQwXEM2I8Ol
rgK36VMw3H98cD4i1v6dFEIgGl60GiXMjW2D1KsSlK3Umzohrl9xlcszApTY0LQD5rOjudbJDPf4
tRVb4324YabK4hCwi2wGC9+0RPJCpf1B0JwRrUgn4HIXOgEsbyVIAyrH9Xy5lAcTm0UQdDVJb9cu
J05lIwPYZvCsYRzy7Bdn8m9rFXf09N/9COOmDErybrrzO/FVQM3GvFhkxK6uS8yYa6QJpWoIdkv8
CJR1Yd1mlK9+KTv0Bqiump+zQvm5x8xq2Lg49hOwu3TpDskgUIelySQ8FmSE8I4N1taPnJ9Z1sOc
nbnzfyX7NUGuMABIUB15fzWpz+tRWCkp7sKstYIDsaDt+ZSk5aOBEaXUmRa1AQqfV/VynKbJKu4v
sEpii4+ZEFS310NAJJKvFq8WP2d8yCNSBNJT5VAcOD9sKZphEIt7eF7If8cQdbdPZg5kpANR3BIB
Qdku3cA6k82SaRit3drfSDOk/N5v/NyykDJfiPe4ApY1+tHqEK04T/zJQ6ApoSr107kWg+EgEgWu
Qr/ZK4Yzj6woaQlImSdZTu7lt8/cqpp8NQIRcaABmCKHPMOjOW+WTbDXDFobTkSfA4FdCktvSNUl
vdy39xrgnMr6N5zwBottQqJK5h8WiK/KaCBjes3I5irxA6mqrXU+OnauhwgtPbPVRACOTE5xoXsy
EhCjqjTqDKIq5vexhw6FZ4ECLh1wD6hQ6Y/jWR6jewRZmH08jb/a+fpWPbDz/xx95uoRxJKm8dYq
y6ntSMlRkuFSs2xr0uu+xttSMpxVu6tXmHUVo1TUA9lbz+fvic9oxsvXwseAG1xJc6kkzlFSOx87
mAAWQnMBOZ7qt70kOUykeodth/6tXvYcqLvXgoP7X7JUebhXlDeUBZd/zH5MaIzat7YUrpC6Goab
sZ67TNApwwnLYHviFn9/Q7P6mN+R82q5jv8bDTLBDQC3urPE8DBZkwKkZvvjPnWSZSBSsByvC6Zs
kBuNCUQ6wiPsiQYMMhcSEqo436ADZiyarffPsARxgWDHEQypUJWUJSTQDA+gcDWpJKwgoLgAh2vN
SWj+2Cvn9B7u8FSNlgXvJAojKdv/UincukBMSeMT0MprCXtYJVvt508c8KCZGnwd47CaZsduDnU5
4TVOGqt0fc4hjeKB+voWwOegjeKkIAf7ilFiG5PchmWPmvkMoIVAOsYlG4yaOMmbBI+0DeN3BQYN
YPFme14H8pKFqXX0ckcYfs8BDHruOJb5mF8+GKE0Q+xbV5seLwztS73clYKeH0AX+X16vBYq+6GW
br59FdsJQHX8iSyLkGS+dAnmBPpEovb6wdQZQ3faDm0N0rQYvd/s+VafNFpaalKYiL0pBwbyIhjj
PYGcQaeeoJcA9gxe9bl6+pQekHiOycwsl+oL539gp6CJpotRMLDqvamvxg82f5ojRHh6jcGkK9zW
keH21wj9uPW/aJulBYXS9zGK+TvEDYNFOjg15jLgsFo9qNtxFRxtXLxhQixYcDThJRAm54DMX0II
gawU2J19QDtE9DQC7acmNic/3kJ6ODqp5050/Z5kOC2Pfh7AC5LzCccdBaRj70odv6dJ+BVsu+qm
86YYMEIUegqe9apymJ8nuOvxKdRSWJX+4Jjy3iDWyG3KXfZA2Ms5n+Y35oXwJtYIvlhBIUWbNlMg
GyBS0q841LqpLHlT0LzlPbaZH9pqZqax6q0aUWwc2pHUKhdTXB++4oT9kqbRnWIkfMF7DrHimxWb
tJn/n8IeyDC+u7awbxWTQ5NfHlS7dNltcnBFZ0fSOTv5JXtR9vMouGxIcwSr0Y9F0QWPvlyradcU
ZG4nYcZke0IQq7TFKHwLmHSyQDYC4tj/YsdgGB2ylqobesm9HFSsbCB+hW3JQHZg/otlncHxg1p5
1t82MNZquEuaSYJIKXkGGjByfVEvuk+443bRaSA2+FQdwh6o8lK7Rp6+6xzPUfOM44Ri/Th80Jhe
l1hHH21ttL6Vy1bJxmZznouDmP7da+C0Nbijc4vWBN9t+GCeqTRc94ri+A3VlUuwWmHbW3iaQ2+/
s9QWO2802joX8bOKAko8XMG0WxuAsKEFbMpzbayqUc0IlpRrhFvYUASSp9Lc2DaYuV8/KEGmyLjL
F3NZb7HY6UqsA3mGFhmMp5D5K3htaRe5LTwMevywWKTs3Trw42VhgaFUemYzZ4y/r0t2DABwSByn
P/5Wi3GGbP41xD4IQ0FoVoT/RQNc5RsvjQcD2nj1Z5YHiYxzU9bG593e4qciJq3LD6cDhDiT3+OA
4uS3iCzsgj5fPdqt4tyvo12nDdawXHqRqXxKppPYB5X0QwiUoU3EgC0LB4d97JIHOFWSLs8pCA7h
HoSXAwIBEbs/o1KHJaHyn9yQ1JNim5zwRPUbmq2AveplIo27pxNGdD5vhaGrg62xJmaQ8bBqPyJr
oXb31uKWVqIcECArR0h0T3gVTtxrKNd/VbT0pOSfQoOH4HfOivVgnuLtbVRfUFFN5gyrrNMALc34
texCF6XPHjzpgCmzphaQuSKkKnjUIjlcD4DXDOz5sdORnWw+CPGmOTAENtb6v+akL48pzv4/p5RY
TeQ+LEhoQolG6vehVRRhCcmm1tA3lu2UnQg+TumBsePAaHqaRNYMlqxMJkNkJf7JV9AswnM0ZZI+
JqM+rtdm6dU0wqiVUibYgg0YvsB75VBtFYlttl8EjgcvBXrDMwKYVc098d/aqWVUHebjE0KSryZp
GVUa8uEK/JkFYxyJ5vj8UXe5A9pRySL45aHDlYTHSGBvD0+Fl8Fn3jDlLviDPJ/QzkUBK3vbJccQ
3reaa/V5t+Bj1TtNhbMu0zwbYdlNYy/rKJqOPw1E+0E7dsgga7NCj0fBB7OGi5cU+SKb4CaD4tUE
hyPsLQKy35m6NyHp7ASYY4q0PbgWFBcFBJaYxo67tcVuRd8p7dq/KT731e6jaY0upOmnT1gvBUTB
1UU69/tAv6ZA3zqHAhanIuI5NrS4r1C1xaIW6nI1Tc/QbMx6IdGGT33qVTdsZmozMQj//+r2CSsz
YV43ER3IbPeMegbNc1T38OoFg1CgQBVRgJ4ZFnSB9kPyCsuuNEeY4EHF/lOpg+LHZj1hM0MJobMF
WVGpiV/8leANhf+eVpEB58DaUdjtIVDPQYRosGUQb6lCXrh8AecCClzrucBCMmDkRreuMps8xFZy
fvVAExPzodMwpaY4Y3uc2XTGiuEQb1oKXzeVvjpvcxtEcZD1Ml+ZcDIKbsnN2Mybr2+NvHZ4YzEB
RTKF/WkaIhpKGO256uSnwerbR1I/yO7hlScMxQz1LhA07kK8eQ208gnRLqYA0AEFYdAQ334U7dKt
zw0RHE1M0sJ61a40k0N2YHKt4YZraN6h43fCNHJYhZ2xdxL9bAc0mRUzpB36kVhfPR8IRw64C/OQ
dC5PMphbGbVCsGNsFnu5Fpn1tosqH2/47SVWN+aze19rm8XUJ0hvrPTReG30T5uoonrs6aG6+aPD
hVQ24VdrGZSJFcWnOYrP7zBFXWtTXonTcNMFYnF5Pl3sv5d7/X6PLWgB2WPtCTvrh2SuxN5sVqxi
LFS9ET1A/XWomx2pTZ3X/XhIIX4oCFTO1EOi020NzOhA/dHkCWUCoI4FZUURXgDRqfYhHy1YcDdg
Q0xlRWNGqgJVcR1smU/RRGqnpdKqEl6zpy9qbC5MZkkvgpebfLXcjWxQ4LZm+WOHjbeYYCEZGESE
OQ0hizTxkccUJ8va4B+nrHiZsz5V7BPBTHS6SJewChTALTFlOtMxoR8TQBmE0xk5loBa4+F49UAh
4Thvl5sdaSjNSgXNyEyXNaB+OfeJSjvgMilZoczUUJh8yhsH1ModnfWBsd3rOotvZjXzK5GXunN4
HbxsWtLMgUQw2cyLWI6rNGgjwSXjgFyLF783jAycGo+atz0/GTvvUFLN5mz76X+IRjeZ0J35wUYx
uWw024c+tYBhCePBSRywbX6bEW4smVPaahJR+8eMzedCFgsKeVBHW0jkH+rbdH1HpQaZ4R/Sng8E
Nwdr6kgAtTZnwiMnYCy6ZPtYdS5p9gOTCqiUF/HVtZMTYlMjXAOsp7Imc6kQk4Me1J/0d5ZPXPRS
XFmTkPqlz6jgnj57N9Azkxv6LxaEjl3KS1seK2XuSklFr8PtDXIlO+F4PLE5beSzxPXq5clQ1jBF
AnVM55ysk7WeBqvBbOyZd+ibkRhC/ow1eJ/KqcB+NC79UAX0vLyTdaeGIdiy1gA5Gxrm1QSAJcGM
vLH5CS1a1R5rUXHtLf3OjxH28WVLFaK0XyPk4ayPm9Q/5O0cry80cD91nV3MtDuXcPYeIcuNrkdB
y7WNCOQ5ABV2NAWuJW3/cdjY9KJ4impdusmILq1deMio5nL1sRVTnGOoZRrsKVRydpqV5q10Umuw
39UMC+eFEo0MPPsktHKLnOqTCaBUp/zI9a6FcSlKFyTmJ5awzadL3z+T9FuBbTz2aiO2BkE4QRaI
TprTSVmpV8lzHpx/HyWfEjn0g5fx/BpKFygwvS57O9k2kPIcfgh2URDIMvlZN3kKf3gdYY3sb37k
rSyyqRDDmn+8Un0RcmcIBerNn2956Cql+5HvfAwkZBWhLUqCrbbDRTWctxjHVO/zJ+5AVCMR3cO7
LGaJP9umAadx3PaL3XYLft5ATzkV2QRwFMxLO9szHTfsv/ldco2fxnX8BnWJLRBLvJDf4KBVlEFa
ZUJ+ZSvPwXbz9WOeblm5v8YIbd4WGmsRrNNe6f2WItO25MaYrtH+kY2fnhV4aDtuEXxJKBca2UG9
zigd/3s39Hwd+Rc5Q2xzY0zcwiv57qxiEQTFW3P7Q6lB+jPbhm1MSiKA2Hep7tAcGfgQadsUT3uB
X40dNsKFWBCZDG17YwYwPxBFqaoPhReOGRsgIaQI89tZeElTQsHtW2n6A4eW9dHaVFnACiIIHr9R
R7q8xGpXEvV1xu3nQ4V3Ld3z+/XHc6mBqTfQj59xUXyMudiBLTcBJTf/bFmN2da2DnI3J+DWhN+l
cnKY+Cid+xWc0hP0jC8HAXB87kUhs171b7U8zyRM8uhw5h7xBQC2Fed6QUTIpOttsl6IdDfKpgYB
zN3MnZtHaAePcEEa/hoSy18V6AyawE/M8qp6o24FEIB+TzbVJzVGA3g+yaA9fa4IEyQFm2FyzXyv
Flr61p4JdZx9Cu+P3me4bnIoH5mRSih5vgB09+uWtlA0wIny9nRVqQT+RMhONu4cQYV61ZTHp6Dz
naaV7NXMzD0GTSLaFEiL2GQWhwrS5ocs7ClRgzG43RjZF5geVrL86i7rAR8PjK9pCTvbuFdZi4qW
X4Y27bLsKG9QMos8lYARwI1TO5Z44Rg9nUUw/34iiKLF41HAefjyI894gaBXCJLC2kwHubU/yXwm
WmAsgfC7vaHMPS2TgHhZsm4aErwJZqGfiCUs4JL4CUIC4nhJ2pm+8NQe7qE5cJ1/rcaNYO8dxzfo
ERCncenu5NFzmQvHwf+eekJ+UNDiWBDkE0Mp1eP19p5fKGd1LqY053HhpO7amaBO3IE2S8B1xaTD
aZXLzDtoiZjTfAN5kb2mAjyB/xf+BEfV5fBFAlpXTBiSgkauWwVoQUDhKIyPzLmIA24C6Y7YkhTF
SYJ6uB7eDDZeHiNXQoN3UrsaryxOj2cp4oyJXay8VEpKN30Qu/kY9bAwaHy5mKnMiLDZ9IJd3tn/
zUhK2siE+ykOYkcjiDPbFK8mFecLC+aIyLu09F8mutlNAWdDTEWn+gYLa5OCOeOGZeXdBvWW0b/Y
N25kcMsr/AoIVKu59oosYPtnpnrIRv3FQmKWgagJY/VnKe+JNWVZ+rkRyuHkq+qaakS2sTj9hmsG
3BntZXas+HCyq1XWN1oJbWMuF/AwnBZzawKLP3Mi47vtiNyvcGyOSIvajee0KH1pb+KxIhVd9iYS
yaJit+6HiR16tn34sreedSp/f+XPS1CO6JW/FBebG6yQ0ilUzNoQzhiwgdyehhZsNo2WdImeeJVr
aiAjGpvWnwWLX7y8GfcyA72IIQYlMGlgX1bpg7bz/FVwhoQLx7ayn3aIqfI63uynMt8ZsThvHjjY
39aUmS896WccsfXQQBG6tlCtM/HWbE3qUz97XG2jFMtZw+5FSAHVkqgUAj9LQht+iau73CeEUS0F
LLhfnnS/qatR1ws8eeNCQVjJWksJsX/uvXa5zp2X4CrOEe2wmjYitGweH+Zg1+7JuW7q8rsZ42iZ
izOvL9vjjdTXslf4RbD+YMDw2UVwkGBz7fhH8agfdRfgF5jCjHBnrSLtLZ/HygRjiPZDtWl3ut7j
gU7cwfwECN24Dkwb5KZB5zmYDLM5ONIBCzptzOKHwhWygkzNomKnomlDljg5ds/A5p9h1ZfqLxtZ
3VVHveJAMVuQOYBAR4ksyheTXgZGrjMxdsOG4601fuIpP6qeWi6fmz12WvtLmQ30cqsidDqjxMdN
uVTVBDjEoOkCTgbzLyPq1DdOw2o7KOt/MHGAMREFv4TbVUNdCGxqnAys9r8nesUv101aS48CckVN
1gDo9eeeWc8+pRVDSVZ2wKThDgP7K8Wrz+3IIsO0qYPkj/4lXHHOPHr0gjovAQAHb2bcAwzrzHBF
2b0AqarLWEe2tuecieKfgGvWLRPVkf4Qb9wIg0tHeidPvvP0an9C3MinBuWHzVje8/gNPqIApjKT
MwFzTZnHVwTe+R4PDjeSeUiqhzxUOERbqFclSZ/sAGVddS66hP+DEpjGeTF1S5A8VMC2da9GK3Gg
VAfPgQVfYv9fEKfjh5bzGXUhq7vvjc4j3i8/4YP3hX32iWClvrLnH8mH7NAfieqbQWdFxvjbDTej
OMTUTKiL5ak2DZVWyvFfSDCqPvVzwUPPpXuwc1ccl/TAr8dn+zE4sGaHRJmQWjL6rFju3mjMZWo3
rtzXwO5Bp/UMgH3p3pqIDwoM3cQ/LcG+jW8IAKyYHQTBZ28XXdJ/GlQ2TpRZd5j9DYTVWxW4yrWp
0TIArNgEENjvfHLMzU2xgIZXIKjEIvnRTHbBdAfrcSTu872BoNWG1XGSiDYAeIUHWilwmKjc3vGn
+dEZcifXfWPTFwGiKdOYF755KzPw7g2WA/shJz+KrgTp/6d2fz0wQd68cBIF7xE6zFOmvwr4l+EF
gCsSvh7bz/1kaqo2fsHbJfiBJmite5MOv1txpOljilsiwlJCHKSItcHpKoTcs7vBYCZ1coo0Uk+g
W7ZyrtLveCj4VE4rsQ/+ZbuS/qXExzlAFJ//p/L2a+SdCubXx3bbqvUM3Zh7C9eWZkudqvLdrAjh
eV0g0NbLCLK/hdNTXKH/6HXwnJ/YKoGj3esb2BmqDZJ1gksUkSWmSWX9m7/ChImRSGSHpXk6Xc80
tPiuijpDdKFNHyBR+A1WT6f8+YpubnD4+UQz7EvuUvfejh326K1ELOHyEjZ4BUe/3SSBpiGZE6yl
PZhmJnvPe+h/oVb748Uc5zb/lgNY2+x52VW013uKTf3oW+8cWxZu/k7MmmSLtYAW/55q3eI3QNa+
wf8Kgn3onTKzZ9BLOi38pf1Ck8qaMRkhI6S59Wz81MJWhxN2NPPuQxgPgcIa2JI0AVQGoAddg7hA
kVobdxCx7ouGHmhgi0rHfaYeY5qY+wrOEYB33FocBggDzvWeg/jtPv3ZFD9dNNfiEwVjWSy9Mp7C
OgCUdWm5E4e77O1GjuPiiCn0OXrLA6l0TdJnNj58iDE8o6dBP5j92me5tRvqAhnxwwy9L95sJ5ze
6BfYzOjfLFGX5gwXKS7Erex1YJH5vre15dXHL1O3hXVcmSKTEZvVVTGfKXSJV/Jn6q2RwAp5kCU0
ektyZwQVqYE96kfOO68GzX5DE+PWWtVXwjMfl9BbFIilmmaB+965MKkW+XJswImSblwGxSv3u9Ia
GMErOdSLdfZSB3io87WauSkI5eUlPkObCVWl54wphUm2e6XFd6mTBODbZU+gyBU8hU78dHibbzww
XG7DFuKzSvD+X2EJBkpWlOwviRCua3m4M3d4rGFHXuNgxb+1FQdsF/JNBDdtwSqjR+9GUfNOXyLI
vHXLu2ocy3BVV+IKp8qAqJyq4NiraRDPm9vMihV5FAMDQdHkhg+dNfVzJzGbxAeFvG2LfFRPT304
zUH5GczYsNp9JAdbAlGQZnb/m5f1pfKSzc8tQipmcr7VJU5UZ0tBWyKb0vo05cCpi6mi3HaOkLWt
+E+T6Se8t4gP4Vxb+KeeWpMNkTzStZjxEkjuJvbSdRdl9Y0hr4/2OBKtFj56r3bcOF2pU3qc50hV
HrxxRuC3ADFzz9DUBncbv9DgJYmBr4kL9XDF7mEjLEyXc+eWJNU9ywgOgcH+43jAMssb10NSI6Qa
cYusDhUGnqlcx/tTNgDFwy2mcsDWt95ex4dso8Ir131uJs6Vj1HkyKue6TYdKIqHHRyeQB9tlWBB
E31sAKyL+/zWpeqEe1+8KRZI17Di2czElUXGcPYqu9TfINgvNjT2Ofr/gfDbb/IkaC25FiEzRElB
LDnjS761y2hj6tc3ZlkstGqGuflqjSsHA61/kQfq7Asq3SOi8+oGHrxOcOKbnClhFuJixiZFM4UK
j8yp07bX4bY5KzZ5r2on2R54yvFIQdodwalfVNzRquJqSNB9eflEMMD2rJA3rwRotsLb6Zr2DFfP
5yqcKfQqxTdbi2QFHDoFYfSMlDsDz7rRQGkFgZI0+EY+3ZRUDUPubyF8WnvKVvc5SDsfXn6iZ3z/
AN/EW91+3cXF8iOhgexd2OsmCCgaMPGFCc+jCfP56C3SIBWpB5TIO9ZiUm2KQyGixL143ENiq4Dp
Df5oNH9JHLMKGgD6D5GLYf4nAH2cUQ93zZIExVzExvmFjEARaGtHBYnVB9f5KefFU7vnONlM6lG+
KhjE1IYSqxrHSPp9x6gz0M/sgTca2jO/kDexCdSIejq8+IAwkHPKH7Tm4Ir7fWTBP/Tspyj38k50
HnGc9CwdAm4WWnj6mv5lOxYCnyX0zt4mcnA9TMOW+Yr39yrJ/ZvyOkrE0ShSEEA0VBctU/j5Iz4W
VpbBBjTLMgssSBNxKqdEVbRa2TrYqZHiC6D43G/YWLUi3cDelQiH49PhvNSbdQvkR6Po54B8FOxJ
b/BaZ5OscC0CB1x0eC85WQn2aA0IYo90LkMlc6U3lw37Yx7HAjpUoVW7l7rf7B134KOpHYP5cAxn
lU/HUpqPeG34h70BXdO44h17gt2dJpD6yP9lJD4s6NUo3CxKdDs1Y0YE86wXHUTZhIsbhC5i7vb5
U3sJpjDnN4IO8VhQwg3N4F757A8KPOBlp/snA5DBihRIkkPN5xPycffbkuH7EcgHoo2qgWLtM83U
lQxNtH8587UXIuvVs96MaV4P7xmD5NXCrBOcNfqKW6FIvcetxHfPYI/31Y/EMX+0nmCU+BHC3dk+
3NcYznI6Tb+xnEttji5SSFr9hp73EAFop82VUOM3I6xBtZ7gZQs4wHZdr7x8zUVMmi6RXg6gf37o
CiNiEJV6ejXtXKGeJZe7PsJRuD1VRlJqsbgEKo7w6A6Ni8iDF6r+h1FsjZMXnEB7obI4KvFj5nla
zRX8E1M5bdTgb9N7vLC2Hl188zHzN4AkLHIbJnipGL4cj6zYhsoxiF2/YyBRd8yExqnGQa3zDEao
EXrCnc+6kMwWuhcPc85O2LvljOVbFZpKiP7rJJiXrLTJprC294y0Qem8XrCOKgS7nMYqvGd2oxWv
hbLJ60kpwUVfi8jQ0vBMK9pqqauY21I4YfwkF0Ji2VBfy4C87XwtcC4An5uQtNAcb3TTXXDZIFJK
zcfhtsXVe+q1ddUh39naWVjwJbyZtsLkDHtJe0UFBXyION87TVwjsGK5BviKdIj6/KbFtO31dxaW
UbFyYrd5ai0iOBgJEA7pAnJvuTGeWVCvboT1PZZuIIpPXuLholHwDuSuKJkrkGJlfs7Qs2/EW+3S
05txBlfpSkEuFpGSiYEl4bJqMdIBDetf3/BiriVocNUtmwVAz3VSBGrD3DsPZ5AP3SwlqqGczBA9
depAmCKy1JNMibIJGz0BifGjaP1OVE2jDL7YV+H96jqex/CAylYfwFvRG61QO6Q2dSKnzdTtcDIi
a/Qffltj98aN520Mlv0zFYRXvAqQUsho2E6rHpO+SG1KNlTdJ3Nv07uUH9e8SKqQIFThg4yVAt14
vCBJMnbmHfY7MvtQpgrlIGgAQ7U7mr/0++OzEkq3rOq/J/klKdKtUpT0YW/2PPvauKLC5on4aBQD
HQTJCassswKuIu02VJM2rHsLDi4pFXV/ui93QKcdsLV7fTnZ5OuRmQjGeXI0TdmlTsnKN0vFDgwI
mY+m3r7Yc8pOPGfX9znj5TIDDdRLqLtKdhZzLRtWBy/J3YgQfvCmALE87O3EprDFHzeT2OMAkS+G
TT3vBp9Ws0GcWELZGwtruWbzlFMKVtZgCGW6XVLrZIAl0pIw4WdGGGjevwdGMKRrwFvbZrg1UUTz
ONs3lAxuA5VoffRo87JeITg6iYTxQ0S+9tAuWeN9mJAYSsfd5LrSYkY9fZxq94EPjGGjZmjpAp6+
f2XGn98cIEb/wlVdI/paFzgc3pxm/lv3wI4EBNeSxP5+kdZwBYnHE3qSg9407cYSMI5a8p18XODj
/qYHBv25duapbS1YrV4EbFWLs76QL8NCag8BTfF9iYE3Mzsgv0Hs/+SeR4eCjFN+wIpI8RTQnlp+
V90idLEA64KplWCTt9wq+GZ6eEYIpUm/WMr0YTHRscCccbrLluq7lh7NkqXQjAdM4pCJ7BIA72AR
pdhglIKVv0eFrEBH9WXD0Wkm4t7WD8JkbvIT51KCIyomFx6c9bPtwshjXNm3x5EBDWhQOaw9FOG4
SMg0fcCDq5ayp33ANP55po4b+zDSXi0F76KpP0hhJRue2WlD3O2Zmdm4AhtVs3GSdNbdeoHzCMji
toN210O7OOLhCVuY3jE4/FIjyWBcMmKpK89rYzZ1PEkQmZLpr2j+6vF/kM21ICY424Pj8qlacoWu
/MT9R3sGTTUuIV7+ztZRmhxjffEHBiJj+vYbgoyWtceFCzBSOdd7hJpKfVJNde1kMvrXOhUDANcm
+b3vM7sTwNWhtZyUtboaeUzWZIhweyOAqYMQyyY4QGw0WJzDdxFrv9O0RkMjhTWAvMdqcf2Z7djZ
o8tEIhNVIq3eLZbkyZTknas3Z474D+g/JVbjQ9kPJvE2F5K4htEbKFR++eg+pf8NFthurgl/mY73
CPt8vp0NoO94DYjCaX7JZqediZH/jFgim/QGCKWDzmvAcY66r92LtOvM9qqtSZQuQxCP/fM3Aq12
cdx6r5C9/fKQMu3sa/ciUKCF39yOjbFskIc1V206HGbX08+KiMtLrKGyQQ19YICt5u3qzz6LJfmI
wuvq9PC+PgjpOw3W738yE/rOopUewWPlKpo+RIqKIwXwVMA22SEw/zqZUsjG2T1gQU5ta5NlT2WW
xFG6OebyTmS7yw0EsDsNedXicOGdt2JbThu6EvfMuWBcPkR9GjODpxd+tta6dHITb4TXgsxFlVJ2
7dyrwNunm9y4bVYe4vWZS5AE/NK9PAT1TZivbq4hIJCmmj2D8caRj1+fZ2jSKtbRjS5V27G3FJ7l
J7sMFI5hD6osSMRrto3unRNFZCh0pjZPBylr8UEl5+R8RnqjZmCLujzWDp1S4NLnSs77/peZ4hpn
Tkx3KwxlCo2D/OMto652jiCuj2ns4CUw8SgqholvbjIV3SNsQWmkj97aOjd6WE1mAzZ/mNFQqqVF
IvsBjrexIsMbRiHsgSKvEyQff5IxkQaluSN9z9di/nofTLwgJqzpUoUEhTloe4WgeghS2vQl0jJQ
tZ7zGyK73o+IcYZmpGyCzxuq3rb7WILStR0EqxT7szLc6pcuy1qGgOpUBBh12g9f6JP7T6cOVZvZ
46njF84+fmYMLVq40yzeu9F5vhDS5crT0CYOU4mhjQNqnbAbcUvlN9GVypbNXHGUhAVc1ovqcGQf
CIp0LzERYpcZ4ZBP6IsmWZLPFpUi/04eB3/amIUYR1el1Yd3RxOSJ7IAYiyN6azXFYKMa/FF/fMx
bPlW8q8vB/V4uMDtJQ7S2w9puMpPVGB9NKvxkhrH/hEGfnLmTm19cC7YZ2UKfZ/SKhALzBd+bMOA
CKh+XaGnuDrCBtojhN3bnQGkp0lC/6yWeVHsIRAAJjdvy+xb2s1omQAY8dBV9TDnMGZ5eH+T3yyn
k8/es0idMo+rmv7lSsKj6kuPEw81t9fvwf5phBphpeCDhe4ChfxmMEObIO7FboH6qFdFKRuL9wor
qmaz7A2EyBJjCHq4CzmZrFqQsTMKLSOjqusI9mErSHeGIUHABqsxYGf3BSMWkZnLMsTO65Vp/iXr
cwuQY3xbXEnJcAvn8kJiLs0N5wDoB+SHpKfMffABi3Kv6/BtDRJEOKFEuaBdbIlA0ixNafZyZ29m
GNVd8q/5Vj/V50yWD6s+oIb7+Bqo6rqR7Q/vaHyOcRHzDvRhR59HaXR6QeKKxuzXc8p0zIPpQIlB
CFyulzbQxCUhMkcQ6lPCD+Q2nQVmKzMctMvStOkflMtWmvJfGCLzMjnVUqelrelzZT65DN5k+LLX
ASdq8oy5a+0XIrX2ryP+TBC06ldpHxrKiVLfTEVqo0xt/bAvwEC5BxXM7l6TyilB1Q9c6y2cX+t2
PFgD5eQY/9bXgMCL499j/EB0/Y82jmwnrPW4aLk33OYeT+LXOkHSLyo0TAXC8ufpSS5xJdTFFXLs
D9Ege5/0DGDJyTGXBMLe1xvv/EklcLn4pVRsGWqLOUQ7A6SkoK13hY7qDlyg2D39M9dM2yPwYDFL
kMwgZrOl1lLyXXdCZfeQrPCchvLxSDhVZLU/yGDDfD7zfvRBC6y9Fw/La2IvUYUFA8NYfBVJovEk
hJ1p5m532lai/3FkqRqc0dR3H6kWFJvbM07VPLa4sHVUJtozoobwifinVnCoWWSuKK3QYNd/KqmJ
QYEr9SAfWM7+/HnRgRkG0D0d+iJ8EEJrnpA54P5WdzLzy9XFbhgbu+uePK7zuQ242zY6BunPWP9a
K4f1M1ww/ugsMKEnx1RDhU7yZee8QqA2vhOgh9Dt3EnaKH0ovKvDohV8FXV5z+Z6kzKnAuQeo1DY
m8AbJlwRlPgiMbiq+A5dwZgq5ZBzZ3wOanFwAc9yDvE3pykPuPjocb79+4+VlNy3KmJNZM/riz/F
xbh1yzlvpdAVwax6X64AyTx8ewS1UreZMOVGIeTUUSIWq+91X4xeVUAnM+BqJ+N3YHoo8dHqg5zY
8og2VONeDclncZYq+E6uLhW+gBMizgGnpJxWTGHqZuO3N5sote+1ARQg7TKKxGVO8i6GmpbCTLKj
FSe8JiQ5BhTlqiISs+KrkZO8F08/LVnmZy4N5ljsFAs6mOmsmatAHhEqQlzGt35dz1/UKd2ZSBq+
XD615j73FTVxCOaQ5aXbdm1eUBwtFMogN6SesX/4xwmkcOfTE1jHVzat5W9yBe1gNVMwj/Zp1biu
6AIPZFnCpw4dSvzXOGGbOkewTRRLy5MPG8I4Q777/cDTN1c45RUPYDriQmPhXm4kE5n++kLxjxy0
FcUR42o8OxkZpTYdj0Wy+0jthevouergDf0+VcXZw2WES5MzUENY8Tit2TA6BeWgKBcME7ghbdau
H7IPtqWyXY7hpUM49w86dxOpnF7ObBZhYZG8KZB5L3+3fTsV3Dt91zXC0fwvFkHt/oRa0spRpcZx
4IhS5M8DImgAzwo+2DKtfaI8k92PrHKRk7c/099N2zq/q7YStwMRiC4IYIJ0/poNWjVTF5Wh2iJu
ncdIq+MksZSpXq8qQjxhwM4NJWoKxPCFZSxBM92GBqJBCXwDw1xkSKYlucyTXfEgeUX7hBECZmB9
nySvErXxGy817zzgkqXv8k++LuEa79ClFNaS1u9tC3H+0I7SX/MMcWLil3Iz/PCOwsuBfFr4/a4E
U1LwS5+VIGwJV2GYaad5r7XFyUZy36wwOysa6fXlIfTpCkrztD7mFd1UYxr1SE7Y/YZfBcSaIXfV
LMrIpaXP8DMZmzMEuUXbr04vDkwP1mw+/880i4puGVWaiTut4rn35vccjMlgo1XSvGUaXsRGi5Pz
YRYU1IrDulHbqG1V0MxMqFabCSQSzf0xIC6HtzjcOGwWkoxeoRICldrLQgrAZeRgA6vFPICZad6n
K3cAALkCd48pb7v7Hremk4IC87+60EAawU4zB4Y5b4LedQoXEALEK5dbLEdfUqqFkz3XZLmp660S
wCJh1IDUkExwWLr4J/jmpmGRS8EUnUv+VhJw3xBVV5YQU49den/lTsAvzmjQJynhS5hFVCLepFPt
+SMHEREV7KWqXAz/YPYdXz1BNu4rWerT92BspyckdPHkm1SbGO+2BFACuGil1z7M+UqfBt/8gJjz
P24ZKIKEIs3t0LFmBudszIeuTQStJF08KhfTdDBrA0mTwhOgiexlpJSexUXmtdpUHEUjyM0m9D1Q
ZAH1IJ6IKtkXghg+Zf9nt4xteUHyXQ6WjUJ3tc5M4mEi3bzn8iLXeUDhOvhp01jy2i6N09f+tyay
gv2fyt7Y++NH3Ric0HBRQpvoVhVkSt+tJkWSPuFgQ6NteuhPwnG7vksjV177hb2yrCL/b1GoDjJS
EwtArE1n4/+skLpEN75seOJwQ0RkyBF20F+ItZjsBtvi7y+d0uL9GC3HwecYishOOkWvVR8Nw8u0
iMXdG8oRMV4geQ/lVq4/f68EB7v2PV9khej7d94EqisEPcfKehsJUlH15kilwM7L+b4kmYqhDk9C
WFHou2g0OS2SqIngHHByRNWgrg0O/qmtb1+8FnxxoIUPfzkwzogfFfwEPu1CgtHsDEWekCgd74m+
0M0McQTxZjxcMZmNNYQOwtE41Tg2G4pX7wzr3JR098CFzQt2XE/3yq32C+PZvOyJMwRop5ODwsva
8NDmias5CVPLh8IucOi+lDOBK5jelVtkhXc+Kjqb7IOEXyWVhbbr8Dsa2LCWOrhYAE9P5fVz7qsF
ayT17sAPMtV+3hBli4P9MsFDaqyMDxT+RTZw0OFc/vO9yN5UG9PCHp+8Gi04cGedE6fJFiNcfKid
On7l5eg7ZkcMyhDNOq5zbTJnAKj0vFXsy/BH3K0m8feWkc19ZOl8SS21hL5czca+J4X+USeLrbK7
ky4SGfVFqPJLPBaPzQ1WYi4Db9IIF7HdjPWqklZNpZnnTG1O11EzaSI5xO0RTQ8zV3ZxCY7pKmTC
KrNlOeF16Zd1sOKSPgiFbFn+qio7Rg4SS0rqyTOlkoS2r1rb3aOVBz5LnVm+c+C+5raoLTVqcP7w
RxTi+koHG6/ZP03T9z2buJ8T+38r4E6JYSpPY45KKpYzvqYuMUqytLcD1aLL3A5NYX2FpGAStJv4
efAY/AdaYYEH0ax3+FXztm93umyu68gpUUI3psV5BCzBue1rw5xlPp9z2/A+66jIQJCcAiwFuiRY
X/f9mLMCX5Nl7lCrkXYoMUxcRdJtbfMf5FqrQAW5z4UNGQZDKIGvmIrFfrZnkrG8iAPSF9Au5fYS
lN8i7LYduWr81/iDJroiUwH4Z9WEWcROI2vFw12yos1OAUuDkBBzeJXtgBNK/ERxvXGn+agVD73M
PHKf3N0VEXsRrhFr23Q38ZFeCc97T3eYmUNIkYAeBGQQ4TfdLkyp0CCK0CfNx3DYylxpBwqEB0Vn
UcXkaQEI77c/0yX6sfq2uMSEXpVDEXFnVB563CVrptsSxF6+FOo++H8VC4vHsOG6N2I0cAP9wm8S
E8ysXYScq8564LS+cF32h9ZgVFY0XylbUKvpT5R8aLLiJKnuIL64z6RM7YMppribuHnQIuFpb4Gl
7Kh63xOaK2Wjd4fJLJnYeffYWowqqSml+TqGbRrYNG721uXyjhdz41XzUZxoGscgnj6g5mdH8cNC
u7CbL/KZV1VqP7gEhIT7zNa5z+HM6MRlJqfOX1HgGsfQFnih8q+RKUFI0mW3etbOCygpoLKz8AnI
/QJlgvEGXQqcaF7Ll4O59KAerVN2fIs5I2eC9dyMrGp+Vphbv/pa4ML0gx8HPpnrn9/NgwedoAHm
9teS87UYC0Q8HD612WYkwSlCRVRn+Ne183GLtAuXqvwaROhT7Yruz//f5yutWF9UZPUDoSo705+v
YjrgQ64zBoNr26zmZJU9lvn0a83qEhUZi9fN10/GRo0TkvYx1BCeNj/JEikJuGO/liEzdjWBEp2I
YltaDZB1JqGAgkMtubYDBFRAkIAatcBaO+S0A8iYuU3fMNhy7LQ/XLSTDBLbbgbaFHzZHeJWULM6
QPnFtVidYWz9mHjMUdWqVJFG7Njm6zv//xxwtHlVzgfKgPF5FdclziFu4ttDcPPRCwzgGRwCUVQ0
7QAxpuWeptriu8GYw76V1xQvzLLVHLx7hhI4MI4nONAkbEHFvfGyaS0RmCnl8tlAJ6FTs8Wl5h80
SrlgvvuBQM8oB9UkWED7jvBzzLzmmsiB1n+icBJ5vuVwqHN1H0tbe9mGybYn0oeT4gee/M+iLMc3
AMKfAkWB8Z0O8+YZiY9lP+td/4OYVTzXYdJNEPI99beRcaJKIOtXYAHBSQUAwCqY1qFLmqxDNa1u
mibw96Fkl3CexQMgrU5lIwlg5HHu5vKZkuGeXLDTQmhxYKifpepCKxm2rcAEVQKUISPzWz2S9YhW
pzW9OYszFFoP4gfjD7VnZxUw6asMgH/ruIr4SW9KS694nXQPctb73U9/gF4xWl/weSnuT0I66Miq
PFk3CN33QDISKnUSl/m9/6nLKzaZNb3JCC/kurboDTxrgJkiqTApdR3IRrEIgQ7J62EO/sGn4GWy
j8wcq5OtZ6lKZ5ddUsgD1s15nNxGG+yackbx7R0DeJLrW3okrasxTg2nzH0kDgj98FwGM3U5JP4M
bnT9HDQXE7iWeIUozcbPhLr6TcTXOVq7wnun1o737063aCNpwtqNRGUjSq9s3aFT088dNuP8zaKo
5z+EaHeNt0T2ya2RjRt/4IlV7utV4pzmY3XuUmkAHc0515rp2/875DgCOcNpbaVCl2fNqH2YXF/x
y9hdMHA89x2u+ghuv3oJKrPp6yuumjY0eQbSs4wK4WYvAO4k0MOCieKGM5gzdMTv/lF3nhCTFWzf
tb9g4lYBfVFqMTko00uNg4nHobSUpl6jbP72Gm05DX2kWxb1ucrzL5W2/v3JZT8CbnWPyiaooC8t
FlLJqozo3GeYivbWwF7y1zRCDl6f6s8wiVs6xZTB7u8scYrUCaEx4Fm+XPo4A608fEF5NZlPcI64
rE2bhrwl196TuSs01lnku/8y1LsoF8A8UUbSsB6FEg80tYAyqMhk9XkfmXVlqTkewGQhZrA7SRcI
QOMnwjBOBmZl4JDZIX4Ex/+4NUTsQU01WV4EtKQOZVM7PNLquFqCrXI0txD+1lqKWSDBVcYSKw08
dG1AgB4HuzIK8Nd4ik0qgb4c8+r/dXCUQI0CAUvtBsMbz0MSLn/+J7wamVLLBA2VqPzC8c4EVPkA
E82NEEZDSiD8+m2lYuqH2q0viDbtVGuJD3Cf0/L5FEl7W+mDUt36w5i9tQ2SmNAGyiXcbCKZH2Kv
FM7c+j7CnpaqzrYTcyfArCYGh88FU+qqzZL1thGqZ0tQlH3HAtm74Gf7Daoazl5WuNz/Add97KQ9
MrvvziMc+io32m2uzxhQ+2Zom4idtVXQhM53Tq9+C5ntb4pa7Sx0w0+zBXbnWxyOMW2LA8MRDDLi
RXVYvKDnn8fi4BdRzFJjtWxJyr/f8Ox0gVqkapH0CMZ82zlQ/Pjg0P8xu4E7/nMzQRLL6uisayv8
DGo9jPz8CQnbQJEuOIffR6cVBKezn6cmJOIKEfETe+8rRzoeRN9BWMsWXs1EGvilaJf/W7cvSvIi
7a7QzJp0fVweEyZoAMjO5Mi/69YJ2abpoaF9tBlmepjSrAnlgiWcSQGyWPNy5+QY8xnevISnz7yv
GLUDh2qFYI65oCTfk0zx8Js9Pgk345bUCJMi9cfkNm1fzoc8YLjTTaJhYbsmKNBqdF+7TKSS6ZFg
OUjki3NCRzdgrwT/i80GKum4fb86v8HMy1REAiAsDx2Yixj8ZdtOFtM83zlXNwwYmfvxwYFhwGoS
YP9i6k1q9dkpCSb0cU6qzGzqXPpV+2sDjVdGwfIPVZalaz0A1xMzk324c/h+7GwFMKL+ELNEAO4b
KNYIav/q9acZbUz1+sTH+0XNaVi/Ay+YZRKwPdbcz2ZLfzP4B8sw+tXXUqzp9lM9Bjqhz/9jRDsx
mna2jBX3lsPh1ozCsZd3gLW3zZ09u7wcczKVmTO4K3/9hc02XXujii9fVFPf0Ug/gjpR11/ldMBJ
OGgt6/3Ut31vzX7e2KOl+ilkUfeygUPzeSLzCDkrWnvGZNfeoirV+D5t+UvECV4klyLAuWxX6/NV
qsM9mlRkvfJQttEwYTQr//STMu10Cjpd6xNFcXrQAElEEn/94M8s4cJhEIXvBTuSSRaaPv5ZQIZ0
EXtEHPgadUc8WMsG5sSSP6JbcjY3nzasvxS7H8d3/1j2vIDbtZlD85zFEPpDuT6sJVy0fgEKOgKm
idzy/9xxZCIGnR+svKEzFsUIQdFRhRhS+MvjiPzFBrPg8XJOtwwUDOj7KD8QBRFvKVa8Rc6CHWM+
5HrLNRPoyEUarmrmlcv+o9AJ0eLJXKLdAyd0aDUbsKSuEjKdt+3UOdJBOjHTTDgIhcfu5MMD5fA1
YlEazKOVkVnK/I15Q1Y2OBXRosUREJA0uHARBQNEnQTrA5w27hhEYs2GkCv3wYsP1rpkeMR6It7W
I0WShDwNxikolBQMfE/IaRw6+ydw2bpFmZ1VmU94/SjZDauiip7HBG4LbPyxmTHbYrzfS3u5l4Zb
0vmQ9ofxd8YHPrgCNJdFsQAeygoTsEkpr01gwQkY2e+OdFHkOm65xErCZnSarTlNwba8E9+qSGYl
RAoTBcmdJqmdxLnPoSz2T75PMU91+cN7eub2CvUgfa4nGApZXmvJCPtzvLmt04PbzM+uh9wl2eHB
0xhvV6I7FFNB809jMlD61EyTmX3wHyOfi2njTNgloxRkaR2yXhMqoETBCGlP6WqcYdhASSkj1RAR
rR9jjTDkKdbhHzecTEpZdtpGVMsUTDW4TOCBqpODfCedzXQdrjj/SSTkGxuGJadVHJMN7HxfYfTq
+wg9l6B+D+rkBaBBxj4j0C6+UKfkMsC5Ao24NCRLa6ilE5JOzNuOvKfXP2fgaNf5jO6o5IQVK0cg
U+moLCg8ajsm1MB4hiMlvqRlhCyyZU1m9zPsYHs20JhrAEpFn1CaLwRBqyeaPpHjaqVj1O3YGClJ
/JMs5X3WMpeZwZpBX9NKzejQckWuORkemoqWZpp2Yf9z1drxsixlmkU9QAZq3+fRR57NqE5arvqZ
6PMNsQmWWuAuqX8rzcfH3Vg4jTJ67SJQBvMj+IOY2/eoeqSjHbhwRP2JNQPKY/27Eaqo5KsOizZH
Q8eB4eroq+knU1O5qeo8m33jyrxas5hzQqmLcLrschTi2c7R8bMWsnUKtcEFL4Jf58/m/dHReNUJ
CMbHmb6MpOHoSRJeKyPwPIY6e6ayjaPoX0E5PZs6PQHW23KaIDrrrLP/LMjhcBqD1OsLsix71Zev
6cmXayF+EQ5WQQ7xgqktea9tp7XubO9J6zFLi4ADn78El0iSiwXRn/JMHs/79IIvHwwK2HpdW2+u
Jx1YotR+eOpcXhiO2un6SPO0/di1eVmbGYhGdw/GOZh/RCA9brNEeK8dmSdSOIoUPtG57sv15wBG
h15GJ3ZgUx34855eDeIVrGYvbsh4Hcq5utenjldCVdQ5Y8gV/Gkobh2LndVL4rIpZuMbA5N/5+by
bIaNALYl+h3ggMT2ghAR0nwKsQhAXX94aHdpA5ul+fXVe47aVfdnjtxNUqkeIs9ZBn6aMpNGx6Ea
ZrpvVVPbwd/lkQQtaC9lEoIDkQmiJO5EyTQQO20PiEiqbf/YtsWK271acVuA1KyrijoOF9FchXGZ
sg/UUD9+EHdthr88UuLAm1Pt5Kt88SiDdT9Y+t5Ue1u9r5u7bwxvKjTGljTJff3jjyP3zldUME6S
qHk6h+vT3zrA9+XgUIDldII1rJiJ9CVgZPc/5ccwNqKm0q2fhGG9doQaS/PvrcZGXE4roI2g5tHa
deB30ilg8S7SNqjm/GTr2Zwrn4Pf2Bz+ar3SLGEhvF73IFIUyibLwevE9JCWx4a9rSwb0V6waqvO
E8xiCCCPZ4koQvZF1vgJ5OcNUjvCLgpcwxW4mRZmrLbsAn5l6to9gOxPZ5cZcw2g6Ay+DM06+b/H
dJ0DjisLpcgX2MLukhj+3SwblhU1xLce9TphvVrJ/tm352cioF/A8/bZXK1RmXWYJ/Oxj+tpbHIy
kLL9QR9Q/DIZwiP0ttZW2Iqy/IQVbiLzVkO2T/wjpsvhzwkzF4dVSesk9kRa0B2TT5rjb9GnT2nI
Aen1STtC/J/ZbT8SFydIYhL41PwUyEYykBYNHBVitQzelarYkaG3STMZu6+aMgmubiAl6sjy1Q3V
2Q6uKvc4sd1WOUiJR/ugIaeO7/POtpD9UcfYTGTJqSE7u3ZEcbpciNeqrRAAogTNsnF6VWexQZhd
bzr6uM4GAJhs7Bt30paUpt4lG07PKuh/6qN9IzfMbNHOPHK8q8K6UAtTimiWoR8IKEpNibCpCZwA
mYacVIFFypJDQcALCNmKXQOIFi+/9YkkdMUss+t+2p9NqYqDTbQUtEk136VE2vv59JwowY53OnKT
u5mlEL+aXWL5otItYEWZh5dkpP6tbRrhWL6DmmO+ZG6AbUELh5GgF9ZfnyO+b7FC5ABbAE/L4eal
pXsHF68x+RveOVABi8wILGsgcqwV/JHtVGhDvchZezH3w2reli445M2/p58EiiyGY/SIwufF4HRG
UtyijFZXf9X283f+B5VvZk+kRqOlGWu5CA16c5sBwd5JK9Pel3NDqX6dqNu6b33Up55ApRr2Oegk
E5UYUVvQ8VNNmkU5KrGLy7UkKistm1bt27bqdeOL85tQTzHs8c0ds4xUxDZsyeZJX3vMJ3hMszeV
9mcGkdraouDZRM2VAzfNEuh/doZAl87UgIjyqRuVmsmvXGXUAzJ9OXhNMWO70Q9QGNg5jaNGqzky
c+OC3bJcmeykc0rflFA8D3SKTV6CoDEwcIuqGOPONICPkJxMHuxNkKzGWoJXMLgxL9TUzzOF+HLe
uH4zQ9ddP8p/NFX9JmLsYcZeZ89cM6wipiUJkJ0xGUWFN3QbHfeD8YXvnzEQZV63QqWv7wKR9HrK
WZjz04eYxRR9s+dyzqRGPdfWNbqzEWomt8b2t7SjqsV5u0WvecsebcDxO+mK38I48nCsX3bHZ/J/
lMKte+oZy2r6qMlkyZYoylLuXtAgRmih2i38iMuUUWQkptAiTQfTqjU/lQUPzmxDAabjCLMapsMd
pUhSbZ5NlUT/aoDdgUZwlhq12TLpo7pWTfx9OKJx+EiLcSBEmSvGVlsj65iqqIkhV80qhnTfglJU
w50+uWmvhlXehw3/Z90jSbh7nidepY1MDs0m3BpZClEzJlMGHZQKrwgBGOAfBJ4YSfoMBNJUluva
3BxhuXAbZXzk0sLQojIMjKbnelkbFcvXkAQPtzYhnfcCWzaIcEiSAWF/Md3Q+SIpAe4XH4p3Yu/E
0qEJX6LXqh5dbopisAL+TJchblaNmz2hocZQXUVZEMp2itQByfFehs7sFBuG6oGQA9GPvMhUaotU
KyirN7VBdlYkzuVfKDAcBm0VnnMyazPkF2Bbe8mNZFEvKTOp0RhwcCPHSC3MJdeI7dZ6FlmS2qIc
MxTLQ33CKfw96XNva5rxs14Lfzc/TLDNCRX4CF2swb0FFYCWHR/kx+L/Jo3q2XeitzBYMceSQPxz
PMZDfmdqAUWNlmlXm2Y9M+/pjsg05oGk647cD1FBG0Ui5q9jkUHijLntEl7HxuVSlnbLwBqCJvgZ
OjKJmfeS3jUHicQYg2jYOETZur/tEl7PYw+ZcRjm9nypKezHSoeC2g3EGm0H0c6y5zTQTYsQ1QKI
Rcbmz2uUZROxmJk6mjyV/+neBWjor28eAC77gKeGR70zTfrgWuBm9SKLTtplvCEk0Gt7BB3V+rpp
Ps7u3dsOEgXVQB1qtlZstgPJ2D9mdCrQNHZOIYqjEywvRFImGYk/dFKtXV4IPsdrJ/6+yGqyP/Ru
f389GVdA6DGZoDAB9WoBo680KPjELykhVMYfGdc0p9TYxyAr3IcW3I2d2JKX/z/PgOC/cqeLj/07
kzGb1MVPlv7IB2bpGXiqge0VjywHNGEPxKNkSNJxjFZOho01IZjBjrTQVm2EQzKI0YoapgvkBHY5
ZE7tI9bmGoFDgH6/qVinNYofAAPyAgr8aELR1JL4YRL5LG2XSeUl5Y8p4YQSxa4OQLIaDbJCbvx8
Asj99oTd27E13DbZ7ZytgKk++Mh3w5JFuMnCGdkBFj6rwow0/Kw8uItzDyFuRnF6fpt620wRaod8
ur2p+kjDLyqmGUgAwdGF7TM3+QtPOFZ861eP/FiKh7pH+xtFMSg4p9rGB8K+tG803eGPtTE1Lc+J
D44vXXuKWasQh3J9vfLc9QBAlGudG+ksHT1nisdDRQpk2AdnC5q5zSy5wk4yJHsNLqU97i7t03ER
cVUCiW23cv7y5gr10YuSUyssujsxqmiHX5UMJFtehO9H7HqPEgi/A3Tk4xfrdzpui/j/ywcsd8lB
P59ktSMMyzOxKb2Q625ATkKPeOz8vkm3CDYO6iWFZV+wNo32YLZwunCIUBc4/5xtlSZog0nkyku1
KDDYozHXrptBCFK8N7OAQey9jqnQgdKLYeMoTZGzJrQJHC9kyUXqi58aa9aT6sWN+ig3ZxDK9eUG
FCsnGYVtpHLUo7/DZfOkgKmqh7RbNvlKQ8Vh5bALxVORpMgy0M83ArqXiTphgAWLT5FufG8xlX5S
Ar8PvUobUs4WFqNsli8JARMLiTmTjNk4yHICFhGzLLVyIq8c4WWfOQQhrVN46UF/vBhY//BlhZ1i
HcIhnxGvZgbxuKdWaATERd8v61rMK4KonNTEOkMJKzWDrTaidwXW30ujP3jJFgFpmPdPZeLGm34Z
015xgsM1j9AQZ07EoNUtC/CLy9YfIrPY+v34Ylo/XHzk9ZYkVkBr/hfB9IXYbqcP0kNOCTa84j7W
ofv2G7a8BWaNpRtforPane4FZBEpZ/M3y8sAWqQXS2Ei0dMdS8TKx7dXk2cnCiFOnfF6lAmtQtFI
KoRvMNMLTd8b7ANOcqD6/WwGhOr37xCWtgKhuFaY3gu/csMfOSxNoW9TOb2/wkmsuwwiGCST5Ufq
l6T8qkYa4NtyYpKHW7ya+/YOAXSqrTY2uJpcgk6MTLXkAJCPmC8QLSp82UTNp2IRhlHucGxs/i0F
Ql1AQzRXd4PZ0ap/IUYz1AhfLNChDfVJ28uV0SV/g2G8RQQf9Z8wYT+pS8PcH+csQLGosiCBpgQk
g/NGzM+lQmnA/T44/tOuDMcyK+D6kT7Ja2W4uDaEmbiUgIvFd8OR/fSLk+xR95S2Ls0uwpJ613+9
VXueZLZbR1C2OuxBzFhG2OWo+cwnUeNaBO7+ck37UWvuDzHnZbfpW2w4gtA15AePh+pP4ANq+5x6
w9cQq0xPUzInHaZtMnSZPZPgT8UHsN9wqhu5abMZQyMxjQF6I4W0XVwMIPfVa8a2MYimjIUxFB5A
TW/g0HUxGAEyLR+WvBkTagr6vcu8EiBIbeYq09pkka/575sxpdKVLHXCj4dhNrBwWjoeE2vkuGst
0hMlHfbQWi9V9O2qNSc16VUrXl7t5gRsTpSDKEOR8Zc+twVMGTRXP/MYZs6pZqGUL4mA4gMMxaom
xW71hsnVZSeLGGnA4o14kPNB/amuPUF/USV7jcf4isMUeJYJ47K7N22Bhlv5cEhsiV1R4arH3bqP
CJ19NuWiHnstgxleun/B65BkZlz9Ku6CZCcMt0Q4iMBQasjQPW7HiDFOnE2bCmqzlB8hKX8whFsl
Cdk1cbuLcICHiRqVVYdVPmteuqkcLPcTODqgCU2NPAhJVa6BlotAddChXEmiLwuk90gRcDlwRTZq
m5NHXwYrolk77R0+/RZUtRCrsDTw6e4c1TjjoyNJJ8ri/VTB9trvsm8jLHa02NoqnrFI77ka25Rl
t8GQICuAddDzEMWvdmN88qOCyk+U9Z0l9Q4HvEemeV2JNJpozlhLZBjvHke/P7kM38ImwZqkWbiH
kyQ6zEqaKKKXqREDhwk99KxDN/HwiJq60De8eol2GyTCqdwKdVrz5I5nfABffCpOi1Kezn/FCPCG
KZoCjpwnTEP745p3BvBIHH93puUU3Yj7jzo8VYpplc6iA2dRvEQeqSungI+Zc/OtQ3/wUy0Z0siP
Q5eaVYO0DoAzgA096Nwt/ukprg/E++5fm2UYpzxGiksS+/taNmcbrsqcNf6F93FD4rTs4ehLbM52
UMAMcQ8m8Oyalgxf7pSFkFaSZXR+DuxfiBgKgaS2oZmTi4EvuSUxHQ7q5UNaqECs2ggazCHMoIz8
8yHP9QKvb9wHibRJRt4HJe6BAVso2gQ1NUHaRwoLbvevtPPnbffRgQt9RQXwnbrZqJCMohYVea3s
eVyHF+amErAytlGIBJsiAu96kN7e87kHS62bL1B1tDelsJd0ERgMP0AvcVdlHaXcW2j6RJDukWqr
LgWOyIfzdeU6Y1Jq+b7nPhvuZn74ILfu94wB+S8LNlGPWRIcdDKUTXQyjztRfefJYSCChPzOhUPA
XuI/qKCz6w+wF0T9k3IKgk+6fIwQu4Wbh9bj2cUqyRaksNuNJEH1AQitYU4BWQD/VitM94bk8Yxt
EzAhf8ZNcqrcIiMu8ZoUKJkJ0uACRQOJ7Th6WiXqDoj8HmkEWhFZsag8b1fJuHjXGtgQrdhUhmHh
Kat+uW476skzM6FsFq9d/KaP6TIUObvq0y7qvRQilglVqJJvmAO9oRU2Gutl5E2ka4G2gQn24Db2
RtqZUNGp5Zg/qBxbU6qGfHAyhvrG8SFKnGDeoQZA3I9/SwdV83MkiVC5fEW+E8Zdu2xZUlMFCZUQ
k8tMJeypcg89/TtF14x9eAIUdS0bWKU2jKs/KMJqgjS1JelqZ8jZuEOCiKjQF5NzxsQ8SKPouvGC
RnFDL7z5+0YoGKPSzZSUvavSMpw4XA7OIiNhRF/GXgM/Gj2U3W8qifh2BtgcKrHM5M5a2TaCZvgg
NEo/JYmwO9y7oRnep2xrQOSc0IcCY+NQKk7+2a5nrmCivC/sWhaG/1bxCTraYr3kvMBC0XT0KjGl
r/B6zuLRxi/xYmqYvuNW5rCRCRMrJfQG2zLs/0IrJOGdbemc8j5+36PbzI76gRcwcqeY8uDdel1M
wdjlw/OFAJbbSlyTSqI4wpcdij3MQacGSlmTxm6PgBCc/bwa89BKhKBFpAG1r6SZle1PBHx3+xWe
CP13lgro5INd3edK0qcZV8Cw46u9tzYlpGz7cnsHO9mT5sK6JGHPBWv99WFhY46MuwIKDvdhll9m
jymi8xnigWALYDpQQ1SGyekfl9UAmlU1sBSoEKxjZpix03+Muhe2GsgJsztlxohklb4HEgcCryOT
2WUV476KJR3UID1Rz/1rIyuwagsOc1B2JwLF4ClE4BOwXKQpZlB18U7sK5tmXzLZidcS9QJwOdpH
FVEhcBE0RL4azcyEXz317hT68ajJP5rkycfNHhBsAyhhqnX/Z5JC98+900K9puRaNrDER9Ody3dP
7p+E5lsB1nYSWjjLmNaj9khVv+A177TcDd9OiFPyBQe7ECGx/N9eF1BVEw2EpwpxdloQYwIKsQtr
XTk6zXjasRPJlQ7R/otcbcgqDBlH5ORcWaWvweS4b29Dx6MtRrjzI5nESxaDkqKPE0yHgV/tYrJs
JIYqmzR6zwVv6fNZYTeKdQluJQru1L52oXuLWc14972DwJjxeiuwk50hDXkS9QOQg6OaE2g3OcK8
98CyRVJ7fmhOx74RU52WsIPGTWrJz7LuoXEfDFJ4xvXwFoFWXvFaI6hEwvPRqOS7tPGhh/5URhkt
VgrFguueKJpbYe/9syGfYkI+vwoWi1WigTDt4Q3TXNcvLSxS5G4FqvhimSTLRCQVY1HU7fuABgIK
luDVLCXt6F/2Zk4MMa7sZBNIdGUYGSm/+kUTsbIPb/EIJ+zE2ZR5H8XnCeqvg/dmxRsRLKsk81aC
aig5jSWQbDtXSM2x2Rbfm9pp4q8xFQV+s37cxQjP7YMed4q6P8gnIYcrX/n1p6WQ65f16iAVgyOy
+NwlIbhEJ4pub9lvUAkWLk3TY8VH31kUAUnRsdbNsVMQ8SFCvmYAk5aaYLxWK2JPRGT/e32wTnA/
xZcTao+h3/9RlcLFQSCz2zbB1LG3l69FcIo3Yp4tdGz1VumJ10xD6kcdR9GiGueeOkM4MhTOr8sM
mMfmeXEn4nCQJ/wOuoF/m3tBk9agnldZCAEwGluNlsh16Jf74ELcEH7KqNd4QMAsSuDRB62yoLL5
oNItgmSpuw5BynwVPuPnMos6tF11FMYIqgu89wnUeY11GgP9oPXEElYpETyzU+qSC7Rcui+wyvM4
GzKSSkEpESIUWIDKspV8r+f09mIHjOcPmn4p2f2vDscZb+xaV3L2z0h01KGlMLu+keWhfIV4c7qC
CFsDZ9NNvNZj0f9mBG1mLs2cUtoYZr5FTH7Hi1+QUCXYkwznG1sV00WyP/Jkc3rQEYdHVtPEfM6k
ZU55SGEXPhU1eRoTbppTNVIVEt4tiYk1xsUxdkPK3MHHHo1JfD6HSA24mf9dsXCZkPVHRMQbYFFm
pNk6MWWWF0iivY9y97JeOghVcXSx2P7v0Phuuj6rdVHKqT6tGMhEywmRbFEo1ojo2B89jvOCtYbw
t23nfu1DvUoKHu6FF6RgxX7iF7fgXuzDToOpiQ9tWyqLGezQnbs50mLT8bcD7UAr2CcUf9kgZQGx
RC1B/gK9dmxA+PlRZ1quPqeSk2rYA68UkVS/74QHGp58z6var+zmVLug0uCUnUsITOEuGQB+lQ0j
8X8V6vbnYrITyx9tKSnnf640ieYrJrZBgACDF2n4z8jJ5vpkI8LsMYlFgoiSuG+EGfGg5KyOHR9O
dzXAiFlKq+tJLzPQGB/CzAlsAYo5Rp7T+BYuTlXltmgv0+RO1ciOlr4maTmRxTulEOIyT8pbX0+x
UqXS0Uy2v/aN4qMVTRzC5RIJh/xkIMBP/k9CuGyxZL9YZyp07hTQZgc00CKzaKtVwCuuUA7tEvQM
5UxBO0KnvoqAdoSipcx7W/6pEHzCIQWcKKSIpXUZOe6swxV+LNH0GT/MQoCZ0tYfu18X9kPQCvai
ib7JIuyFMWZTuPM1E0xSdU9OGNEPemWYWxcJTIY6JBsslwFRaH5KTxXLbkEhaFrIYgNTkRr+UJDs
KR7Wo+3Z7TtBEnT0lxdioQNwElkJoqkhSEuGrOOv7h+peYX/WaA/v6d2zTJXwvgv++TxozVsDIdF
4d+kio/t/WpFvp4GYFQ8atY9vV6LhJV52DGgTQ3jTX7yspDmJzxX+K3+MMJXNM9XF1FoJHYEFbtw
6TMlGIwnrcWMu9jAtoBzlrL4YcEWUC7n6N6c5eDyU6bmYFGPOo0OtoNX/hzOG8isTe00Z9OFTJkg
R+KQR///LRFYjaaoV9qq/F65LU8SwmFymIVVBOPvG0UxOkorekwoMSBvNHBs69+nw2B4z+AaUR/r
1qgzMsLic+Mt+H1ERKQdh/B4TM5HSXr+3LUx+FRcGkBo37QX6VLE/wD1WpnTuRJF9y+8Av+WBUeT
GZzfLfj+99oy/enTdYyTy7WxVEzGlXyIPoEGzXPP9PG6K6+uLzK1N2SMVG47Z775QGU0HARhG9/p
wAp2Wnq7lfn6XLkB4SiQRAtcNS8F643ISlRAcufAaXdFoqapUWiopIKfcEXKeyL+Xgu5CDUMYU7S
EwDsXWBhlJMRdpNJIPm2ZIU3N0iKMJCaH8tx8sH+uQUgTgyaiP3PJpSJ3JLBs1PHjWyZuRaYskbv
R/pJdpClN4J6mVv9KMesIdsU1TxbyGXDL/90OKoZRP6/T0B1Ni0ILrckoWcKmrI9WLT0GrG9xE+H
kOZz/OMjL8yzfEuWPQxoklZSunsFDGsScB9N1Wf+ZcH/C+hfsOPdWfIprTfbVwlqhwoMDiYumI/H
Pp2uw3CzGSTNXB0syNSoRG4UwAG8AjR2D+TJcNeB0IHb4HPGExhwRFpS/fU7hFLcBDmVBn26rcbl
b+ntHYJeI6F6wnpjYoqhkZsDwSqBm9WlyrvOdetbMTX6eA9v8cFGSTx65BNwKjGf7WTBiNbQ7uvA
xnfbVdenBJLC1xF2PqETrz8PucSq2EDilei3eUglQ0tg+/JtKNv64VjLu1ecnMifi5kXE0qNGw0t
GU1beSFVqlmeZamPkTuzYn/W/JUTqsuDlk9x6LYfzn6ZhpKQLw8aAMDgaDdl6RkGICqU/92WS0B5
tOZaakWz9KWco9wFHkXZbDDb52VswdlB0Xrvus8vFronVSNh/KtnIBI5RjJ9sBhYF6rbdySw+5Lp
fJdkVRRUz6/AJrn66XPEp9YkgQKwMvhRoAecsiPUeeaoURZHz5fVkonh7owiUY8THg6lVBmTbb/X
meDh7d+yOLPbVZdTOGRyOjDrTrojJOQ1f8r0ADWW6w//7nDyofq9RCc37IIZ2ks4w1rx7DG3m12Y
maxItpMRt5NyRt2g5iueOVbrUIuG9zf/vm6zIy5pRi6pUa4/VfrJvsX79YocrVY0je1EeXy+WmEi
SqLzLrhhhFhWU+3ouJXhfHRDX8zUYLQXt2lm5y3H35QyJdu5oMTSR+2WtOvWFLDPW+ptaSoIhSZJ
SGwjrkBkBQA7qGfrWqg/LxsNa5pmxGwWciNZCkehy2H7lVtDPMNgoT8tZDUjjqbNXHkkAoAV8f5X
uSQXg7KIoaHgY25IQMHp4vRkhgR+apa93/d96NsRfv6d0sd5HljcywuIn8umgcHBSP4QII6RCMxq
1eE7/xDm+UJGnRIslulS86O1qRAGXlpJzAyXv/cHMcgx2NA8F/Uc8fIGdFSp0U/0A8E9oXGxMhe8
kM+tp6tVURIisQ6YsGlQmWonbgLORedBiGyTGmQ3Ai9YEHfZzasLmLA4FPapSYR9Q5wOJxijyxYY
dUyUd0SWuL1v1pIXh/28HVZj7gOmmmDNzIluCqNyOhxLxvWydUpgNMeIwj30YWVUu93STczAyZ+P
qzJrgvbgUEcGvRBFeXrZvUDj9ceWTwSI5+sBqsVJ6byiPWxCe+KCG9/qpDH01P6IO2i1rqOwQT0r
3a9EE1fZNBCcl4DH1VipUSfPB3Lh5og5YjtPkMSJhmWWYIwpGA6J9ptbP83NnNOeDvf72dH1X7bA
zIro/K+sRmIN5cgIM7WcPZpiIK2vmbuV7gLhgFo/bvzcNJC8waxlhKsc1NLZTip304PEvLfo1n+x
QpvYN4+7DoGQd4AiEmNEEF9nmoxP36k+6OtpXKRuJzOupq1kSKeLo+XVQ5PAOnm3atHE46BTfOUf
z/CEF41xCys0bBldjLMpmf83/JbjgagjhbzsQ16BPf64I4AlpfkmI4r4U/yCi/KoyLn6PZg5dn3D
FiU7QlTw91z3sSCx9qndHblBOUkGzVcA6byae4A3UbKVyNHfokGy2xjzAzRV+v4Bbp40VUUtzEH3
4FV2057A3RFRPOomoGoIzP0W67zcfX5A1wee26pkwrm9SG8AnCtOMU2/eRrILVGaGhFFvNVhvWEI
MNrh8U9MkUOfKg8v7+R/BorAF+OXefNxj2VKOdT2+r7uVRSygwGOQXLspoKYvKKKslzgJbub8CIP
NWxo38qXg1g1EKZ5ZqBTX8+sj95p72Qktxa0bY41K5zwi3keXDmbOM/hia8Od3UcFMkSnoqw+ENk
pb6J4WTRfTlzkNCR81RDfXcXXns37E17wlXj3IuI9nUEgfJVpzs3JPpD0ozXVTb7m+D2w0ym7AVy
3dkd4AVSb5Ajy22bBEGV+m/jcFy+4pKbb1NBTAWHr2RPKL4hTd6wJZ5PgPhQRUMtG1VZMWp2iLUH
Iun0aPIHAZWgv0KH+W7t2rrTNSnnQqmzYwJM26XBL+hN7v8qdpOcmkRLEtrhSTdPTnqNLvP+23Mw
ZtxtUgCverJKWwsXDA1iw27OO/Xh1MIfk1TXZwgaP2/LPkBXM29nBTrY6nANTZpgRq/ki49ujlow
92llx28cCXFwEizYUoVoMQs3bO3Q/lwxCTbOK7GObGgXQyBPDgWUZ1hng7YlhJXVKlTg6TPpWTAr
lq8194xKAZEQCB95Swxh9Cq4flbh/o4Cv1e2lvrlfB2I8njWh3IP20sSDrIKoTVi5Mu/g7UTNvbJ
V7VZwEbFEzswS4NTvZxfOPLEURE1CTQ/NhiL965yT1yKxacmzUxiA+5fDtQJs2qHxmTY0XSAng9K
Inewx1gQM2r0IrfdUml1rZrVJORwgalluUH5WrctB47uJOKVnSNKHHBUTLS9cO+aAaZbDXiyDyHN
xSJPMLL8snT+qh6hT3EaO5UdH7YmIacUPWewJ8ZPeoKzRmbVjQSKZz0Av+4Y+U6gZ2aouXsenPTA
x56wGVmQLJATqmtSB6z5vRBE1bEZ4qL00OuLKeq06h/UTzy/zwrg4KYam5Zq8YJ2Rfj1uxJ+zZ62
kOMCT3/ZRQ/89yNK13VMofwgH7tAIP07aAUfMINDAlBkq+p2s7wX0C9cxVlXD9GVGHh0bp46/JXy
8Kgac8okb/vKVecky6XjhDQOey8S9w/7nhdH4Y3FOh2/n2X682njBo+Ga2sGPaaFsX1oxquHBkdG
gs+F3573zlc0efFGmGAgwaYXk3syJDP5mc94tCOolxNgzKhO97ckXtsIrdZJRrbndSM/EHRXQW5X
scdSVaPkGFw5WCWU/y9kBv0Slz49DDRPs139tt69THPqmrWZWf3gUTH/VgrcHAsFoeiZd8BRR68O
Qp4VIw58QVuxqq7kcepBZiAJee1LwfuAY/iFBMUSFaBWT7xCoAJEAwMAAeFVzkDcHJRGJVKYdcFk
SPHU9Rj/oIwalWzx0L/9ogU5oT1i3Hcd76cBRQY2Bv/vYbobPm9L7IfnBW/46JJKVpAGkmPaCHGR
kaVMWGWhtBBw7plMDI795qS3lDtbst7glecHea2wGQqnBMc+yLEAQ60w05AXYiAJgY/Yq96eFvTy
f0LFPYUGky0ggMtnVuIGIHyLNttX8UrsWFNyB/cfT7Yt44fM7ir75ybMbSg6pcXzpsecrp2KmgOg
aFNC9+Fzaon0vhr5ZXiyCvFix681VrBdvO3jKP1GT5w8aQIqCFEpZauX6iiFqlFped4Yt4i1LvN1
ThfLIeykAaKH2A/k/e7aWIVEmFJylbOST5CIaQlS+4f/3R1O8F0UcE0ZP6HmI4znAnFu3G9fWZZQ
L890qFYGZ+pHgTBacGn4lau9K4Iq4148y0CJEFn3Fp95BvDjpiny/Au18oYOXQEY6oC/entxeAOu
10VlPlsnZaOsGrV4JtIZeESinfKwajrWTlgY0uov68SwAGvbVD81D6/UE1Uwh0WYaXY0Er/B2yHh
5mCQ6KVD8BgGNyjBHQtjRLhbLU9EnumuaO4M8oWv1G1HLuMAvLLlKbqR+OROuuynrnM10DCusbNw
sRvwfROYGixT6Po2nByg7yFGsj9x+tuMAlX2/YdCgZDs6/ztvnmvqQi9oeawavT1s7cVNmik1Dtd
kZKRKhjzKW78gyd4EQ4P61dd+Fg4RcJ77vDSJuRwP1yI9fTPyAYe8eR7k5m1XOj9Av6vJ83+Os92
bVA9BgYPAyZtxVov0fT+gDmR8xrCib7oZQBW2pahTbUahddRTglPRGuH+Bi9XHQuAy5Gm+6U8JIM
7CWoEiCel/9JC+lddG1YKbFu6LKwVRQfni7j7pPNcQzjaThkBv0Ey2CH+GrdlUmDhUu5AboNxRLA
ZXA1sMfKhO97i9QV/Ynfm50uM7YvHN313No1TUBbkdFE4UWvBZAIVvUoqQiS6FFuMjbBoF3HXbDF
GXnpLUC9vRf4Ph8lGUIUYjxwt2Kz5ESaKM1H2ncXSLnGrG414JT9iN5NnxjZfztCALkz0IiK96B0
crQHul3fv+7kPFhAIuGQYIgz4KVzp75kqnaXCP44v5bA1zgVTgu3rl4jMjiBMzQhZyh/c9z4kUTA
cjJAJe3sX/ktEFr/AzjD/cKL9VxOjW+xHxuxawLQ3iUdaPAqw2cRTNsz6I9r3ijCZ5XOJAm718fQ
dDND8anNl660VDLcGTIHzjX9Kh5xwOav2/09SGOvq2WBZRnLNB7RSjpZi92lbVHwb3iZ1/erNL9r
oJExGWPr2YsS7KcvPJrRtl9UvpanVLerOkZzr0QdblWB2jaKmrIDrpCVP/sKbIWZG/2ASjkWCpCW
/48hQJvOhZsByl3mQsf2kyS0N/8ErTNa/1jCpE43QJeoEWwGZn4/neS848MfnoR0IsyRZ7jNImqd
DbISI5Xes+/Kogn3Ebuk6TzWf6xuCVmtCZWVEi7QOx3PYmPTYwGqe2kIOj2DN9coHVXVcw3rtf0w
XmfHDHPc0oTLqFKGKcTF6My7v3Zcpz2sahv79fDgvOe/zADmfZelRrC5PcoX/mZU09HYXhZchB7V
kEWvrkMkWKtC0tqaFsjpa9IrbEAhspdZ5yTBvwSSPHjLLNKGfNuDG29/ExL8mgDqTGG30RP4C/RA
cTu0hIeuPFll4l58w19uxFvKalZ9fGjpf+0e2hN098yPrywpVMVPGb//vcZVppvIdnlXMDLv2o07
ih9SSzVO3lbXrwE0yL/Hs77Y0IrXQeGAoQpGx+L1pnd7j4WPPquJfAiwFpTMTSqA9LQHwz85duGQ
jgnJvMSwPHvYWDfIaxt5Z702TVsGB8dkDOFsXNG/EA7XOHXH2JpQxdr38iL441E4HXv/hKQG4aO1
a0EfxvH+8ZMiVsySF9BtRpOjmzZ+FQf+OkqSbHqlU9ImJXwp+qZ0hL2iyClnKV0cwABKmhiKj51k
mFWh6UpFtcSnYDH1AB/bV+t0/e7uMlvPCxr1RBGK+NJbXt+CroGBcg5wGlU+QDvu+DJWfd2zwpwV
J85M0x8YyXSWwex7IDPpJfIg7n2IMyROJybsvUMmrKYVHBw0vWG0Ko0cQ972csI7DFg4ZHPq7CYh
z8Zqoce+l55PgiODyYBvNGUTCTS5BtliKtmmXR1v0oJ0Xe5F/Ltid45ZVbQRyLtACHSOYouN9Iof
IHJaCQaUI7NJjwRDk8I87rwaXNrR7A2G5Kk8OUKs1+Wh1RYULZ9cVglIGT9MW3JNKXBw1dJoteSY
ecUQJ8VehR66bwl+uOXDycUfl6DDwBheYNh7dMd1yM3ONt0ZY8R0p5T2/IdC2NAFrMEzCC9PfYjR
NiorUR7SBB7PPcln6kfaorfAJQ5FmaMDIhO4n1l+ByaokvN5AueRPxC8U5K6dvn8r53D/RUS/83R
eNbVS28EbLvpZaxN7M5RH/a69yJlDCMzjawXjCASQwNwyXPwev6URPa6hDlbqEOPIppEXRwZqhSM
hY2DCAb9W/6bhyClgZB6UFSzvsLmWvSUcc0k5idVCfGZHubTHFGYj7eP3Jfp4D1CCUDhlIY635hF
EgaSNiMkX/1mdpn/IIXfZth3mYOYfxe0wI+ZPSeZvj2qIp5Py0cOeD7ysneB8JvzchmiCUqRKf3H
fjjYARAJ5w3ES1CqRw7d10pqX7MUQWcFri7QDA2TPfFFas+gw2Gl5MzvmWLnV3T49kj/ktN3WoFi
fmduKKfDsP9avH1lujM4AuhmEHNVIGRn9gfpeS6woi1Dsn8gHfSYzChaIfWRT5NFz7lf4qSChSb5
3SUOYTQXYGyqtwwHLldsqvrsbxPi1CxOcfVpembBC2KQi7/WtP9jkVCdHLKjFPQdIAIdSNu09vbU
dj7OuEt16/avblU1lWmUhfjHpdmCUeMpvFETHdP0ynYwNcAhIdB4hrTHhVKL+deGqD7SSXw2j4zY
vFB+uop2bOKJS52NPdomFX1yAuA4Xcv6VEOaJaz9OZv6Cj95BYYms+Ylc8MpO0LFr9c9xaGgbeW6
sCA1EnpwOWsKT77w1w7nfErQhS8eAhEeDIVg1N+P8sDvIqkvli/1gxsBzIWQdAVUkNGQEA9Cs7T/
FF4OxfAkHY110dUso+fzX1BLYnA6PZIZ4cOAR4qX0oN5GWlwXZmSVFhLy+6lUXV9ihIALSr6pyEo
lCo2+Lp0Xs7CnwWELd5nO6b42jsuucyJWRkhVLmAD/n7qBwcUsy6K3XTbtRbE2dTBRYakMR62Jrt
Tp7MFAUCWrN0BIW1uG5ijXXbUjjIMTyHUMPV6S2pE0lMhdArPqk/6aNg5ItxVY9mahFMO9XBALSW
8yNSy19EY1IW1JiK2BKoahyv41trjpSX/sCeiIovc8aYs0MYW1IX/+hFX1i63WsB8Px5WZOQuC5k
PCBNph38wJ7podoTige4cSQlLAEMcJPYPO53gx/erjlz2Llxb+Rl78krtPmNYbutM9jx8B3Js0LR
3yAkvS6K4e9uAOKvZWDZEaNMGO5k98Kq3TzEjB/FqnWNyurUChHCB6eym6Lj/VKQ/PmA22U1FOkl
nucI0KacgwPGrUt0ikGzEaairSxJEgPq4jTrQ8o/Tj0Xc4C38+w8L1pRjzb8OsMMvKYBI9cOm46M
wP9C+mBRqa6wlT7g0kxxbLa0Xs523jOBGMBGbV8VABON/2U4xi9+QgzG1TBZVbSaR+hVskH5Bvs2
Rfzq7+DRMamkarJpOI2Z1gpxh+Y1jh2OxjPGYL5tgvrWMtO2NrkOWJi1n0obOjH8x9ygrlQyJy4S
5yq6Grkr/anxDnPCX+3rNS7Re80B2iZB6fCJPx76N1qUGA5x4mQngMu06CfX5Q1FnySvj+vXJ5Ch
f2klFfwVNYou19hQ8BphVhCy6Rf6uAUEOvl1rRBufW9AYrartOkTHmuS06rf555+s6Wf5Vs0TQkF
e4ECa88fAPJTm4QXNeRrs18LuOYXC/Kgxd8HoLFQyUoMq8IYLMlNtOtYn+xuAFxstk0Nme5z+3RS
8NHdVe6P+yUi7oKTu38b0HzHgsBNa+l4kJ3HWUBt+PgkMJVyyCSy4lcHFSA5IP9nq6Zoo7IaiTdY
xDLKKOX96MkgtgEMu0j9GWHmKXrd7qhn9pD69Mm5n4JLPWevkmdVYsQcHIUkA3wOKEyWqjsW6g9Q
Exck0Gr9EvUv3giFs26iOZtlf5u1dVlFzs92hDygfBM8T62ZtopYqHyq5P4+wyf9u/E7UjgKQdV8
2vFVsU+dag0mhDqB7D83q+/MFWkpHVfGrBa1lxtET5G+TIq0OE1SFpKkQxe8LSE7JgG+ZKZiBEls
rHfYMcYVHfQ3b9xg8x/SkhDGCkfFeRHJmteFtCuunMVIBbm9gvFWxVsobrzSJxBygTM0LedV3wzW
9irqfIYp6D17gKMUo/hgbYDbtxWvtvN9AR7NlMotu95kzD0Kcui9kgch/x+/gl9J17FXmZlexpgs
8j94claY1KstLKRfkX2ObNjucG64Xs3xY8pSux2bJTHnS6nUVQJBZR41l/whxHDLMpKG8eSZPMKN
c9J2CbZpYVXbeuSNrFjvOaEjsrcOs2+r37icdn3JEGz9hUSxJ4utDXRuplVLYzH03Mtqd1agRgiG
axxq9dBiAIr17qzvwcArzg2KDnpoE5vStOrsE0Hc1tDi7c2ioEXmTgis1NzWcdcls4zHUK324dSa
hG791VtG+aQDBPG+r37vNoWsIT/VTjdJ9uwcE4I1GU1RAzBe2y6GkuC5C4Us1/WTQVCUuPSJFvHn
PaU/SARNbh4epEnmxqKtwtQRWW8un2MNYunLG1q12el8w317sgzzGqqxzne3VnOz52tTZAzucGsH
iPXHflYdjP6uvgLEZtem9DngWd/MNwQsQPCjnCW+F/6iKrPqQXwIhJxe5WfQpcyayyDcF93xLmyd
ETzvmIdBqFMRUTL832nVVX4Fv3AkWrNamp9+K9UUSGF39aCmYzFkrtsSQqobjmPPgrD1BBzpGd0z
kcDM1BZ/URKnphgW/z54qGlSbJrFLzZ3BzBYutvFZ8SaXBLheFaObBoSa8gRhWIMnMZOCrxHS02R
HI1gKvEyfIBDm03n9YsL7k3kZJwqcBHDNl2EvnMafVMvcwPjoV6n3lPgm1tXlWH9I+WfQMgv+y8T
b6mqVLzLJx2azyn8aDzzErhdTblMmG0Eh8xJDBkCYlfJFqmMP+L4j84KAwx4YQYWtnCqO78ey8YN
0J6ZGL8IBl0IXDAmEXmBxY9p4QdkLMbhnYNJSh4Nne79+kLuC1HyAPoSxuCB0MweZvvrZe/PrSg/
ASZjvN38tRYkz2z+SmnuQyHW+sFKe+qLGcfhVo0jQ99mWOLN2ETfskxocUdmJymCeD74NGOPhIiK
hWW+BA/joefKqP5bPdE3g5/xP5bAEoYDXQi+Hy5zBMgAFiCVFuKJFVRhxpiWKYXFBQ2Z2LOR+vYn
QZSZqLr3S/z5s0Rl3ff41T0FSkH5L6c/speYhH0W8fMUnmYN5bb+qvb2rTko843dPGOVZWZVZQVy
Jwz6fdCQrmTLDMNvrB1aAZ8KyEGQeg1BYF3VB8idYMFj/07LKagRX33LCLcurAe239knGwmxZZMH
lSGGUAnYZlH8QSZHk3UtDFncJmEaqqF5XZUsqbnYO7ixLQRmOo4YPgzXSFSsTYkX6oG5cLBcESKH
K8P2egsVfB8lD2idOQF+m7RruF1BEG26EAzxh146XJI3jrGMio5c//N9pYQDUauCZVVRV4/AF/61
Y76twWXsAyGBMBy6cvyU6wX8cJz5fPslCq60JThnQIbcKzTMMuhJEHPo6judQnNcZQ6AENkSMr53
taWv9goMV8nOJHjleGCcJg4nQctNfNQCaXEgS5EwP3vNQnYTotk1QQCMlYueLbh46NpD5tjQw0it
IGwNLKb7h0EguCfYJKqWsxGMC3jn1ttxx37E72cdQJNLdaXZrXTlp/E1u1+lzZu5Z0uSFYCLWiCJ
oiEL1pnC1mP1koQvjqipgNAhlznySFFk8ieFGlwYeAX0/ysuJYphUL8PPyeKiE64ewed31hsQghX
ifg1wFDqfz7lxrL45kG9q6a0ze9dEfpIkeFbkljrhvTcEW61ToCj9u/j533PHfwBLqn2/C9XCD7j
S5GexX19TVQkGm+1nRrcN0WgVZ06lL3CGxXLEoq35M0cwqzUor1wd12sdSzcS0+kp2phY3RPmq0t
kxL9NhHTv8UCplzZMPhNcbLGmA3ZqmieO4HGvgPPwluWvy++YHpP0UU9wwpyV6tt+6pDhgwY266g
/X2zboxKaPrMAjH4Q46+2MYH8OfrDbjklCcuV8gYMiHd/EqXirKKhaLvWEU+TUO4RVxdvuLIXSu5
F/eDDMPiWleaTmpKYo/sc9Xy3VwlsBxsVuHfs1JcXETnDmer+sIiI11KCqpHocs2FDGTRlsI5ON2
nTdLeRnrjqR/jLbvrmmdMSjLA/5b/uY9zZKn2630QzmdS1GUt2u3jk10MbBCLwwbHrIZI/GfHv4n
mhbOa5vrQ3Uj8vPytwgUrqiYbnNNnewhnC+yvxLGxIwpFVB+eMxHvdMSiEFaLGJQsmvxDhSFCc/C
lB3SzHp72cOuNLh8eEQG8laiNPozdNlnD2Ja/Vj4C55Eclk5Dz5yEsbj0NrKodJS2HfUesitTkh+
UHV3Vuz6nVxSX2BIWcU4khsLhAI3urTAaXFXRtDdUYNB+O1yHSRjzaMotBblHFapmeAMc2qUFP/g
hTcTygDLwQTjORad6nnc6K6ug6AbxrwMZWEUsilVsWg5yJVxtnjeuYdiwLFp+GX3jYlAa+DDMkl9
A7iJY887CmB+fFahUUc2NPebXLrT5X1Nft9530AmYn1+CDp7zZysTHwKreZKScrMO5G9GQUbUuVB
q1BVGLFJLI8aHJz3b8pCzYzM2d5iqrMD62zs2MLPoXkr4jcrUS2cHz+r8nBuBdElCvfSy/3VrQ9A
7YtNRpvqyt3Ga1iE40akEqgvTcYvIzZ/QcTjr5+G1DWFDjAepbu0k64PGYgDbt0N/kSOYeizQGOY
blvhZ+h+1WRpfGEQeGW3Sk6XXtoEmlQFAhNnzfhsFrzYxKOZts0j/V/+S9rSPxw+7lrrHHpQb6F5
mwCM3gYWttm6GUmORDmJjM8KtmxP05T/xncAU8csXeKF2LE1HAscWVVnv8XAsqMA4AQAMNm6bZWq
QSEkFdsPK9mzVVwfdNZA8jsmK2latjnyeuNfXrFARF30YtN03UQt21UwqHunadrabt9kKKJyX2ny
gm2UtxRXn1nNTU7P+s7nD+LUr78m1ZnxlJ/AAw7Yi1fgvMxo3hNEQnCqGlEdffhzT4W30gvi7V2h
tVByPsXjm//nCE6KEQwKPJs+odiQ9wbwYwtbo5wUz1wXJrYIh2ipt/UYJFM9d2Ts/h9tUHEhLJun
WhCE/Z3KS8XWo2DhdhGa1vPSZ82kZfioBCSYmAJ8DnAuhHFgCA8HaUvn/lm+gPhFv9Noh5TCsxEs
orvCdPrXOA0lbsQWKDRlEghrCpeumkL39N5LaFvmFJEjtORDmKFstWDgDLBmrgu7Ci3uToNAGGNU
gFWZEKvbJC6s8f1i1/AlFnV8lLLsNYo1oVTCfY6/FkqYChtvbobfQbeZR31g3fjGP2C3GKFr/6TR
3vumyqu1iQyRLqKO9jN56h/1hzbj4zEK+QlfQ+mkEbG7r2InarEXYpBASgLd3NuTzSpRoQ6XFuBB
jGMe8jIQ+4duqKCF4BCmR1vAeCxqTus9cg5EXB0ld9MvhD9ZrrGZQAe/3chkj00jB4JsiirfZ2e0
Utn7ewm2NURUxSmtLVxzQNq4qBRVHM3iu8It4H6UhMwwwjDylpx/hK4cbXbtAoMiekyvctffgFfJ
ausdnAWVGPK1c6na9WzVVqo6QPYU71Qh67Dj6ORZUqoAPNwAZsU+ayl5isbmzFE9IWXATe/qF3jL
fhsthxIQwcoGH/ma7u8BDTZVt3GJUl2mbY+PQ5a+VYZCiiRcyWlnWHhcUjAYYcbIuim5LoNKzU4M
MiM+O5zE6V0cNCzzg21lS5/itq9OoNXunkFfKOROE1uyDLz8cpLDzINCFGHBIlEbGs5OkSQLwgXs
cT2mb2Z0H2Sc2h6UOEm0PdEjvTlP7SFPDFzxyZcueaSNB5R4nvPXak4+Uwnn2It2fVDjkiIr5gq4
uRI93WqAiNWMNPH18vR1BFlH08sF21aGK4ylwO1SaLa7Vj+3wIuBhTvh2laOxXeDlPiUcU82hZek
xh/idCkHrpOV38QbgbS32N0o2zgNi1sjaFaJTWkmrImG2TAGFoqoCh874ue08Dq14Kcgf8QhbLr/
AEYg0XP5diQHJ37y2SQB0hmCCMG232tsERA/G+2YXOPpVZjHkb6XGLss7IgamDbP9ai/h6oNg75p
05Olf7n1oINCI3rEyej65RuLvgqFXb9ESVpo8KvK+OYfCvZ9fY+0o2/cj5+8QRIQvfvVIIusmeaO
bEeNaeKSGObt66n2x+ybkkP+RTQiBjmqc+HaEjkBobBoZHiVrcyTXG61cUsCCScxSAIVErgWn3Tn
8/ADN8JDJNHumPShof7rlo6VOL7t1NpsmVzViVs7QytaaXbuEJyxx3+G5vUSgK4bNjVP5/QE/vUl
rI7W4cYy3YG9tPDiWeMa7Xhu/nx6mBgKo4r2GClzXFkZF4gKhgWJYQ8jk/zNeITZyKA4oxTSEWZt
4cAi+TJJalXRopWA+0Bdl0ZV0AxluAYl2T4sm/IEydWExzjStnUkVOsJ/3Rtz66Ra0G8omVsJQ+B
djD3jS0hQB0KV4LdxD2uV1d0DWlZu8KrF+6Jmvkob2awfgHnX+A64EVM17yVkHamTiGUaKp01OGM
WKHK/pIZDEw8LxlCW85hkhtSfHVomOH6NJYuIwWo3sSkgiSkP25zJZCs2rjXwgjIIoSD1OKRZlne
EC1HUfX19OXIiZBPYrfWyoCaaH/N29Yodu7ASMTc3iFSCpwpTUtSGYxvrExOmD3tI5v77yeGIxah
VLABGPLx6ugL6Y+VCImQSWuAb9zzjUdR/oPbnCquSYma8+tC1KY4UFB2lVhdN6iLHCM0aFPYJO6x
/pLHsAgI3sH8IK294ODRUunKcND9ZxApcaoqNZasNYLcJtGI7WI06QJt8+KCc+fiUtV4m8+0qBG6
WQ1MAEG7kaCRd0S+g/D8mPIIDqRDiNBeEwhYt7ShizLdlZ6v2Q+dewyMQ94K6E0gz5ZLuUi/MYuX
sZy7woDVcrA4w/tpp1nZf5AvQqgdeFMZAeIGG82gtpxa8ntfuxRNA2moKheBX593senEjFFnGgOC
0LUxUM+4cZQS5ICNy1lh3qWH4T4+axilratbLOKWGwDyD90k2UCUnVW7DruTImz72/c2lDVxsxnB
phjEd1W3/F/3VAtfuFhlQ0XNSujXh/Vwa7odRcLWa1jybe+rbD/CqpGUf6zbieyfGxWdZCMnowZg
+f33nA1I0an+V11FM41HxT9q3up8oj9EIpNaX4Uvsul2aqXTJWkHleRoqCLAZ6R9aNJXsBUbd2Ea
HItWG3f/L1hZUIIGUibA4bk2UtaxlLr9P9NlQT+jpzlXveRmvhZ79aZz9KRTvVA6iWJf2tsgy5UT
JWnIZVDGTFP7NGPWyNgBPE8m8DTT/g8UKTd7FgUrfcpZcJ+ZMif3ARcQPU7k7MPy0vab2f6r8QHW
16xP+CCZk7Nb5co0vDI6SdkRHYdAU+alpPvseRIef+TpRbF1/W8zWaL2G3DM7OO67d+QhwJsIMnS
PTdZ+AAY03ce03O3LVZJ7Wf5ysDwZB2uNhmAC1PPGyR1n1FEVMZ4ZK/mJT+/mRMwWD80L3rg6k+O
Qj+ZwggUib0fOr5x0KJrfHVPiqcpwRUVkPoBrBSN2bV6IzmE3pS/K1ofVV3lvOgPOdMUYrvwrprM
xJcfOA/03j8TiQMV8UficjMw9XMLGELYhWqt4nCsIGydHOvlmNb/61QWNRD7Rk+VKiZ78cQXAhWu
YhrOwLx47jVVm+2VQUjebuoznQgpbju4LDbCmf2mC3Z+pX/Ye7nM/u/C4Wl/HsckchuQO90229xp
RLR8HSt8vRKPQd8BY47VFJahhknngkyAzh/6h12VV5isKvKBTYY9iRgAGmLUm5u/LqT42RjKpusN
CHB2bKakVg6Sphj6XWOj1/4gowM2//pxPFoBG3wRXAtb3aqsgJ0dlxonPKy4RlD7kfyPPz6lCA+i
SYGWVw6AtSxJfHAUqPbMI76PXhF6EuttWhbEUdJg7g0fzb0cL3iNbx6CRZYVy7dt/QiMj6RKdnjy
pC43rtqd86qLUVXGVnKogBd5zMwpSDb+XDTZwOXRkEaSFSKd53rMmC/cbwIOE2U5YQ2NreJUqdXt
fVBhGRNvu55u2Ya8zGBDw1ekM0YkNsuUSF370tAXxun1NL0Xd24BheB4r8y3gRZCl80kk9vS1nmj
24ZdlM0YNFc85vuwpdDHDSBAhv0dfeDH+MpC/3V6SAqrOjOmvLF6RuFpeF/8deAKOpjz9b8x/wzu
KH9JyxIln367H+xYmH2iMjhuqorTwBsBTZtT5ghgbDc4MN/Tz8uO5OThADQqGZejopws+cxnM3yj
A35pIOtYDAPAklUf+c02OffUfavNDGR1mHOaaH8EIQ6e+Ca6ACetseGC8HKp8ZcdzuEL3cqQoFdZ
4W0qsGVQHdwoDBLios+077o4VN6M+W6GsC4oK91o8weyv/EEV7r571Ep+xLuvNSYTReEQ6qIsd1u
LJ0nvAXK27AIAWwRWpdgC9k6zSffYd1zk+nl0xrMUfn9E7d3Qy0Vt5Hjrkw3eZ3/MWv33q7Fp6/e
AFdzpIWfcXSoKo5UsTyDNsHMMyVWHqrZYc0miOZjvrruE/TQtYilp/YerK9qaYgEaeVBMJ+mbczi
pbH9yPXqwrzv33I78PXxmaabhOY5iR2RgxlyK0tM0/FUqoqZi9sGyqJeqTUKDfPCnEHCPKxts3v3
KYXGF5FVKQdZMmsobuwQ9USyZ/JNqE8mxbt4m/8IAedqiC7jHuY8LOhdW/Ayz7JF7FtaG5Qe5fKF
4MV6ZuGWKaPq5JUtUe3b68kMxasQZ6ydXb/fpYgqnURStvjEy6tXZzAmQd9wWWtYuqBz3sMi22J9
8+uwMZacLbspSLX7H1W5dlZAnhrWtOYucB+0lH9l7zzCe0zfXC7HbxInVU04mdAFuqeypdWI0Pp/
Fk20z9ZhcuMrwJOP1DtcoWgDY83ZIxy766pthVlgxRN4uwkMAU/liDJxr1TrQCR/pimLcwW7jj14
YGwtsqzG2qDx0rdaGB2RuMg3hc/BHJpnTRZRaQTl/wFflkcXlEp2dpXRwxx6Zdym6s1lZiV19P40
KOSvs2bBGZX2QB+gjsQb1bJxMWFiMtQlJ+29B3MX39WCNvqTlGDdnVvRhxCkiDoqmkp8JtWUejMC
OXVCOUGSdup6r3Rt3qsSHG5gyEd0NPxax3tKCG7j8F+wYho3LlCoc7USsE7ZsckrG4vUHJukpm51
8Qna+Frc0SCWaPRmdFjMCLafD3AsB1/ontpfeF+PSdv5hi6SDR/98DF0reLQ+6944NobLu/beK4Q
R0WQ9iocYpn/hroKwyi+NfH34mrGI7BBXo4cx40DVfeO8rK0e0ZiKDIlJA031CDpA4bBguARvYXf
gVLSkY/UAa6JNh9Ecis++wwlHy93nBBtmjVW39RvbMjTLlT0E9gTyseLWGZFgT9CLEQxmu8GUtb0
Re3M86OmJLsnlqSS+NxfjdoBn8qz5ftEXqXbGP2JJdeufFIWho3DlWci1fovpFFU2BZrVC9llE+i
2wI6chRkdmsM6q64rF+y43Qx+UTwjFPOQsMuxx/LBnbbFI49gXTbK063ldMp6Ls9e5BIyG8yIvVe
SKsLLZxKLHy9QyntcEY4CdWldmlJTIdLEONEU1n70ImJfIu4/LXXT17bwc3c+/BcnyDanDRT4p1w
51nm8IuxE7pAv9iVvkiukSFzHHr4gj0XJAJhI16ndiQC2pgvlouCZpLffcgxQfHSN11+FS61SotL
E5gV1zjhAwXB0tCCSdPls2adOKz2WtgTHdAcIoVzi/30QB0bXo2zoMoQZ/Shc6F2jigX1o5GvBKB
rnWc4iPqngNLpJlhFsNZyHyg086OL93+Mc615yLRNC/ch3GEmy+Uh9NmB8+6WOv1tB59pE4q50+J
9eLNPuPRsOXxNT6K68oSKZA4H0bt3nPYlY45ZR+BZ7HKtC6Wrn4lDPdm0AkDn0xcY55MDLiXZuuO
qCzAaKXqwhIQViq6+SicKrUZzwsXO1RKnQT6MQEIXtc1pKgcqQEM+IW5Moq0uPp0fKBf2eZup7bn
R0cPpxZc1PSsEm90ZXu9cDrE9lMS1JOnXGCfXyExDJ9J9btnPqDjeB3MYtJAhdeewRp8b3tw1khh
R7y/+38DMbl0X9oGlv0lZmZh+XnATwyrG/5rCeAz1lkrDJtga+n2TwnZ4ng+KO26+oNKc+fZDRG7
hQ0TKbdRr4bi4jNoAJpC9kTX+vH5TVZABCN6tEJJdodt0nlo/B2vwmJyq5x7OvWItJQxnBMabhGP
DuniePNFr5WBmBw0NdnrSPAL1I5B8y+oU8p3BoaY7TLtzkBmQmayES/NAfMetgrAc3LyBw98iBJK
MVWD2zHXSmPMZKhx5hIUz+IBwrTsmWZ/q3yIOWmfSxfeu27LKI/bpwFQylKbd3A0mLeC9wlUAFQd
tiS8ANkaymLGl64efvnFaxok4cSGsIbL/d77ixwl1rc4DPYozNdSNwtXUMsuKgmuhdUbPcEuebLo
rwx9uoWn4Jdw8a0uVIkdoakMAzbfhNdruqstMG3G/j+wIpUEpE0wth5rvZMN3an05MK8HwkUtlwM
6TSnIo6RN8eS6stlAEmm17LQJU1UKFJctKcdYU5Vqeajv7Gw+IhjFNeyt/5D24udfYtT2UKWPCKT
eFN20/4W4fijq6kYlx1JqPi+mX12h9opvJtQWRJZ8pZ2eGa4M9XXPxrJN4p7KSRryGdgVsH3UEsf
7/6QI9K20A2kmyN8OKDtHNG5vk6lUW54bSZkuvTNhqEb8pjI1UxduY9v0EM6bKdPriOLGTx3eW7j
27mlhLZutOxNQ5IzZp8kImJsMNLlOxUBlHlddCiznfAwqrMeQ6OhA3XrZO2d01y8G/eT7kUjd1CS
3LgPdz7LdFVesjRxNehHmXbXg6S1BeKuqlQFuTqVWeNywzngD9+wxu+dbDT/CU1SHB2dZ8Vz3HMw
6H/aWsjEpzDZW46NI1A5Bo//8MzhMxHA0GWvMkYTWq4Bm9TFYr6xZl6BKCVRYvuaeuMWrXSUTYwq
JPmpZpwQDsFWhClquAuewUWZ+RF8ra4eyfZugLkqHAUhCcfs7qTRGnJa9e6zF33B1fmBHdWZInQD
huVsmA2KequXKKFNEA+XQo1Lqpe7R7VpeOzRDe2WbDm+Kt8achafVxI1Er1JFQItRbJRJCQf6AYJ
xQsdXWPW/zYGK9gd5/jns5MWiBOd1E5oB/RnGfEaqJOXacxYu+X8gv5QGHVU0A9HE/Ccu6SVWokE
rbBGmK8MetdaoIjffwVY5lMArqeyvLwUS+JkV0mbxJ4O9wQXBxRPuhpjdm+ofKFwOK+RRyxzXifr
wVhgOW+AQCfQ+N0nI0BZ884YqFl6XMKNdWF3C6wfxUS4BbZ/Xrrhqs+8jLDiqbGpb3ukv0ex/pNL
dNQkRUwV/zuQ2e1ZbeeVPGZWiuOaVGFayqjc4YRRlHdC8QRv8pSA65iOYvjHgf0Bebih5uQJM9rY
FqW1i0Za4XJifXBj/QfE8GQVaRADArAllO19zk4vKP3vm1GY4iDFGjX0vAv0FYLGAVPSMS9MpFn9
vx9ejaBc1hRU6PqLjk3okxs+aY+++zGKZUnb/cKPqcI2Ex7Q8OpaG4ZeevDA3t6DqvlOp1h58ZJm
u91OBHL0FLwQWUn3dVCtpzOCu2QMP8nx1p/QPRM0LUdNpHI9de1Drr/9iY+FFbrc3TGVcH6Iajhw
ShShWJ9K+VjDnRI4WLRdvlYTi/HVikqlc99qJAaa3mzaBHf+QnuF0g8Vf+kR6Anmy9ZYRIQGJkQA
f4bB/C06O0IihFJCSC3ZaCyjxe4j737v6ISbMd2Gm3+sGr7eC4B0m1zoJKlC6AixrzCYZjt6mGMj
WP7UCxU6w/594rqKrsf0+KldbBm/FtX4uYP1NvDpgRO1QidzEfhcGp3Kbh+CckvWh8yay81H1XI4
o3EUNv1qDpqaEI5PzOTP9SYnVWtwUY1RTJCPOnsX+GP0aiRl8jDpRJQXyAZKsw5IM7XP8x+74fBj
xOTDveziv50geUrnGLqkP8p5bwJCJ8KVbtdsbIT026B2GiGWzf8fd+Hdiunm6e/lGINFkbr/7iHu
vkoLrOVXQweqVJO6WxPixVg0NZ2stTyiKaulM46hI9yePUTkSfUpZyC0HApbc++FnjYsFMmUU45W
U9rhaSqd7CXm6xlKr8nx0WCI1pQ2EdaLhz4TSdwtdsl2+CPGyF4hPuVa/4tL4vmGzFo912Jwi4NS
+fb10Ed2VRNsagwPY9k6yCcettstchsQYX0mcDF56efVQYvQCq5w7ZeAjpS8WfxI0Cq7Qy6lp9FP
G155Z1qfc5npE5uu4fbFIjuZRQ8YN/t7dbbK1nX9geNclX7/BCtu7iNLp7PeE1qiwHdsJpRUq2fY
jxqF5Ga5hJddA5JTOfHABfXWH7zmmWUO5HLu/q7lAoaIlpy95rWoRll9nxx2TpPA814nAhywdcq0
Y1sTAlz6rc2/WKpN2t68AB/JQWftogbvQuYG7gDmP95odzZJzvLUYIotaKXTeOcSp2QCnre+YDsC
4wC/Hw3OqLaRxri05rzYOLMOn8uCXlOQKgCcbqcF7T9m4svHHQ1VkXthL3jf4sZ/O769Xhphh1BP
dNPMvyeuloFEqh9i7mm5kVRaAdKlDrN2w4nSVNPRRtSxNAN7xNzrsDJidcMQ2Jd0mplrJiwGIsyT
QmsTdaXyy87ojA1yaDzrozm+mz/LvwGrZYEPMKkyKP1JdT/WmgS40SFw+NfA39wygDk3flJYdwYw
u59eGMs6VzsK41kl7wUNNtgDdfJCqF5FsR6SVzxXUemMnUPToErvHumRimC5v6flwUxtuPO4YkAv
RTsFM0DScmHm208apLVAF29M3xVHqN+jNSWuXFSJKeQSa92G0wXFcjSlWNRolH5i3GSLeQRlgnNJ
000zqmkogBEFAzeKAJyDwNpwitkUz5m4cSXMRftGOvXRZmuG/0wiJ094rMi2vDff6EuG4on+Lnhk
ern44BeQFCo+J7Ap0c7tiKwm4uuyqPpIqN2hf8VKRNpCpYS6mT6x7r38tHrHQ+1utU5ofRgHgIx/
2kTbjJxCQvJCmbwqQeQjiqDx3n4dx7syh76KnKXWMJUpKxNO9PraKcB1fONvi74oQ3zU7vYzcvnQ
qLjdWQ7fG1t6W9ELQb4SREvaCA/iBuAC3hKdbg4YWU8vvPeFwjk5MZEuRYXaZxb8l2vaRi5Dl0Ns
QR7DUPsj5Q+yCxVrksfM2PLL6/ng8ps94jJNTKmozFUdAA0L4bLa6B2KnXjKlb1gNMuKUUsLT3ng
hfbBgu5m6lL3My58nnWXPvGKlgEbV8X1TYO/IgSHxlMKRg6nnwOVD1hqmr4UzRDED7ipKencK6iR
6GkTW0sXm24W4U1Col+dW9TB+Z3sRIbZXWXvgEdpRiW3MqMs8366e43LQ9Jo5Q+mzuxn04vN7Oj9
HZocgzC/oZqpT+0CERv2tT280GMCF+a09GBklN4WHoPbKZVh05oT23/GQZlFJs8ioYFZsV8576SB
AQ3JNYGw7kzLsCVbPkr0dXB0qTmSxlIuINMCmJGHPgvGBRqutMO061sq2nH5BJE5r47rCJc0WgBn
JDPFMKjYhbNAlsLfod6/UiTf/KxDbmeEPmAg6XZE0d3DAheOUmLgAAOq4RrM+aO85IjZkcrBVQDb
KhN/8D7yAL54qGZEc/Q1T56YsdhRhS7ABw4hyfCR/yuzrlmXSBn+r5105b3dPBhCK9BCqxVoAPnR
Oql0BvTmCDOtjumbRjq2IWv6/98nVxHFzMFUe0idOxCZHz3tGXXtOoQ0Rz7ihaqVtv3aX05LBX+Z
gKNzEbmKKeKD4DyusNfQ90jIoP0vZdwHzZLwUCSkjCA8ZZBrnE7iloDOH5Edu//3rF8/dd8zJVVV
ScfCh46ZbQSz+ignTkvnPGCcFnRuGQSSLfKsgLWsBepdRVgnfCpFNz0lW/GZpOSNTcreV3IApuIp
oA+ZosCsn/eXOUktdjo+5+dcSCgakz5q2RBeQ0y8v2UT8vLqXi8gIEHjeedWGQmQvi9FwqO0Ns0I
9izm/V2BYVBNR2PRR1VS3i/JJ4I4e+hBOl0HUtH8B7MVDaHqkIJxuknT5XQ990jjR0Ri9rTOTs8N
CTV1Lhd5l3QiO/GG9/bin201GNqzo5QCpriNbS4tiwAgk1VrwTPTiMquq73ZhHOEX0foj2qnX6T6
hpK+Es4kYr0glIzlBWlcKin+nvTjDnmurYBeke4tYt2oFPCyrWcsbwkv5TUAnwNOIXgVEK++WeFw
m8ysGrVgLOptyHGgLhnHxtPYwrUnAMWXSa4e4TDE5fiz948wooFsyfnLavuyMlW7LN3jcKHkFyOU
Othtmd5IBjx0Qw4VA2neduZs30lfw+WjnkVTIxJ6MybZW+3OD7nN3F6/GtODsTzz5VonFcxIX3ik
oKqXwyovGi8JteUuWMhODUUi69nCUzyHN2Af7DuN2IXociwrkFySEVMIWaByctMFQTC//uaSjBBI
TfipmA0Tsgz8m1PbAS5WN82J/1XyN5qVizh4pLmNnMMcvgu2PYya5wfUhVRJmJS0KRdbfo4ULqI6
wY40mTtusP3Op4r6f/t6gdYq9ub8GZjA7v/B10cVAb3/oHxijOVEWC3uv8FOCiWt3sz9xU37B1Qu
BEoZdOD+wVaJnckR+Cit1mlNzL17AZKQs6Sm2dd8sxZ3fAVsVr+WczGMDGc20gU6q6LaM07vxqXE
fGt1UpCJSulBB2mWLxePks8bgHqaa+cwLSTQnSMYpnMVeJyFNxGHCbLEAM3b3R/BlAEHEdHC7Bpo
Z59DAIys16D7fcj8qjyt5ILK5pdT9vAuNkcPickURKRMo0nT1EnmrLnNRbb94xdvKjBNVPYuYRxN
+bWG4gIiZktQIbjg/ebSH98jdpeGy74x6AY8oI46ggdL+43JgGYdyx3QHF3J6Gxm1t3dikZccLxb
UzJYS8UXF8XjOATKFC7EgtVQXO+sZ3ftzXc2ixWPVl7mISHxiMvb8wCw1TUgkGLaxMAVL9wfarBJ
dYirEM96qOF3ynfsRDir+xxgDbhewL6k2+XyPMmvuc9gUoMbEWgHBOdf3KgNvsLCo4G81XnN47XY
19Y/FnzMZysFKIXuDOBUAbG9tH1W0Ro/oK84/T4nXp07BZo9oJChc5XLEGm8MpuCUIJ2c3W5117H
z1K5fawZqGR1lpIk8kMRouSyHAz8Eq4rXZ+dcScdCPir8erfp0AoywVK12/McOOb+9YuvAvUMdep
02VZ5dTLF7v1WwbBuphY5+vNJGuvn7T0YC5Ms/3zU8v+REwoClS34SXI3I1r79ZTmquy/N2lvsWP
7EJj6QFlxw/yGgEQ8jSMMZnbdnrHvOImMd2AFFS+MdnvdQbBvOn6Jm9Voq2CN6Cxb12LcxeAt18k
J+36/Uolr6Dg9LmsIGxhaI2L6ZhyFZsJSmnq0CRDgQigzxccd5BurN/v5w3Qv2UY/I0KQ/gQN+lG
f7ibatruCNDlVUomHtZ6pPYCNPn1uny8DL/VNTIlWwJ1nOHUT3yYYOqKF9by4g2ukxaFV0PDgtEG
I+i/bPnZCOuA405ZFCVT7mLi/UHVbyprFuV7hVgN3H3SQelYaNDB7rpT/Sp3H7IUqTwfTJ6nZQaC
25FVF82GEkZDVRV6OtT9e1Nq7FY9mRB2FySDAt5WFxjJPfDnGRdIOh3qepuWZH/j8P4vlBnyH8u5
twG4jAzLofke5FASuYmFJ3O1ma+5VLqhCWB5ZDZb5cODso7Y+sML4OeTmTlgeWMx4ok0B1sLBacD
4Qy5PZc8nOvwujEBs9MkUZPRCFyVzYb4iTJ5mBsiUz4UmgOCVceJutP4bAEE+pgsGmDqBiZd62EE
s7VG9jr0F+FHanLXjIyEh9gupZA1wzjnrzu0sXkk4ab3MddGSNpXNci1BYgbYWf0gz4pOJWkjrsi
TtBnIsNprfcdV0vY3h80BU+QcS+qwvuSDMLL1NxvSNNNvQ5/I0/YD9vyB6Vvi+4SA19SxhVpWkz4
bWTQ7AoSSS+CrRijW7Kr9mGusA0yCQAq81NW2v8xntNzTrLgRsuuTkPAll7rrZ0i+IicHXVthnZi
oKH3hBgSON1wb/FdNJvXUxkmgukZhfH0GaBXallbRNfQWDWx+RhvLS6xO6WarWbGvCeBSD1/59jQ
JeDyYG19iSNc7cbCT2GEREX4AJRc4VtPD+ba9fJeqNhdMH2TzKGFuDdqa6epT6LWxkbS3vu9JC+z
S09jftOTZcr5VJJ/jPzdrF/gSqk5AF89sL9uK9E0BdlMeIXC1gWIZ97mK8FjNB05fWZP5w4qeGDP
OAKXSItvFQZDWd8X+7uqnrZNCwsZIvXVy97egvdIaRBzhEc7J+PsQneDn3rej+UX9BF6tHKuvr5M
g4QBy7JENAvguqOdCLpPo1ng9OdBcLYpw244tSxOQYFDcvl8qa6RTETWPBR7amt6Imu7WIF3iO+d
nlg6EnzmcGt8vsfAmAZhYGZoHvEYbqrdSpq1kVQ92FvsRmbcjNzTbVtlwuBL+6QrpYYvxeYmqZXs
jXh/XkrUbAatid49fAStEPn5FeDlQy+XchPKyG9I1Svs3OrVpqQD+UYF7v7DYuRrC15vtZJ9bhF/
0c7GAkbD5A5Cwas8/S7e2WpDPcffKu2ntZheFs7kLKLPNsn5u33RDnDqHzJ5xRGB0qjOVDu04D37
ZDGLQztzxx4Z11wJKz5u15co4uFrVnGxCSP60mqv2LlhV0jEXoeVOJAbpRRZxxsSf/yg+zfpLXM7
/NWsohMvAcnlucyupc845jUHZQfhh63nCV5nlkwXQOVciaj6UoLzzbogEvpUamYnk5c53ivlJCtG
npUduXBvex9pqKC2kwovRjV/mUusaPsxZjVquj32tfgsQhLTQKbWKFoOdvo/y4Wvy2dSP2uQ1lCY
ZJV0SrEOdqX+6G/k7QcQzHXFa6DMsA87CGLVLqSKuHu5pWsGlu7Ddj7o8JnhuebmJ+FNPPWsV9Sq
4EalImiTFVxy96WjNbrFwTY1ejI38Gw648tPGbqPG9fxGpk9qVBo7w7pSmi66OCZ30/iUj+7cihh
htWXvWK4vMtv0O5n2HvT0wDUs/OGmwQujhNJKOWOMdVqKOrZeL0MonxcFp96LNDfUd2YEaYlBzei
CAXNweN2v/foWp/ycapafdMaAfpPOKtEAPC1f2P+lkb+zBg7STDY5/rqmkm8k9vgkj5N+bni7a6w
F44aH24WnTVTMnF3sl8d4zgcJTnlTw7S0MsRYbJcLjRXCrj0nkO6ggQDXF3SSqmsB7LsUGF4VWEG
MM239ieN664rvuV0JKuxgpataskaviTtSNIBhsByn0d7iTwxE3X6X1JqujPGEqVmgFimEHpUHeGr
Kqsi4RT+4Bf3ikLV85JDIThGc4DEDo6nVsMhLAU5hOosmbFRWjix21Dc24m0XNXXAF2RXQlpUiCs
CD+N0U0TOMRwiELR7ZHaXyh67qfxtgH+6Yv3ahOOGJ49ZF2lwiATF57b6ybeJQrWhg6AECiR3fJR
SyD2NTdrbo4H6QFRkSGIlUWoO8iaSxmB4cTUtAIa8l2JHhXPmVc4MfwNv3efAj/jaKRrXWumfFFz
xjY7tXOY6yRX4otS+/z9fiCcg4ngDu66nSiE8oZaNlRdodEzaMjr1g5ICv0SdD0uNJiGLNj599WF
n2f42Psm8GbJEnW/GtUS4aXuLqLqd5r6MSDZH2ZaWk4kBrEA5a+SZyY+qLS/1dNCgNYRIVwCaSdG
pWsrKo0WaTPwBrduKS4oBl673kBQguazbmkkDzaF9VPqCdTZO8YzTANMlRAVMrjJoWhRZT3fxUYA
uEfsss6/eVN+CBIVmf+bXwy1s99GEtt5ypD/qzrQAHZQnNkUqJ3YD1j5TZwAtBvUmkYO4tOo1Zlc
mvjuA44u+BwHy92I/6Hu0pM8qoyYxib4FnwelW9TDQqFcx3LWxGHMrdmSAjShV5bkoRhL8HiitEW
T+4ohcJFJI//mdRJMpuYY3SwRHo4ebSWwWqfFl+FAaI+cdxllgsl562+AsPfK4XYiu6PBWxOp/El
BHUxuc0TMj4RAIuB8PDRWmRlfup5VmQhV+9MBIcpR4JAU3u3if30+N+AmFOY+lo/07e8xlYXYH+p
UgkRWVxpnp813+3KhJEivodzdCBIQNUUhd6wGKX8GO5Hxa59QeNpaSccGUpBenrNN/KFaNAtNd7O
3NsYPXoWo1/i1Jan+/7V1s/g0dmenLHbtr4MYm14rCk/RzHd8MQmw+bkDiCvcV3ByasA3TsjUQFj
gx9u1sviYrFgeg5LTIjdSA1SqssHETgD2XxxAKUXE7SYu2W8Yw6OFJ5tguaE2U13kFb8rLtBPb7I
OBvUTA27XDPkrUy3twpHzmpd4VRvqKI4P3y9RLFBc8TVl/EzkOvUbTPTq7yzNLUuVYhj3yodI+az
KbwUnUVu/xZCszHFEQ94pdWoEhPg7IlaCkjTtTp5eVimvxGL4JO3crK6aNsdEr4SoxMyFMYjKoyU
p0IFNPWMPuHYFEdIhN7p2m2SC5VengPNyiLjd9hM9OO620p+EaugiOYJAZkDSAdrwO32TPqC1U9i
/ZJuF9qx1PnP79p3dZTDe0Rb3MqCZCijT4JtZgldjuqJZaV9QoYtL1LrAvR6V3fB9+069Vfd5d65
B80RdNytf7/xuYKAMYeq+xKWwHa9tSNr4q8i/1jEX9DOV/LYWhqCNAAYq3C3QfHShD7rolSurFCW
QOPRlMccQTgEKwudAsZYYUJ2UyrVruAa3xxfzpS1J4Lb5p3bzh6oHgOVtF6V98zK7hkBziRGCDbc
ma3SrEuFstrfiapybBbPxMzuN4LjGgrtLAfUvmwlsGtl91uysa75vGVH9FdpRy8G0LudKFf5uSvy
E1j5xFPByKegnBqHoQzjMmcoRDT3afx+z2n9lETrwsDpgvjAxLgc+waJeoCZSTiVDl1sz9/wcNoT
kOi+G1pL5KsIrmGrOeTC6jgZ+T3q6sNE8s5OJasLAder/ET+q0LqVFSVg4zRmuRpQIQ9d1cHJAmy
eT/rSTpNgmO7iHJAaF/Og+rkrHuQE/OY6QOLSr2pvMdnO9WR8y+f1+2pxNdg9Rj8yFjOAdrcbcwl
GTDw+krOv6t5CbkkwllgFZKjS5sRIJwWtLeJNOunSILPxZiOQoFuPIrnRthvEkAzP8HGqQlnDl3i
c0U0Vx4tu0f20GoJnswuGrcBqsMnXQI7fKAEUt0QhhyaLUmXHShBtk/IYqO/9Jw9ruOIOYeEC1y0
JHopW7Avta+ETupIUNVO8jKPGM8Ni0IC0RZsq5SefvcQ9ThxuFzUNS8HYFNwBGugFX69ZlvHfKMN
jYxiIY10X8x7voCdz1v6EBOZlwxJTWKO/5l7WhBVcMQ3T+2CS4dGE6OKC7Lm3cg1aQIxuFJYou0h
Owby4TPI6w0zMN8YfUf7s5L1Qe3RjYmsOnx7FIm7HYMNxw90hY5+sahUHYUe9YA3kElrtks2rYXE
5aC2qOurV5PCJcXL6n8bRlKnNwRzl0UaC04tuQWoYueEBams1PLKkDbQ0xwb89LkZh0wU4dP2KeL
RFfHBHEuLKNyxUA3VLCxKDkN5PcTU2taqLwN7LUElc+BmkjPco/aLdEaQsciNBxRL1F2ivZIlLfI
c35hYFftRBpV6UbV0IsCWFbbpBBKJXqD0ly6Q5qIC9SotPUKDVhtfUhYJ1aiWEJWCCuOR/wTh51D
G+kKdKNdd7ltGGX/s2XRa5T4nLdJOTReMQFUtFTt8XxsSoiP7nB43IF2Vj6Uyfn5wxy/Xm17h+Ej
mRQdE7ohnUjUAgqFbFG1e5IvoIo9pdDwrm1rjk4WhpEFNXGckNYMFCh3mpUD2Tedup3rxDrXP1ql
majl3LcVBVLSA1VDwWZjRhyjYQqA31D+iLdb4m+TwIN9BPPhR3Y20tXOife8mlqsNUzXH45/GUVC
SVxEDlp0WPIpDvm4LYju9fS1tWVEmtvIB+DzEozz/etJcGXJtkfRYAEBggEcOu0GSXKPeeX2ymUg
8lQUaSWV/8q7UuCR7H0hUsQ+kET8dKrGf5UO7M2DtIcXq9pkEgXKMp84H1uyygH/feKFoQ/dii9N
nAAk90ECQ9CP+Z5DP/AG0fezP0MRctFYgILFdlMCUTWmifCPKqnZRBhmh8mBVfT/6A6stat+mK0A
hjGeSPLWCuFSZh0XSk4up1eZCjhorWVlrCHyXt2cPjPstXSAusrwYFfbilFD6CJ424CQwRJgDlh8
dd1esDaO8vlBvU1V3T76JImWIuDDvzw8n0r9j0m49sNxQxPuUcx8AXmXMzWX3qhBoMRt1mSe4gXs
8u2UQZKvhvenYPQ2aWMgA0Bb1ACCxgFH9sdkrTK4l8I1P6snJV626Rb/RxCfUorRpiqimnEaSwoJ
7pE4Zm4ck5TM8ETEfa82XUVYUZzxr6uedoVowgVxvzH9m707TDULSNnEdUZxi+zWFnQk0079Ll7g
rFG3cSbosFuzmbWeLa+uON8vIKVuxh3o3vFpOARG1aeg5+H51Jsve8cgcpW9R1LrfYICB9i/NZo6
hrvxyl2Cje7iceXEczj+J1+4za1DcCVCz5j/GXdPrD5CR4gqvjRr4IzPEBXeZKzGsI8bfNr9fd7A
P8PXNKq0mi6llBbk8yZf7WhAVycHIfUURSIeAYKFIMIP5betA/WGd/lOLL+9RKr3WxJRFnBLfPNb
gJYGnxgmsY43tvQmu/0CXACJB5ShfjlwMhZVjQ/3+LTCQ9f4CDii45+0TnwzZVay9wt7Qpqz0X6+
uNDk9nkW0Xgp80xH7wk35uyWKdHUJDOPs0X7YHTjLg01crjlwIbyd6xIUnmmytEyurMLMsYg32/L
4zWDN8kPB58lylWkxp4uAS5qRzQyjoO90RKHmcIibJO1V73LCbRYq+elRMSlZLU514yD0dVq1YZy
R2YbXxOgR92g8VTk1SuMSi2uf6SNJ6A/Uj/c1XqDpkW75ufiASFc8GDb0QzVuJcSdUcFZe6RkxOB
ZHWHqnuUm9xPLf+Br8fb21SmBR/SSNKhqefSO2eY9bRTadm9hfpWIkj22n3XGbny0hyecpDyUjYz
+vQhMTXFK7FCXhkR3PBzBYNlPNP2XsS2XtxiBqT/QaH1SAv7ekoso8M5JqZQC/bBCPfTmKNpcseJ
FnQ3ioBRaUvF+HGnpU6jyjxuST9qFh8787dgfx2CEta92A2cTe5V5u+5t9BxteWxCElEbJV1FQVM
Yq2oloFN7dC8yZ2IY79YPDq/7/ms/R1Z9UYGHzCAJkf4Ha18vNBS/7EjrbdepRM3cCmwb4xkpD8X
M7ww7ujqgWteYPr0SjIKwDSXZjO5YMq7VYgtqq00zsau97twb6Mq6K9zn7bLJH3Xz+MOeF+4+ozv
suq1byLnK7kQWhVsEWtnRXRTfTXqj3O74EVzWiXuKthNEbb4T4xZRJ5ENx0L4cCnDNgjJu4Q9H2n
8yMM9TV8w41qLyLDwMb8NF/RyDFdSwOpuoRgQQn+lciPW8MfBPPjRP/7PwPhloyanDrXDqeAycjB
u5bLptK8UU44EQkcdlhhz/A5D/nO0SDr1ABiOr+EqeRnKemgokJ/E4nnIVUt2nFfK/U1NJkqILBU
Yk0MhD+FAWAkBdGSJ3OKITyslGo4eJmY3K5EOwViVM9Ori/JWyQoEa1xJUtGTZM/NLwgeUGnwBW9
koeDKNjS0OfU0iA3A7qMOSH8k6fu5ZFdq3msJnoBr4Uh77vfgwtUczEjik61RotLZEnGQ+q4hoWM
4TNWz+L46ysuFcJGvlT+xVi2/uN4S7+X0mHvDVsyhT1CwALJfEC+Or1NeNNzfkOREEIRYqAjc+9p
9Kz7SosXPM7Y+9h23VjmyYtoUjO7dZMDQMRMjY4f5wLOiom4vLLBpdXoYmsv3UUc/Lc425ZNrIgO
QRl1V7T5loqnJ0deXs0ezTI+WRvEM/duXsxBpYZ2f4a3YRLMyIh033QzBrGyTDIjTwuOYcpdGOOF
BoY+md8SBDbXVC+zeXIiCPHhHjbyVCChUwg3H1gGWiGj/xhNuJmDhvazykJvR/zyhnEHHXB6gl8y
wbXL2QKH1kerWbJbMNJLKvbXJVax7p6THWNYeT9UT3bL8X4iPjtxDI9GaeFcIZ0j18qu5Q60mVvv
R4UPtn+omxK/2i6rPrD1O34riP2fwLloojrkC30FkflCI+2NBLyu2P5JeuudLpbSwfBKSwnM0tpm
U4UkzocXmGwih8e5yFL2HQkJn6jcKRV9ZqE6UizfnDfmnHpgOBDsni3/YLcfMFxhwU5XF+k0IxOF
Fxj5KrY9XEoNj+mYu2Zn2reF2qOGAdutrAEdOZLbnGJIgEfPgxKG3yj3okTMSA7+kwVh9o4KXvT9
FOLzAOrfbgQAzgZI7z83HOEshrqBfFGY0mN7pmR7FsxHy9y25H1uug8L3NUNi/GHZWzoEPXUFmN9
xxbcretAbfZVJfPSUB2f2RDp7+iMFrKUmMbbkHvZpQ9yKBt/Ik+XE1VJ9mBSuEV34P481wml/8Rq
ujjVI8Y2qrS8KBkSvfJzO0KRFB68PHhYLWYO2Ff4RNbFSil5NAl7GUBUD0d02APGDHZmVtNwHnUE
dh+Eihp5dqBEO4o/KC0tGyVn//y1PbcW+dYHn2x411RittpKNV2KjBAA0GtO7QzpO7Js+7bsxZJ1
5gsUzEyS2/rh7Lxz8GcLrTbhbnjiikVGFvF/x9rnzHtJYNj5a8oP5DQ8mlN6art1E4pqAyUazGIv
dgeGuHjnOoaejBHDxAprT57htpgJy1WLzwHHVJM+DjNvWArylkwQbcWmtXgeEV9/tb6mmfbA4NEB
t8Rm3STaIRxG6IDRL81133NRNc8xta0VPCVMzexrZB5Aj6zdiGigYSMbYTBYeEL40ukViNoyvQgy
9K6iEUo+xn/Ak6nM7e9omf6T30NLECplYsQAhC8bsas6zcwx+e/6b3/TWEejqRQ1z9pRm58Q+6H5
6j2mkMLRJ2KtSpQpJiurG9p6zUlJCqiMqUwEkeFGNMBySU2mf0ryo0FICTKJMp6gCAFiOa5FUic6
jAozTEIq33v+W+7219rFFyW2l6r9pNIx4Cm9MrCuzr5rVlLkRQFqJMtDheCueUo5Q8FBl4JtbiKF
zkokRYqEm3Bw7TzU722NQUHRJfHg1FBbuqX3Ej1QrohAZ2z+FTSXjn5sW66DWC+gulye/5Z2ALyH
I7KxxS0Tr95ZaTz3Wo2IDN4fCarcpRixkyYwHmRQ/zMlZA/AoP58zGrM70qNTnbDQ2NKgegH+YxD
wfLBk8GPIM1N4LrRmUYvAQ5hi/Nr335zF7FWS6SpxCD/ENXLZgxo76QPv51hZx4GOXl+hEnnPNb+
R7mixEbIRSRdDiEAUD1O6rnSk/Vcr7xAzMNZgxPwu9xsAKPdrIfH6VsL3n5cJfpt3Pyi9ikWhNEj
tsIrwXtlBj6S+s8khKERWk3hWkb0GCiywMbOSu2QS4jadRdKSeAtxXdBFOTQHrYT4zBpGP0VAtC/
gvHS7UNjqtlhi8W/3mOVYMHH7ov8atEJQe0eD+LhNAVb4MKSnEf1DR62m9GWo6E40oPWG1Fmf3oU
/ndIq9qzZRLCml+6/NzvYJb8H3AmtGJkPR4yv6DrLb/13Qc3Zfk7EyOmwnNXc/8qVjlQqFRpcvUc
SDdzhYLSv+K41hmOKwlWygz5S9Jj9AfU/RVsaU5lLpH7hyQbfq2BgREqUkOAE4lcVcTMVCZ//lmW
NTKSj0nAEUtOic847FXlN+dkdQLm/Ml9JDti8x4s6nOCgaEdm3KG9Ghi3IWR4sKBtvOidB7D7aeU
Lsaqixflnbdh4a+5Ke3ut2NTiIfNVG3ZWnLlHHU++7iXPP+hIQfgPDToyfku+L1V2JyiRYzKKh4Y
DPS+6HCBccBkNOIECcl/sYgYwbDskH71m8R2UJDQQjS41HdFxOlpqNPtJru1ZOw2XWZEvVZThvj5
4KcvGFV+NENia0kdiaeB6Z/n60xzILlyYWDLcmczQYrFXxgQ/ORnDCw/jBpSFpAjnDdkG+Aczbmw
lAlpVIvJMcDVyr1qdjKE41RhtTTFnUK4qY7DlIcPPUMKzAsQrg2n/zpFSq/EbL6mgY2/PangsSa1
tSDVLd+05dBFD9WEqsTO6Szuw2Hsi2SWwHOjUWk0dYZ2lKdyH4kmBbT3AuvVszkuJqtJSefQjO2t
AIUjUDM3gL19ynVFxhLtuWks0cICHGoNhnhK8IsosR8n/FoZk5FiNKIcnVd6e264K0JwK/Nn7mfd
o5nANSyrrl/K7u1Xwj6LwPstjCnjuxJpkx7Geg/OZCQQAfO82pjqHAppw472LyPgi1O3Rp61Y5uY
aBsBDgQZLH+i8EoB7hTH1h1lYbiAd6+XN0wv6+pP/TKzWyVQFifJGLEtiN5yXSP8qkcDKYIM7FSr
Vjc0mvVN46O1MYbLGHVwtMv1xbhiAwxW1qSJc+4E4/b8fWJ+AoQbJwRMzxPZlxaoXfIKSpW/nLFW
7RFHVll8EnfOAcwLjU7bstrQ/IpJCSL07zFeR6ytM0Hdln8dbpN27L1u6zT9on5NdZhP6KszC0C4
BVdxrl0jGM/FjxBTH6TL5q/9BpSB4DGGaP17f87pKH3M6jMdpQPJuoS8gse7RQDx64ZItrJ8coG2
D5yPDJaWzkQ4eOSIYyD4a2/BvmP3eb+/mJN8mhV3yKJ2vNwP6OAizvUGxr3i8RxkHJxuLFvM5Yvm
sC6kb8CW9Ga0mqVzapXvWL8RLuTrP8/KS5tyhGSG/sRlKp0Ad0jqIKrhouCQw6b7NG70LS0gPby5
0hY46JfYilNVb957tVrLmFwwXvB0Tvxkkymafb2tQ5j15GDlaiKO+FImxxEFTlD1F9PkAE47MTu7
Nzfa1F86yIdfUix0hXQ+S+v9Rdpw+nIm5b4OoZX4dB4J5gPrwIKW2hvZKimqwjGBeDw8OzJbVdik
gmtKtl8v6Nivz1qu4Efsb4SuciLM9u1+xcw0FminAZE6SKss6GQyVByzgvGY/CAu7sPZvxQ4ZPRC
EZl0/ukiZlkqu/8JBFnfcAFR3WlcnqDML721+WpyuT0x4tIOhlT+I7Db5B5p7ftWmSpDCGhC2AK0
S/YFvbvP/GYTnvxAKrIWVjLXG10fn5CLyYDS/64ohElKusahsmo9r7bC922e7CiQqSLdMSPN7AVg
2ObpJgwHgtR/uJmMIfOSWp+RvMjgUjdyo69cVVnGSDm7qH+6XXxsp0wpAqQwrEKXgmxkjaiBg7t2
lKWEhdWXHo7pgbe6rzbVXpc98Ca7K7jTxqPyUGM9DMldZDzmH3OEc6FclIuVWf113AfHboCU8Nz6
IBvbuHzwEugwYywJOy1HnuEvhWkrVgi9B+4QKyMaMlCp9PsOV0reDyW89Ec91mnes8HL2EMmJ9fg
1eghX14UD2kGDkUPHMKFS0B2WeEs5dvOy02cAA/yxWnjX+rF/Ue6rHX9tpXLUnqZ1g7k9Zz2eDtU
0hJMm6vWKrJmDpRGb+FwzQ5TBT4Ju/uraVb54m6ChsNu5NiFI8YBcQ3HheVLIEXzwOoAHqeLDRLI
55QPUYXL5smnAl+MDajytGbCn5bz4TS5By2Z+0+SJK8bRzE3iqdaDv5Hby5RXXW/vveryetm2G8x
z4+KVOvdGW5qGp0r3wlT0rYfo86xm38E5gmhSzyB4hAWrFFo8yWuxVsKI3vMTIe3x+bRmeJmpB7m
v7DSAjKxOCzqxZ6FU48d/KS+o/sitpgRuB7P+Pm3B3VaPzhraN8wbFGBA6Ng6JFG2wVpwecvzgRk
JZVa/rfsz4qrDnHoQjlQaBxJ1eDDJKuIAAsMhS33toypWsGj3rzT7NxBiTNbIB0nbc+jyIutVQBq
G/dG6VjfxtmkqbOUe0ZfgLnPjIL5cnKldj7erNyXP7HqN2FMaBQ2kaJOzHgl63B5bSAeIjY+9V8U
qM5KGHQricpNtBMHKrNutwoSBPgc9mWd7iIwwKjbtRiRIw3bsr9Ca35PLxdTr4zMn3QuI9/+N68A
h2dPZx70JIXlh8wphwjxMfMq7vnKv5DlZ98rFkexzE/RQ4NgNAx3VO0JgXgBnxI8jtItGyWMgp5L
bXrFZmw39tFqiE6HSFcgPdSPM3hZwHkASa/bW5ybcEtJWnsdZWRwH6rRncPlcL37sbNSdp2yzil7
BC+zsSOj+buTQ4d+R4JQ7pBqvuGImm8RgdVK5GlP9DuOEe8wMnaJUdzrFV5k84zDCAMXJc+4xJzw
v1lYrdu5/3kRgFN42aEgFqhOHpbSYoGo5+8TH5xW8sjkSkmIIiJ/BBUivB383EAoqRftdl6BcGt5
Qf8FoysYuCiRUqvzowO2SQ+LMATIR96R7k831aIXP4XSMXExThmud7V0HkXyoHU5AhB5Dt0ur4kt
U5AmspgJ6p/lqW9KeATuK9mSzsokgqqLH01dvwE/Y87m9QFWFjh9mJKkM886NbJSxNm28dh71IOx
4oMYyPEZhEbAAm13MD1uj+ozvkE5Dn2RJqeI+OwPITLfvJowUwBvugi43s2D2FJpW+YtvADd6tmf
s/M5Y8FlEqy18IWTIp5/g1YuD/z6Driy2eQaQQWFEGuV8FIPXyLkFisxK0Z+4YbMGkse0jz6Z5hY
ASwsb51tp90TBsRrtohW2zMJn3KQiYbNrdfFI8hDme9rlzbUpj5m67TKNv3IbghSOWuufD37cycB
NcTFHM3Btss3amtUvAUTLQPsJax4Gn0rIV7MNjJbE5BZ5haP1pbK85tU6i69hgLt7q0VJjH5PNLC
w2RamtIIDYrLvVKICmHbbOxRm8GJ0UwZjOk2ZixGDuew8W/5L//LK6rY3Fuo+Mo6ShPJZ4FLS07l
GYXZeBdDwUxsdkzFdOrTOoQD1SvNGv+vIMYtGWg7HlX/hKINJuVN6cMIfHDQf0rARxEoFrO7cHiQ
Nb2wNruhF8i4edDQs/TCPoTVSzVouo0GiSecsdiSxOgy54nMad+Mf99D8a5vSAech3Mql0S5LsOR
Qq/7soMP+a0FcHcqCYWECJlu7eq04rYqOhVfEGhAa0X/KbfNjao9C3CeuvkGLLVYdh7Ueem94cG6
TIiCzkZ4K0XM7bKff/CmZVNCAxWUAWjRI9+A2wK3SrFoCr+clYYGE5C5Hsflb5+M4sTEBxOe04mC
+wbyMAAVsCYQxGjlmS6hS/HPzXeWngbrtytFUp/HIQF+wUu+hC7SufqLZajDQ4R7DUyCt0G7+3BC
IzBF2jd810Rc/Jm/hR+xt1k4o/XxWMSYYWjqoBzOtVYYUBQA6v3w6lVvLVKnep8q+KWHEJBpgkeZ
V1yM5GyYl55pD+HwPKSdIhvCd1bu80NwxPgCvRa5qISvSq+XUyf5Po8ei1K2+SwZ5ECNVHKd+z5A
vbn14bL9DGAJADu1bZX2AHiAIJOTQX5tw8XafL0ntZtsNhETe6jnrClY6I20zRNUHi45qESgEwq4
iu4ce2/SuDeq2Hovubyj+IpZm4NA5e8tD8OgHauumXij5JdXlXZlaRKjGRFclndmby3Z4B9hMUnp
Zqq3dyd6XrfOWeH5bCm67a4Nuu33HfNkPUL0zsd6AxdhkpUSXFXq2qAUrED/RNDv2Pl9Mt+ZQlIT
b23NqhB2hW4XhHOhZGC1pUzjKckx+BbB4XgkpzPuonZQJaJO6gJ9RpRY9rSgh8VN2KM9DZTXO1Nn
Nm4Pj88iWMSEj/oSUN1OuJ3jw0MNkRFQGIjwudyL1PYmutf6WsoTvcrU5rl/F6oI9npen/KHmed+
YHsz3YpCwiSoYk6bOuoYppYsXB50KbxEVgFZgHlD3v01uWAKeaiqje/GjzsSVu6xsJixeyCx2Nw6
8Mfcd/pVCW74v7yEKUAFbn50TucAVviCEZ+u8VKza2WngemYHaGOWIhBFh//rbWXhO+aVXmGOfNi
HR8XPbj0GQMJtucrzXQ/Uu0pubHa1GnjXIsq7UNYMn9SAF+E/63xfjiUsr7J8Jtp3K4tJzfByR/0
e5YQ15RYyMSsIzlLV5x+AuxVcXsxhEP6ROW/BuBReAe9pYu4c6eBJu0h7kYyJxemC39DgddCewXs
BQCWRHx1ZX8YHLLfJCpaPSP6PeAVGKwUGP9z46oX0NoGDfDEzkJeHk7CFC5jRdYanqFaoumgG4iz
jWosRADkwpDse14WXWj7SgI1WWTDyigw81NKLkr2vXs7qEO21geCLDMxOYSxpQ+NDNpXKn6Qy+dB
BSfsRAJ4lwr466wDFoO0s4SKaRPwhSu+O0GjnYc+nMuN8/aTOMYMqSZsMUsLraO56uVK1d8qehTV
XlZlqtMr62SI8xFxjskRIlfIfBeMqt3hhrkQ/e4CvsZWLdfij2LclaJev4hPzMe48L3PdxzEXsqK
p46jZAAYyiOW8jMvnfmc3I4fOehi/o6FEmBhOo66KG6VNZNveqFS25uyUdv3VYDjBb/eNQrRWwGq
NsOXNT9wzC5EQAQ8BJQVSMjY8qhLH0bNklWW9SMJYt3k9czeZutoegF4SEnG86GHS+CUeU6FuXoP
6HDJikctg1pttT7FQIyAt1xQ9seZ+LU3E0+bhDtI0Xfyfe2Ni8WFJjuf/WCGD2KZx+1bBjgTrJg9
RiHLpjUloTix8b6ZEdXNE1RRiRZcOIten52wxXd97qQe6ZQbSQdCo9JmHuGKHdZEvWXCIBHLvlHa
Y90+mE4i//k7cfBTiS2Rp3n9CIWYPYpgR8eBFh6R85tKnzbYRFdtUvR2iQrh3NGDiTtGYKR7qbg3
+pewnQXqRyW/LGjneOAFvlFoUByLyNxEaGoWL1S308DCFW7vg5RPOh0OzTlYeZI2rmCyWI8SMso1
wH6upsNEChSUlYjnH81/x259dOR6xLW/BHOBNZLJnqbiR6lcTJz3vK2xwYVX74MhcCMQqBkQR9pQ
ON/9tohCKMC+6B8SzlBonTXzW9gnJ9YbyHK8M8lsj8JKpGwBA5JwkB5x77vd9c604zsGfPF8Ocsl
1oG18WBH4hgOKcB5Vl02bLlQJY94ZipH9EhrF7OIDdy99PeG4jRbvIW25ujA+wmSUvLkze6se391
oxlFriEetG3jLyhkQz+T4nT0arNEAuzMnJ6u9m57ECkub1QZHXotCE1cfhAEb3+HvfvdJSjZEfDe
xHKpjJW45u5nCcDQ3sBFXNs2VzFXhfdFldhVfwhrJwxO8KineRHN2rWTBE0c7Cy4J15yf5EuQ1rJ
T4qnO9n5dRGM1XupjHGy3qB/3hefShUcvp7vbWcHaLy1xamyr16MmmV6BwEe9xVmTBpAZCekAyni
AnmEJlfc86nZ04S6SuJSfZ89QO7IYkrkUSeNRiq6WEjxJWh0mlIhW+ubY5CqDWOJ/8CTspN8tQ4l
sUUUstS3Bi3p29U5G8H0dOOpEFujATljjvJdvFNZlXJRlHtwrKFa2GU12yGoGM5NuXktVUbsHQD9
NWMhoxWh0AImCAIw3kmFPwn0ph8s0WiZs4AwpV/qQ70CW0vbdgIXs2bn0IaHu7qv4sN2Di/A4Z/J
71a03Ym6utHdYgJpjJkPVYexnpmAOIod+3xUG1IwWVVD3iSS10Uz2/mKmJ+CMQp1sw59NCRhQ/i5
rlK6RxGas1JU8/MqiseS0YnxokPTRL+gGc5EGimpKkfZYrvNYZd4hG06EfU8/LhuRuay8ZbeqrRp
eIE+rZh3qMTaE2j0zWrWtrNPurqHOZlyOKsfngf0RGDU7dwcsGrXGbFOPZfIglFoCqSL0K4ur2yG
DF1pz3jQ2ZwSL1qyt0xNza8vfOVBaItd6o2xnP1+bhZ/qRTTVP2y9OK5yNQCKY1HRJhdVi3eu8RS
oDRNQYQugdT+eD+NGvLTp3RBCrqr4+INAL9R4eqxBFOaWLuJxjLytqGWuA9pQhmOqbnUdpDMrvjx
E6AR6SAfabLms4/ryL6qrd1VeJ3M5cSnrqJhrJl3yCagv63CQQqkRQJYPOM0gdJmV4QNGGOsiXKn
/xOSYjJX6Oy6wsgwBXWwTcBzDvny6qhCr8rp42tFAoi48kVRo9adKyHyWfDUZcKPFNTeCutzOQ6d
P4hUrAXs8B4Q7B81xegTV1nL6HPG1BnA5rekHwTHAedNbz9O0/QjJq4Mq7/ID4trkhRZZYacILiQ
TWtmbMcP6w7eib1qa/TiPqN0Piy+5vIq8Hip5jX6DVqQAiLg8KO1w7uwbc3eA1OxqBcvJJbe8V6w
N3j9BXtTO8mB8nFltz0XeE5k7bLWiYVLezyxoUx27cYYVS7svgKFecgYdOJZYnF1yaBR6av+YcSX
6FJqqvMNoW/IGMM8dAJIzboUYRpD/Xn8OP8pSzc4ZlYP8b8ipb58qDmaWyxrWJx6M0ktLDN9bPTx
C9VKiaxeDT6c9c8mfeq6jDq2bhI8uAB4bDr9MnQO5AQcEkIKOo5mFKFTqr8ZNYbGPINsWJv5Ajt5
KZbAq53QzMiW6iDMNWHhgkLzqOeyhxSAn85Sh6Ms0QzHoqnkAbe/95r9aqzXsBr6iEgN1EC1rTo0
WA3HTCm7IIzek9aag+6AmxhQr53sZWhYoR/at9Idkeg89FSWj6fuYUCHESOiq0aQk6WKCDiC9S73
Pfd5udPyW+kEWmCwPcQ2TSqvmXyYGF+fgRAR+RXsDRb/UMNFXcr2jyumLLOp5ToyBuWm5r4wGY8s
kkS9VmyhlkmgDYRdBi3hmq/ONlcBhsdvlnnppWSg+VS/Y/3wjDG27niF43rxOHJd6KjdU3QyA+zf
986C9yvjGaPK+Tq1GZS5fSYvcXfVZggki8B73wrXzZVKTFJvlfCjbdX3xmQq31hZq1PM2TQeUGTj
OthkT/6zijGeIt+P1WAQPFKOmef2CoEvz1e2Hl1jVDE8/4lfgWMUDD2kavlj4Ey6sebxR3TwpIj6
iAAO/hBTRx4pj580PL5oO5vNrPaD9E008IAPmwuSRJAQQuIlNn4HyR3ZlM92vWK8OOF/FzeXjCCV
AcEfxzGEhK42UPyT/XCSrgm8ecc6FvCYmbo08i5me0P9k2M/o21wI9u/v1wFFWzoU2/LFFbB0mIJ
Yy1U0Q/j8PMWxtluFpOSJHQGg9wAipgeOPgKXq5ZdR2gvoldy4z5XJK7LBQ2YSWfBgGmJLfixwEN
hfwEDjGEmbewTG8pOR4R70vBqOF17QbZSIETSE1PtHhQMRqsnnkA2gkMvEq8gB/9GwUEo1KYhWUl
AD4NAHtf32F9Dojt105T0QlXSuHfycL9G3YeQsAjBB/6JFp1Llm2UjjW/zl7lL5X6CFqBJCHugyl
GEkmHgDwomAJxBjy0HpOc0QHi3jyvV66XtoEeYbSLhgBFjT17nJXhakPO2PxKeayOUdgSX3wQ7Dk
op5IFHvpSkj7hLPKY6RYybS5PVi1rOYyfhllsAgppPz0ezjYQKFlLU2JwcOYD/yB5j1zjkHvfd9G
kVhl0EZ7bHPinTkKYR1bzEONwoJky4yTVxFPG3f94LrwlO7v6kqy+NkO530J21h9Ty1ZHSfUh+O8
FMaO8ab8bv/tdbVlfWIT4tzaizrNF2qrmkwPsoE0n5mD5BMji0VrWcvVWkB8q1o7edAEeH+ozsvQ
tgIwMwvUVTFat5JtfrTjRysmRC7htXMh74XNYLObud5lPNlwreT5WzPcdcabNaNdjJvd1UG5VlMV
qM6jMIwt3Opk08zIJ//u5eamFmGxXiXkkKAZxvs+mMGsGegSXLN+IyhjhW+R1r98XDqLCLinFpuS
4jtgP7pCcPGO3KTVsJ9ThBD1djWuQuYIgHe5W2M/SSVpWMs05xggR/1YJhOMzBpuMqWPq51pS3Ve
DXByeExb+g/BBbiycQZQgeR/gC9RckE4Q5OyiIHv2n6acN4RuamXAdAkCuRijdnybjJ4RX6w1+Lo
hvwqolYmb+2pdV9QNRrOnV2Xc4FBwMud8TDhjnFIwaigoQCNBADSz+tDFGDEaIqx6T63SPC2q51i
NQltsxMu2kjkgnwzxZxWQGwjz6/KuzRRayOM9+UjD4ltEs9eKZPglm+9tBgP+dNoxuwvA71R+3U7
AjjUust9SJPVC9O8JgGx5FbDwqBVONGABmpzXIdTdl1KU9M80E9WXfhlCrhqmQVA1oDJgJXS58A8
wioPTkvOmza9TCfY+D1HPo8FGnFu9eqjX+gRr+FtStZ8DhQWcCWPshLF7ETLg22t82OHpqcSHTcW
8XFfrtntlAfdJ26eMiJAo3vJqVweA9GvSjyiVYN2xVz9wnhx9+t13gli3awUTBhfNkaXqJxKM2US
xZ6CdvpbSwFulKn580y5lQFKsGQxONLMgWk+NaBsniW7FeOSNC7GRoRQvGkSXLFOk0zHhwNY6rt9
bok8bDvWr3EzPBSJ5Upjn85JsTWKbpWw+DHBe4Lv9CZ/UASklPjmnoTYgGt3RHfq0rIvOti+8wsH
jSMQ+oZr4V2yqGf4AqlndJ9BXg4X2M6QW//VPt2lShPPtfZHw9zr5Ump7H9KVpIz8gYMLGyMIax+
bDyIONx9QQOEkzRvE1Fp/UZZSGH3wQ93+LnPQ4Knpdrh8bhvVn1y5cjjgt1UaaLivx47ygxnI3AK
rIdzjo1261dt6Ro0rmuYJY8RYlsUU6ywzOG0Pt5xnjSttDSLZNg0RPbfIrh0kNPzAcshKTzA5jou
8MGM5mbkeXcx7K1HlKhfThQNq8CyxivFwQp1ybxxlC4WFi5rOggtY7P1K43kwlGUIKNMSjACRlMh
czNUXJKQtu+aj0akWz/5KzZrScoqrBwkzXtbJDUT/lvTzLUDezjRorXM6ZIzrxbgMXhFYA+jKjO+
UQRHOyMQfmBnzQjDTM5xceowUjeS73foNJqDUVk6FltgfHzfN2N4eKZTdjkf0pmavnp6Lp2ZSHNU
fetrOcwsi0yp6sfr6ws1oU03z9hojirKplzVW+/3h8roslMga0OO14HdWuy1ZfxvmQJBqMCMfRpK
BWnikT7wAwC/NKbExAWUIurX8PR/M7XO7tJPKDQ2aYcGU0+0hcK8nRyKvZ7y4HpsWqWV1ldseUUm
OQadven1Kdt/T5pwzYg9XwCQvoQxGgozblc6lMvV1jwjyYdHvXVu9VkhNW1n0GzD8f7lTn8yt0M8
IH/lI6HqL4Mng2HDzWpw9P1wZlDsKAZYUlQAgamZAQ5oH+Zhi9FFYJK8SExTKGs/e5S4e5TtQnZ/
yyNx1e8glKMoJ6ho6EMYxtrXbHwTW2Kd6qGTiem9ohhnhdcAMwbY3l1jfTf7P6u5pAkwrN9IiTts
wBrnNe8pBiTyIIIK0erHdzXwsnFQ/Zpc814lkVhoHqRM6IogT97w+J06ceGE6vld7+H3XE/DvQ5K
CuCXLVRc2VCbEjgxEKquO8Y0flk3i9oVY4NyPzSUTxxNHHAXnQyW48oXjQCGrPxCs+clmoUMf4tb
w4tqzKt0HSTLfE9KWbllADsIlzKtjvs3pkKlOWbFjGT7WHKdhQDKmEUu0xcgO8/3zWXuJUtEaKAP
uItXN6+0LMcg6Vg7K+QJzcATt09ow5767G2TaGAH/fqZAJb/z478U3qwHUxTAEmKqK8mTff4eV6T
ZTY+Ty5P+t6bGu627SXvGpBYlNWUA966N8OR5WIrjiUyTjkT9uONtK/oXiNROw4NRSgjDAsn1ze+
jhDQy+zZYLk3J+urH+bnBZKii7PNUStZElQyoIwH7W5GxTRgRZzlx2krsGC1FLTI9vfpT//qhRY1
XBuvmqwz1CrrI1aAWXCKhvKWDG0Cp/0oYIkFd6F5rMdAb2sWylf1Cxu2a918tOk0m5712rl3+9nn
2QYUN7Ep3mjkgnz80tb2fbRUaR7mI8e992X6963Sal/wIWrcolYEbFUKtAcXLC4RNDYohRtFZvcm
gV45SgL5wztb8nWpR1fzsvvuQQvaotbd7p5mIKpsdSBfbmpUPoYumkUrh0jt36LyHKxSxakIYYqN
8l6QLTPBsWf4Hg28NL9Ordek9yAPayHTf2AmsYiD+vtqftx4dmU/4yKqOw5fPVjax8iGoR39AKC6
I+qkwJdSgmnUeTpWCvJ+4pY41SZK0ErUHwWsqsVXVZ4s2cJnlwIKIQtwyEELAuFx51hA+Xik4KNv
E36FTkCcoav2gDXrxFvcS6p4jvvJ4cF9kuO74b80xvtfk8j6jJ+wbv4g5yw6ktqJ2gn5X2vBxMyW
cL/PEcPRxjS08mym/ZKGCJTUeoYSMz1VFJbEL6dU4+L9n+Q51aeZdlLOZECDk8eD14t9sH9RlBQ4
hD+goRcUj6n3BCqVWxCRi+8obWD7tqHjsXkbtOoMH+KGZo+r8C/AKYOEVFlH1wvBCJYMGqT7/M2E
J475Yyri0GP4GwEbFGWEEnWEPvL47ThDJpPCOxyz9Kvxo1F3EyiaEmKymEd0HKgR8rTYrSdr4Vbm
yUaA0L3ztAwfEB5alENthCDl6ns+UCPWdPqOfrN5Z+Y/rV/CZ7rPUNjWBRlCVocezV43mNOEDJyq
s6WOdZ4dTHVqLuWTugDQpZqxKuSi7XglJGdGceRdCAz7VPlieQZcB3uvax70JA2jSg5bOKbjfthw
xHVQX06YezrTizVV2TfAXLV1T0pn6BlOCbqFfW3iW5BeHwHV/8o4OYyPvRZ+71Cb6Tkq0w/ChgLV
JDQucL+xhCA4Xox+qrXIk0hQwGygpwBOf7iaQGmA71TPJk7b32gC1QSw5jYSQB0MycwxYaBdqi4w
n4uNi2lCDa4S0W3Ak5B26j6jaPdvFlWMYNUkNYWTvaaCdDbo9Ll0Y4SmvV2P94pKTmYcuN4c1yLM
OpXeFXQrdYbb6KsUhk2ccpv4wr6DiLK1jeGLkigHqP/Bpb9vJ9a9c6hHho7j9gulPpBaXSj9bHP7
yj+OG2xkOEr1cBu/dS34IFMbKIrTZZC5xmTIg2s/PQoVY8ZC+4qm8fQqawTAvGpsygzLcnv+t9X5
xJyUpIbzl2XUkkQuK5uXk5RID33YTCBknjic9BvY7KSy+yTzmF2N1/stQVbjHbm6nhhaVhi6MWfW
/LMJ/lxy5nsz8T2cZcmkpvgzIyqo4P1xGsRVlVVF9FGAxdioG5nTJPW/SgjiEmrxHFsDtLzHVzhB
Arb3MTC4nrMeBgNFmjz7S7BNU0T+CL1h3dQrfrbsjso1pN+nP2OurKz76umy7vP2xCRbuResdheR
CRpGIku1C0IzXOjVAUaXJRTQl4sxs4An2Cjz9zOxlbqBy5KyK3bKqeU5F4Eb73u+765pz2a9aQ5s
CAgH72pQ2qNOHl8Uz1OeWpq/iT6uO/LVnfTOC4SPasU/V6xhd6YYTHmlxYW1U55M9Q/Bzs7ZYvPx
z/UdsBR+YHRRMdvx/KiEX2zCdkAkxGsiJ5Gy4N6hWB3WgPcnfF/VM1YjSjWmh79J5joyPhEPvloT
Tpg0Y60eSpfPLBHuNbm+k5qwSY0QTZd9k0UxA4WXZy3NnIm2P+0PvtX9R90stHxElI3sfnGrrm4U
t9435FCO3I+ZP0jBZki+RTOGmVtqmtMsLbpTkTJ99XAxj8IiEb9MXPGmB5OGBZ7AAZgOko7AQb1B
4yVUzYPYX3B/XG5vqBalEn5seAHZ0fb6YjGxRjhDW78fA1pP2pEE/bj91V2r3c9FGAfErYieIlCQ
I3kCdV7WZG6oPa/u2IXi4/FN2/pJKAkvTwMms305IbllOonrp7LYtvEiZiPv/zgj4znpKBSDbL+E
dobcTcx67fBmkDS1bTR/3v6D1QIzJ3KGMWekeOcUiGiY47IJNgkZbV/4nqrXfSGzNusAjde+oTwF
Y+TZsWaFwin/A+ZkuD9EgWOngvocMu8qx9GYrI7/CooeWMB2UQrnUjDKOnjLTUXZfp1zSoy5Hwbc
C8DTbLJBEFB7OYICJU12oYZslAGGokdTngEXpqrWI66AEMKsEl5l32aln++S9R2O6d+U//FZxTbE
c+qssX3e8QhYKgVK4C22q4inOBcjZJXxLt7jU8LdIyKEY4nwcXQwUQxo0SxoIpx+6idQoVaFpsjF
cXooYB6lK+MpkmU0eDSewjFy5Q7qB6NDevMK8jvtojL4K/qXJmN3+gVP/d8OqAuqHynasM1+vtFB
ohNie5PchDtfKq/9bLXUAEwqxCzjcgEWaIvL6/OAiNsNfK1rEeQ9NEKJBrP7ib4cgcM3Fd3C+H3V
OO7xNTfjfdYKtfysTID7kW8YkTb0Y+dSi41HDiLhqJy+BGH26OEOWuvF97bvkxSlOOWmY4t/waSY
tPkD6VXhhliKMbW+TMI+dkgNovPvfFMrhcuYbHu26bjnN7xRbQoh7wdvj/2dmhFBDIVaaxcOrkc1
KbFie5b7OSGrzL7TM3UEMZoo2h5fYSHQOASk25uFFEgU7TL3KhuQvUCWNa1fxurhSZlci/PXP4CZ
HHIGt95AyIcPuhv8WIeu1nSdJa+HCpkF3LayvyAGSDQ78P3UmYClBwE2mGwpKuomIXz5vRpOkQ/W
VrmmOuQ6727hcdg1/sUABdBFoUClWA7CkeG5DSGrVFzPFX3D/mx3f252Qhz+tY4pU9hxtHiiBNAP
nzOZeyQihqhXtYCeIn6uRqYwv3SRy7/lwDqxfzQDEOFNLBj/gzbmmnb6rEXxpAe/6PcCnEEixSx+
uHMCpnxmFVGqSEfcNdPudzUE6IE0rJ6MDOBnVdVoTai9vkamO7m8by+Jnbap9Y7sGSwt6Whi973Q
K60u5RneTomm0UE38vldRVqdkQ2BMQR58teXv0GzftuIjv8fRAf+s8R9W6q4ocOlzOlecfeOiQ/w
qL5V6Nm9pFz8ljPmi3XDTbWAwYix5O/GsG+Mgj6gdoE9WocdpCu7xo8uwO891oQL7e3cSNINOBsD
NX4KoloiOOhFMBdZ4BMx014HLzvyeimrzrj2qNSiUE29RcrInJn6OEy46g29vOzz9RCFUzyuQb7p
EA0w7PVKSGzjkALKPFAQmbbzG+Hqgcjfha5dvVpCT18lQX97YNlIyrXahjicWL0qwh72l/X1fhtl
x1jwvHvPVNHm2TsupyI/Nl/TXGNoL1zEt4+izF/iHgbqd44u4kBPQDXWu+HidfEAZVW7m4vYSfWK
JBBmif+Io/lYlGxj5nKJk2gqkpECRRfX3GyD3Vti/XdrxjN/RZAj6cjPO0AmB8BhSn4JqPdMBbEe
Rp0wOYrskpRPIkUG9ekfYb0mOzSPFtRiAsW2oQ9q7kbEkLTVzB01KNE4ROGFkE0/bPGT/UlYejfq
kRXLouUP4i37fQz3CJia92QTSOHcdSUKMh3LtEACZbG0QzwB9fuMyE2tVv4Jf9SgkgUBlTwHwVma
4ceNKzK4BBNd6szET/i7EvPr8QoS0XEaoZA/y7QRWeJE6rW3CT9fIWfyeiE/kNGTTInEZmzDaVft
ocBGjMYCsMcaM3V0oURapTXuRuFFCYQJs7xnwC4fglemcr0UZ1qzLyWWubN2jUwyiqMWTfavB5Fw
PemMQlNGZmhmKtfPfvN3h6jU4FKB/P4Au5BXFPpZ49eRId8LJl8X4tTt8+AT5t7S5fN5tf+pq2yq
2wRfL/FT3iuBDeWUCpk7TiUqeXDsLTt215od4jUyLiv4+bYkWkAYDO2/WFX5kgxiTd0/ssLfM3dz
WSwOhnBCZSBcScLQjIXoCDn6naJ65dMw62C80a6t+YyZrvsrPVM6Du9qKGuvnF7YSQw0JYTX3Qrd
pHwXCB0nzXRQClbLvjAg9AE8MfPHjhkPNMrKe96zWATwZlRm0/LNYbXofVLXwJAdqvAWvXiCLyTT
5Zm2hJUCD5Uf5uN8grRBhaMeIFvkoxZlS7pW8YUQEh6NJydRe3VURDYEGkVGUWzQ7Bu7geRa1WFR
jOLs487SpSCJCffYBn629tgAwlTbrOletBGnYtZukH3nbz9SkoSiPy4foiKJKAOopvHJbfYZ6w92
/2dDv5yOsTqJByBkOTfsN/lmCXbtk/2iRNdWUatS94hgr3elzft980Gqg6G5KjLRO2rPprZDEcIM
gRMXMaP3DQegHKsxZBFjd61zpJlAbiaYc93Ja9a2qIqZRzabPePpyIj2zfxJtXuFpaILZOzsQmWs
Xif3ViVO9R/VMFFZ3dHqxOD6aIljNZtxYo+EgV83ofnH8+73ftkcRpSnf+V7eOsa5mWV86JwZ6rf
dyqYbWRi07S7jatFtR3BPkTd+QKP6+to1SrIao/ue+xBnLrfZSZQzNXfYvSC6pU+vwfba3UaR0Sm
6iUHd69PzhCCpu/ntFly/2jzDELABKiXV/CEqXZZIyzOeIHLwcJKHFjuV5wvC9hDa8IdDUeQOtin
2vlrAir+29HtDR1Dmi1usq91J4ITUPXm8+w/7MoZXjK57bIhCDVklAiquuFmzkgr2lZLkK0pTWcy
U5r/lWn4dRC7z5Lrfgoyvh06x4jOeXd6xFymhUQKHI13nYAYL06l/q83FX0o9qrBBHgipGFQ9Zm5
Q8Q6q+cjZBYHv+ke2LX0B6D3XcJWsuWxolcMBu1EkHVY4dwH/nfBLvH7kFpevr1qTq4IQCpqaJUi
0ALEG2HYCHFqJqgolKJDHHr5RyUvxq+iZ9HD3Cvk1Q3y51H7khTZDuWEQbND/Clt9NixJa+cXWxJ
nPds984NYdEmGvoZI5n/SiJeVNTOvAaZwmpFjdcH6yeUUySh9BWJMhv0GEpnC8FwsDsjUSXUktt5
GelTyU6DTTsxSvTxZtT3TtSiwIBt+lK4Y8s6SLclMTqqJfqBVu81T33ct9etApexh2vYp5SOZkTE
qc8So3NZAvosqgCmqFARz8+2KEx9Qv95VCGiuth0xnGqv/oi4EZvVt3Ra9M8MjBQDFGlmRKY6UzY
jgg8UgRT25SwikO1OVd4EDXWfKQ2b23QYaojx223xviz2gTjAQTc0lVMVexjDPlbTPJL95Hmwa2p
XrUfVZRbLJlsU2NoSbDmw0fU5Vq8xln59WUYA6Z0mnX0lPiRksJReg1zwNyODhfkoidEMo/qW3NB
13kUR7VNG/4WU/8LYTNhiznJhoCYpSxiEn41SH+sqiJp2T/6hlRBrji8rfg1n1NAwtTyeZQy87sz
mRer/8q7ycGMhVs+zcGQPYCGIlGMYeiJCWgNjjANmKZx+OAKdqxPxxBXGHI+njqifs7zG0dTXyIE
Fr2m2YI3Rb5FsIQmMrUl03Tft+mXFGbgeitcytF5kqjUhvhE3c9vPlk1cfVs4xZ8ozmd9BKDVbSe
p2PtjBAKITqJk1B2AD58ijKSyuskgJNzqcI8UrFNjDmfTBGx07h1nk9LcJdItt44zuyvdDgA9ys3
AmmOoXaxybKvjSQibUcY0UV9IJH/LgwIsPdWDg+nhIUt9gBUAUKE06gvHZsNH0V4+lQ8Ie4PyzQ+
llQX1RaUuEPMCDNIopPOwGmgPyOTZyZl0UQqWvfHmwcktxmSwD3vfwqk0J+9KZq0t93SsfyIpWKu
j85JQOPVpzYjMoJgxyCrT3wc7rPHP9N81ICMsKSMFGG+i+DohfARy9CnNKZ48fr26V6mbYASWU/4
fewRrja2N+Fv7+lqlB14sjFnuO/LJGkbWKnuWRTqMGgdn3kSV6+8vDEt4FKL85wj0j+Bfm1JkveA
KnCFlKSG+gq2tDXW+VAabITkwgkQgKtXNpku5lr6GEu0/g/QkMT6N8dcXTnuum3GHYOScu9eg7s/
LRw/gGtnB46ROrD+8nYYVbZPJfULpM5wrFTQaUek+BwcbHmCaYknDkQLsbf6xY+P6cjmc7S0fDio
0PjZtUbGBJ6++YPxxryuLdkQeOhfrcsUICZa3Y7dAltE3G/G0FFjZf8Na9H793m0TeHK3lExmMtu
3qa+j5DoHi8uDqb/aciqOHFkZT/XXFsSF0Rz5fYw4JRndmmcJN7JoDqSQUW7GE1luXb7lYk/7Fe5
shmtJS99CmQiqKoe3K4Dn6KFulN32VtBxuOK/4pV91JKFUAJq7T2ySDv7oF6Y7aV4ryMAJvEU4Rq
zqhMeJLEGjonv5/xVJsVhmZeG4YHqP75IGPSQnIfc4U3HkZvzJV5OnGIvDi6s+3FIJTCXZRCnoTn
WhFGrc2GIQKlseI2PwCcVM0lOuOgW8pyLBwjiV+VN9HED4RtOqC1zMlaOl4zdbAMyIZf4l8a9O3y
qrld7inO6sIBebOjR49HICVchJCMBm1QAX7YGeTbHtYqpev8FAwY7zvsA8njhpHDqL6jvSPDK18p
t1j/XItjSgZcpznzr5GzoudHjkcM99Zz7pXOit5zjF1IFmRz2xB+l0+i+G8kh9+Fnvufi4M6lbLV
4rDZ4XMwEKn0ZWIMY0j9py+EnNhQFq9Y5rg8FfT9ooKAIYuUuYjsz9JmXZS8RKhxQIH5F2YNfeqY
yYbkNDsgixSJEuxN3ZGQvasOaW418dIDZE9WcLsH8XDjDhFMCGdyNyf+8GZaIU6Ll9YhThSZtW0z
wXNMBjDELANXD8Jwdl6sv4f5b5StnDcObuPBVjOOozqy2KYebrXoRaiaK8SM87DWxoxzenKBb15l
lFAS86TAlD9UPtKjvOZKssCPrX8ZRSdiG54Kcx2JNgGcBnOvI90ZuMWj+tqLVmigW025HhJsLbrS
GORM5FDdxwtIFFX9iDHGK4vHuIVltijP4Ib4gQMA4GV94SLoPiqxVABI8/rP1L+1HG5roVeiw+T7
aKsALZEdictKp/DBoGaFDGXzjp72r4OcYiw2c54WDwWuhHqlpr/a4deBGskcHxf/YMFUBOuDunfc
KJ3VwWQCJHli9o0VcdbMasYlIkXnd4n7v9us5x6P0fVbVo0snyovzKze6CqzC86MCV4gLZjKqdve
K48tlKY8QB0G9115lqdm6xIuuz9zrun4g2a2xwuy39O5UCIrdfYGQgO/rA33W3J7bxalDus3OZI9
34ZiNFX8KPsM4IUF3+6TRWwn9/7kD7rB6j4TC40sYbcstbHGmU5Bl+1IeadaCp9oE8NYEi4Y8bJA
75rWTx+9AxWrCULt6n0n9mKYlhLGZhef2kz0+uM6nXheFsUuDrsukr33OYRqpFw89n95xW7eSFOa
Ok/czFgb+KkC2DM5Cq1ataKsEdrnFhX/LEPHbLOtqUV5WYN50ek/U1pvF65MLnnCdZ70Mmm1QuGH
NAxVllkhITPmCSjcjdnAaLIinoxoDTO5/dda7mLZqTQLBI6kyrfI71qtSIjeQQUyebO403JKGj+H
I2FjteSnOiD1rjf6QvsrVetWovBhAyBufdClgNdvJTeIa2vkmam0V20NT5yyBYpmoC5mOKnq+cqC
ksp9x0n6FHUcZj7mn3Lx3U6c+3nap2hqATFpkzDe8XRqZz2kLkJTbbhI+2e3wA0FwX7+K9KlQ8wP
q8hDqjOywyummxNlSEhA9UKCmMxBSN9kPRVY3glb6FG3mmjouOWue3+93AvzgCpSQ07rqGGA/nGA
h0qD6TFc3S+NCrgbIug+GcVQ0C2suzu+rvM8mGLJOM+odJLzGFRzAXN0JvoqtiyyRbWneB24YAZ/
rg2IQObBOBxFwNKY4mpfQSZvm4Vvph24YVEA9F7h+ZzKtHPMqb1wB6Yvm+AbRnvv8PgGMf7dVqPV
Ly/lBDc0EmJQ27ZQ95/AQNwqnnLeiHuIuY5OeT7HgLAwXCwI2q/HHfc6aEKYudcZ2TZP5Ic1ggs+
Hry2VpjjtlgE++sceVFOG/P4RdXXtt1VtZbq8eOnR40oCvpuZoe6I3qvqSUoPEw4rLCi4ElYJYCo
EdAKHDoYRFh3apWCCuQFISbUhm+nEZ1G5RYZoxRukTtWp3bpEmyOZ3e+8TUYaAyJMbr+PfxLlBSB
1ZxGOwHY7NkWU42GO9aiB1+rApp4iZhewjhyrlCsdCLdWspG/cIRjQPm1vJ5aNxKz3uG01Q7szbs
c5ulgNRIis0xTNuHm+MfDqt77cc5YKk0vZQCnX77VcJCFaeN7evyOpL8DZc3xuxiPcsZzmIXdNHP
TTZ3dCTwtwrluB5x9QACXpqjB6Q0Fl/Me+u4C7iH6aIXgkljbH639BAtE09uBbDlseA2Bvc3ZK8X
Wy9pTCVgFBG8tIRY5dyNLcqzWc8BGfLwS3/OyVJcBhBzmVqIKmyZwXN3JFsFhJU5UxyLZ4YsXMIm
9YHm8tNTE6V8WKC6XStLWGl3AGD73uTelNegxfun2pgQqoFnORI6puS34npQPeCpAvwv2vUOVFBQ
So3y/myuAd4H38JA5fmch4ZRD8rsxio5w3bmmq5cqNjuEBtylyVQ5kFcwXIArPCJ4fyJ49JJIaUQ
CGKWmaPu/eZGCfBnUJM2cpHunKgdfuJ69b/0xlCr1of5VgnigrLxHGwSBAi6mdzkZsp5IKnTlOqz
rxmydT2m1L94b8onJ49Kuje1dibHUVzpOXodIEF53/n6RLylZQJpweyWKMbF38LH8UNd0NTnaZiG
/7JXr0Vqe7r92zmDW3m7IRkmDb/fVPp3YM/aQ6YHklHUHGl/PweGCZHhkexZ9iR6g7ZKi8egVXbu
M3DRULvRLaKgZeFcXcM/jUnJULRlWIa6f+T0evletzy3/l4IBcPL4Hpt57u/vHLx/1J4KQ+oioXG
Iry7YWtGP1QU+hRsX52fg5PVSOOAqtRbJgmDNrhV74bOBMyhDy+GD+2lWBArWKppJ/dO04uXBjkn
Y/+yRiDxcPEh6PTmv+988jovJDpjpdJhKr6sf38LuV6nW3fk7m1SO94cctjIu1PvAdJv0IXtuwej
NYNdwbrK+l6ilaDdSD0uYfty9YVRxBROIeSPZTi+jfoihYyi1UoZlT2QTzlBqp8nRBoAUQYgQnYs
tXJ7o6e9w59rhF9ILBAa0KL9rHqhVySnKtL7uKwb3bxB8RLr/L2/AGM2Fd4+HiOwBCxCxBO6hW/U
7M+RLb/Av2epuYAI+x36nJlji+pyoFVw+sYA5/ynM3Hnlrq2qthNA6DOWfAbBHdz8ELZqlttfGVB
VxVVoaLRgzMuRPgqgdWA1UIDrf4RlyooZWTbspB8sQ++ocN9Y+R/wXmfeiCjI/FRbiQ4aJF6cCvG
M1Wlp32lc9zmJjYTMWFHrERn+wYf6oQ+oH/zHWjkvD6a5BiBxscO80uWE6OkYTs6+t9GUuIjtYP0
xTEzJdIuRAKRKFdiayu98W3kswr2CYlvS2916HG1MQgSkJcLtD1lVvRaBqe8SFAWeKU/5rNTTN7v
I90Lbpo0JpP3nlmoUHS8OdsnYa8gs9/xF61s5/2CTwfSusTpsdLBPUof2JwewOQn2qWx+NvFZf1A
RZ6DmBGFR09Wu5FXvMvhqkfk2LSW8cr7g+oPZlswrz5cv5j6jFOst8NOBNYkK7GnUrr7Vy6ZD6ZM
pBnhoDuiRWeVP61CFq6zxMu25pYoYUXcLsSr+u6A3GUXbjh9/eqTr5qaU71WQq8UDBykcvsyNww4
WOZgZ17IFmD83peoxP8r3bNIdpmvzvfqq5SmwEogeSWAIyK3sdwMoaz4UF85kjOjYq6+DWMdnTyO
RCBW7AJmojSQwqQI21/q3VgtCsITZhpIvjkR9nLfSPgK44drKnqWC1MosKerUh/kt3r4yu+bN56j
Mk4c+ybz6JO0kT4vEudkNeqO5Elsg7firgta3ETlj+EJMbJ5vNVKBUIEFqLFdjM7oBGOc/giIVBl
/ZCG84Lr+GzFgj/zIXgL2vcJ/QiAMxYDaOwgJPF7V5OYpAV9ddF1yNv3xU/9O4dU6Wf02qjRJAr/
0WOj8XH2vAjYgSt8ZaD6gW15F+bv2qt9id4TA/7G6QwEmaJDi1CD0JPdAgEIa9hUcUZaciTBnqVJ
LHztz1Hs+ysgccWLR0n+Kgvt1/JtfJVr3qTBqq/F68SPRF6nvI3FBi7jXqWm/OC256uMfX5OANud
Ucx5xUJi66f3qhpcjy25ujdzqbtxZqOr6JFpQKZMX6P8jKUJ/8yX83FG65VND7/QK2jblwynAV0b
1Xcx/FTZVYxWxUOFQusJpHUGg/HYvWViIy6Fs68TzILCj9+fWUhBVTSpPTkE/RmM0PyzAaUIimY+
AsRYNaDWw7MQ+taJei5AXkIjuvI+EFpqJCV28tlWzKa797FG5PgGXWR9oA9QpfDub8IfghcrQ6RY
fLA7oAUwlPfZjemOn02kXU/5W9M8BsyXCcczu/axJS8Cil5BP71Ct+8qX/OeWuDDSJuDHKi1oUnY
d8FULJS2LdgN1xqeOD8ahV3XhDs5TVEV8u8laHxrUxAuC92LmY1iMy7gciRA4xZNGBRsC1T0OqfM
joxT7GaA/u+itbfhj2aFv5dFk6OucnmybJg9Bf2k31kulevlxr56wRLaiA8fbgLENfv5QnozF+UF
2bk69kcgn3QOsBKfk5BvAKHTA+G5WWA1UP07U7lGDFRzF0Uk6EwvZmHDQ5KMGyyjZJdHthjuwvlc
jk+R3deOiZeDjv/BAa5AgX0AwhcuP3VD3crwCCBgmCwyKHwLgn2W+e8M2fUykK5LTiN+DG4btsaW
oHz89d3QYJMQUH7f2OzFepu/YYuVXpM0wP2PSiq6Lse97K5gnMxw1lopeZsLrnXP/qJ8LEMosmLS
y4AmOaO6R73RVGHiI6AE3dCrC75pXS8e1s2hzHu/9j4PALiswrbYjrbS5sV4pz76YkRoq+PUip63
Iw8j3Aj7mAPZgl4hjq2F8rBk46qAvg5bzWhUhANehSzcZIpG7/mH0di09MfhOQh3qguBmWK+Zh7F
aCXdbDi3w9N+iLauPkngR+orK44y3ARiRmoTmxJURCUY3ogH+C8cGt3TId1iFZHjIGdapB9fER5w
sef8eLVhmtuD0Vw6/bosoH0Hg5DmNe2pVis2iNk7opaLG83yVDc3KdSFFFKBgUcvHogB9+/lg0Xf
jPJbIs83LUlB/RezYMom3sSjFoDlWvN+I9aodGRMxQJEIH6OgA5OEmjZOZBf3c5bXFD2z5QVO7+s
h1hMEhW4NR+1KEJXdpm0AP2arP8Me2MjJ3wSewgk9nWV4YRsgD4C8ksRVumMI+ErKTJ2RXeTPaiN
kKjfYMs7FjSdnMofSQQ7WRQxg0q9ATHpug1Yp2w9KHPqlFeFkBUrp3k2Z8QlKDwEdFo0oGV32u4w
x+SDjTjOT/PdNuRZqCOzHVL3rtHFiMTScU5391rJ9pTM3i6NwuZSKP+PJdIM8afFwoaEvQFF1/4u
orHu5mwRctS4jYBOKbNNyxz8xwom4RtzfAmooLZ5cS78xbh44BZ20/YPfx1vkfyyrSEMexWUuQuf
jHa/VmwwMTR79TS3wT8oXw/Y6JT+cZsze1czfpuSj2jh/hHSyxEuLyk5HwAXwHz1a5RlhoZWyccH
1Xe8Tg442NryVGieMY9sIXw+nJW58iVaZzAOtEmCmz244TsyS0YfJE9Q4FmR678v3ndQRc2MjCd2
qTSYwEL6F2nr7gMCWwSlewk1H3azJMf83FNb5i5vLcKvuUsXuU2k4+S8sftVSC1AAp7SGAFgBpZn
v9gnM+U3OTAJiNrbhIIBXt6imJsLjh2uROJukjHY4hqLIA7oeaD/wV8vxItwXCH5/Nc7tM5Ek3wG
GMyZaD9rITwj0MSNbPfSr0vUWIQz904N/sXRZW9f6R70SN7uSfCelUFGfxyertfG0TTlFIvHBqVC
8e4jnY7wm0wV8h2o/EcwymhyHUDfTF9H/ydw5acsJMm/pUJVnVByfv1OE9lU7yeOx+AT4M4mBAvc
/Hc3NbYrukMryebatg0oMwAdebomlzDi0oLVZfT2lukWQ6+I5k/LsVgH/gpRm1QVayXAmjDKUO0v
Dx8SBFTxRjcN43DsFjDqHpA8JWWLVDsQKpz/vvUGXI0xBiLqGVlhPm74JXP1OjdwlzA1wnuE1IS8
vp5UoGKMrc7nYrhUfIpUNbDQKvqi0wb/J0KdxlPBilGNvkyUnw4RRBYV/bNLjesmpm9ZKHI1ulE3
MVId3feTcgRE9RCFIzuZ1V57rCcXM9gkzq0eU/pcMnorTWE1eBnyPzmr/e/99Y2ntR1nn1suWifF
KLioFjWtn2eFzCSJ6UgzlLnjtKQdNkviYa8GJYR0MG7K5khnTnMPeCzn4mjDHL/qjJKDnWqXI4qJ
l6bHM6Bn8M/Ybyqraq5gVG8QxXmGTc6kgsuTzXxApxuByfCm9oS71Tyvl5bm/++5UsvdK9Dj4Q52
vl4TC1Kabb1h6++rDgkRhTpCa837dP4A08H0hhwN5y8zsrxWkKiroYOkmqEhoUwvBHuDj7NdGrPs
7M5M3yQOnkMyBylbnbUeBq2Bh7k1/dcOXXGiWbYGuIrI96xjFkk8YIWHM4tHpXrZYTxjiLnxuUW8
ou0+Ip7844NYqHtdugrfPtozflUSw2xA/oTxZAhgw72WACwjW10eMyt1PEb0u05/PzLnvVqeFMyc
PAPirFGhERdVsmMRqR77eT38jSVJff3U+Zq8Y8ta2fE7V+UXZBFlB9FjdrQZ68Qo8KtvGqJ9X38h
Q+58NPoEmF6n1+lb1J72tk3XnPTO3/dJ3Y/aStp5bZ0HaUfXuN//ADx73iDgx9j63FuOsq9ts7iz
ZKPjufnYNHAHkIiqMxXHl6FhTy8g29UpyWapvrHVEgwfqqXkZJyShJnhXefXOC7aoK+yCnONM65u
9+JyHpzteCopTTDIim+KcNOIWMMwBJ05ktwwNo8dqtO4g7qGwL8GTov/zcmH51JQnQH2AUM1iD0B
2QXl8ymUGH185z/9yjHVW+oA4A6bDZxReG0inMRSqm9QikimffBzswjJpk7BaRXcW9sdHh6LfSDJ
scM+Lst/U9ALm1B7ZlKNuwMvlqlaQ/5COJq8HO0EgZJRHS7cSb6kPwQEWJkD3/7ZafMQhuhlwgmo
8RmQpZfPf0ciIYgzg3/VPFSILnUp7tfmT0hs2ojw+US6At3ZCfy+32vAYAzBZL7p/l7yzR3nHSNP
lSJTXeouZBQh+RaWLEjhWD/a2jTHVIsv2UaN2/xoqVGdLtdN8E+UsM6OmvhVu+v2Pp788hX8DJq+
2OaNgMO1NI3d8u3/X9bTStAvOqtvyZ2BFdrce7Ko7MparMZfGzaGl1/QVDqmJ1mpj2KckTMd3Lq9
Hr+WLUP8tI0h4TPVswFmpsUkGr7uA8yWyhEgN4lygpux3V7vM6QHvStD6xAfQLoHEYTaID+lT65M
oEvHGWG7FjrPequ+MepA3oBrHltPjz+uDjm5NGY/igOJiCeW9ErUBAf4QKCh5Ed7C+ZaG9/mmODp
k9OisyLpiPjz0KsYKefQ+qtdwxm2/2Blu/Ch0MBM994G3QMQ+NX5Tex/ecETPMMHr8qUqqYhk6ME
44ATTPI0dt5+u6qqhIwmY/BSnSVEwCWsLQumL1DGsnNmMGf0izJTvslySrgXaTF+nnpjXT6+7MvD
bm9vLPFJLqvkSeNlx2coK6eGh4aJFUjCKmN2N77pgUhixOcVM03zGBT/TnvpMRpz2TlOAyjwa6JX
N5MiyderdpghRBKbd25pEKukU6jRBDERcCmRpVQWb1bixz1HAS+MvHKcrk39EW4kPKrIbNop1nb8
JU8Jq2GKgK5GOXjkhx5TOass3fVm6VOeOX1gpCsoq+oYgVVwNtV+/58Mm9EV+y4cfVSADKwjHegn
kXPLWD2JH7FPP6mW5QtRERzxHbNqYJ6hUpuXQQZ29TXEtMbgZcQsRyfd2Se0k20LDrR/muJdw1R0
94VUW6wLa5c0goxN8oj5R8gkO8z0WLK5OxYg9MVUKBK+H8gczrS1NNyc+nKzD2laNh4WZcuKqE1p
aitmtGF2wd2c2U+4op68PqtjlorJzk4+NMWXaoujirpO5zA/+SFtLR2lwZlnLqFlqxlL9c+dMQZu
J328am8nkaLFJmJcitPiqm3/IKBy02hr9n+Bev0pRFrEB0vfUKK5WYTEzugnqIxZhBrCYa0PhTfG
8wo3K/stk1vIjQV6mpsv1v+Uo3hLj6DM1neay09tH+0Rx4yLlHIWxd82qFJb6HPbzM/tUir+vbhh
5orGpZYwbrK7Kf2k7ntzdA6ZtO+78UQi3rsYEYgibtcjo/03MowcUiz314mBAg7PCmlS/wQsZyKj
iYPu46ERN4q12jaXwJLdSseurOmub90KgoMLn69p2AIEnxim0GpqFBwSiYmyMB/x+TmzCjR88/hg
HXSo6OLJK3p5UAV6YQTd8kXd5wHas1xhpCcQuJEb4gHqXWrt+RgCBwldWC4I87zwYCInAA+JQX2x
3M9GzMq7Xg6hZjYzxVWnEBIrftYm0VSkLUNE8xkjiZthP5n3wX4ZFBrvrhVv1mhmFt6bNF+KbGN6
qup50fvF1oEj/foXgH4P2QywPxXP2Y369O0mq0c6noTTKLOdPibPuXKL6ndR7+7YBnON1tVYYt7T
3nACuzt1poQxjVdjQSAYJqRTYuzfUVXxK28mzzYVe5auB/YsqOmDr5PIZCA3Ky74vC52Y7eMxuWv
Gn/tyzwplhdoasqdJUvpzoWMS8oLy2LsAsh8TNBsidQZknsFs+MbvjxtXx38eNWKw2DEVrATbW3u
AOH8uY0BYAmAT6hN2GOz/gWB9W/sAUJoMMLGmNi+06yiLtTrip5qjDk23KYmArXlt6MZzjx2sBc1
mRqdu92BK9i0M5x5x/dwEfpfEf6DJ8uOcgmt8/ix5B5SeJF5VuCG7zB/6M3dWVf/SUSo+FTUqWkm
ijPe3y3ydX+HagvVlmTnd4zLaiZont/biIVuwvO3xW1UemU5xCGdIm9B3AL5plqk1X7Lx1h8BXmg
IYFpGqBI70gXDzxgdauEamQYvx9nUN8UBXmWuR1EOlpZbY7A2Md7uMallQwkRafngxrkx1l6bIsE
odZCSWG2Fy7nW4IICZp0gATh+GT7xB1vBKswn9kT7GsbLquZN9EXUMAvmeN3OWJrQK271Md6MhYB
pW2jERqtHnrONtDrnVZ1ZKfkA+fRPsjZTR+jJd1VgxvEImWuIY5lBnCZ1pZKinLv3ivmYp3XlpmO
wJr0J7KL49rFRLdhnE/itl5FMl+TKnrF8Cm1CISct1UPrd8tRPpHsR26mVzapx26izeDLREn8POD
dTvxHg0f8qKUDpXBvmQDB3LoVbqwO5j0/oyoSFE+rUskxAjirNSWGqFH2f88SmdhAbg6dTegm/Ge
vSmqAa+n30DFGzROQvn6onWCrEus80VyQ6dli5EFKlwR++oYdcuXToLM9mMLgtMVzytR+nsR37pA
gfCxJEINfFggCmzwW2PlnBexVLSQX52wz8spw9D4YfWAoO0hiHkIo2CFpALUjBInw41oHIH8y4CQ
Hp5IBO6Uz6xgwo4M+bGj2ug9x9teTGFmx/zScyek2YXvTJgQweWltX74TjJiQ6vBC6Q7AwkH6Y0N
5Td9M/qjWMDOL4ZQbSFkkMm2aoMuX0iiHsY9xxpqCOBPeec5QPgf79b9S5irmIq8MtxshNeR+8Fv
YUoAAQ3OwoZwxFTfi9R/uLiJ36gXmrF3xDIGQobl+OtjSUD2DoVvpfwRHBoXYX8WEy/LcT7rhbJe
MP1pUDUnGrtDCwjUgTg68Yuy3NPxXObIIX2mXZ7VQMPidvX4u5k43HsRMu1IvFEJNZ0nBSnWsMrn
n4lCyM0atPFqTTvJ4WL87Jh7XYublL/U4gZxRE6gQePQHR9UUoQ1IaGNDXVbG2ZLxBnrXWEMid11
8xY04dVQqfRzidx9nLuZgtX56qnILUTHDEGzuCAaJ6bkcjdEjmzWeQLa+9QUk3GjPQOtGTZ0YSWP
vFr0bLGPArFxxTNYMeTIFvsezx95WVnIZL/9nMqgGPrO+TQehi/DAIG3oldQqoCajExbJxeapZ29
M3PH2sMkR27SSxSJlcjD9zR+SfSQXqwTGBxgmBK+7+y9DBmm2ZZshPhSX/ucLanOHxIOVk4fL55Q
wiPlfcWlqFYPe3RqEBG6Cj/rbk00l+BI+0h5w/gw1mkdakb65LFwnHBgT3H3OvK+rBE5ZmKmywif
RSFUqUEFJtUR18f5xC3YXr8qI+zCOSUYjNr6jS39bpjf//iwMm/u2nG2ubRQwDRVZxod3T28ha/A
QK647FBAoDBGcdyBc49GR3mLnX1/pWjcNEF1QcNTl+j3zkxWkl4e5aJmpkH8LV4sYp9ZRIiixWW+
v/iA1CVwItSC2/RZFrmS4mekf8sSpDvzE2hbcOj/3ZzwTzyb8nQ5vnhCfee63rQRWPffvriu5NQe
FUHOETRupwMV+8pGIzZW7I9Pt05t+eamUL6lb9VwWtojZ7B4DGaV6twUA41fCZ+xAqqbE+ilH7zG
I0KZheMm4+D+oXwMkdm8GSfcS/fxJoeUuL+K+AysIaSXCL1/7DXWM3kDMPpSHsmKWWlNzRSRYD1E
2z8/bBnjCJkEdFelLegQMW1gIiwkGOwAUszd+Kq/K7WALCfvC19Kj/7QC1F7au/HD2dy1+hy3XDQ
qXB4qz8DZU5ovRD5XFoqnrsJnAcTEhFJynLtEfB9WZ7nA78UHcan/C9YKxjDlp3YkoQEn8c9tR2s
drfxjlbidW9ahknYp6R1JUR796Fh1rdm11toT/MuKXsSuH5mZw/g5m93wKC1Kq1vHvotdVLb0dSL
zuRhvznsD/IeE93M5XmU2NOVVy4iXVIMmBpwJGCg9/9o+7Fs5oCtBlHEtw3CMjGM5kSDlga60czz
1loQreQEpLhtEBstyR6YqwmaTf6lCvnGdfQTf5SQ24DeMTnND5nf3C+983166psT4i46QvzG8guo
+Vwzp3SEbmUfB3Fi2uHcKDCEGFCKCBbCOzZdNs1SYTdumiJ0eOZsd37NG3bt7424NqrWR3KqaUwc
ldqqY6kiBkzDs6dwZpYhPuCLGuX5vdFXhaHH5QDioz5S9PWwfehoQhv/l5Y4K0eBHwRFBDsUEkP2
AiC+BgRY87IWfJqD/JGCp4UUZV1RLOPGe9O1VRH/SJdffLQhtsX5lwBWLr5cg9yDUEIVInX4E9is
/wQUu5HenJTP4BqcjRuhCzNb75WN3hogdgMjLjCeBpcxjiOXXCq4ICneOF9TLscD23mywqs/LrWr
+BS+GmooN5L2c9lGNylWrBgdbiKPUdLsBxIpzCKZyVX4fJqQR1q4RYCStp3Z9H5+Im277A3C6dIz
AT0WNEsIveDRwEkyCUsAKlbZ2aCGWUzRIZN+kvXdCGmo+aKS4v9OGs4dU0e5t4Ic/j4ci5ScM7F9
fDxO0WC1FRrcO7bhznjsOGbA0a8jaOMEYdoQQN0kCZFgbcLtNLFAtm3T/IaA50Wc+2EcxGPiVapw
2mJMgaAPcVKPsw1MaRkQPjK8Oe6UNoz2fnQdnipNjx7c8O02HtYLijTaPRgIYHfQ5uQwy1sGZ2XU
Xtzh7nqGWQhWhM7WC4bWo84x3hCdZlbvXC6VMGCYYUdYo7c87F+Mg+VcoEQFdvu3KpSzxT7okESD
LmddYU09TOUe10oZL2Ch9/lCkl2EVFfI+8cb4JWz/m3kbk9QVxTo2n8Gv+svAM1hasUJ8f7Kj/xT
hdVD4wT7HE/9yuMAZ68mUoiuLO7Kk+uKuFGwGBJSY9Q5kum7eLvVyzLXahZarzK4TM+uXUW3E3sx
TpVtwYyd1X8OXcggDKEIM1S8/5zWX9Bjlhbx0pbLPso2ODHXod1ydxtR3iEyfBGMHlwAiSYtNsD1
51nyiy7Gl7yewSfulUWZ0ZzN6GS4BWdBy0PmKGmedKzRzALulkVuJNBJey3RLFOysPhhum7xAwoG
ECmpkhanIr8P107JjqAGkj6QcFNjCq4wJgCMdmfl5Dyxux0nQZSBn+I931nqKyLEws3O4JNDD8iX
EuFdLkKoXxmWgFaqOsd+FGCG5yMCHFT7pOj/sH/wZ/s0+gYOJKAklX5xdVkFOZSXZPFxkMZXX1CM
DCbNtztv7m2oTFK/0thX2RORfPi71dZD9AuU4Koi7KtdtV9bCoSv5pKorHo0FTx//jNVmuOYptoz
+xTNY7xB5La6oh0avAUOkllw5gL/h4UZfa9UPjN8v1poq5WzLOKSoH8CuLEL0wikAYkjw+8WayHu
9YDdLvhNEXUiBej5jD9IqHL3f4eJRnRYJnZJv81SSp2KhjK7u/vZz1A5nR6B45w/GwtOVQD+I274
uXcNjRFeePIlkEWZNZ6AxCBCYbCLoLeapJY/zFGMxNhketloCrgwvpz0PG3/+JggPY9FHDTN6j/K
OZuLoieAJ9i0qSaAwGfUiWN+R5GmfzGIA/+mPutEbUbQ/yA0gP0BBlThVREvzlFVivfmD+VhA74n
57KdCN4oRdtKnynnFGyK9SafTXnsJDI3GbZ/TnqTpDgMOkooD92JtXPuqYbgqeMdJcOKWdFjVy0d
CN5pBHLc0Eyuzewqt5NpNStKqepFzhY9OKeank5yHKpdwR2KVQMf/Bzp3HxcsL17oWECVdjXk8Ce
WanuhNeiXm824lQORDwy83RPEE75CMGmPWxmTL7JzIXCBqEGOH3QIprXNijm5rueVTngPa9mirym
LLqcxVQtLe3fJknln1WrL6xYnkigJ6grxDZSH7Yl9lrmsq9qKwGR3IkVT2P4LF0j6GJ+mHERtohv
H4FF9BCV7pMinewc27XJGyO94VuIsmGThHKalbLMhJ9m6OxSvVRWix5jqgMD8U3JAFhUdLz7lMbx
6vTrrTS/4dFKDi5qSXv4R8TYQ/i4hqFPRo9h+oC1zk2fTOvbgIxdziqYAyWRoEt7z5H3orHkBmgN
k+UkPemfLtffHsxgdIStpX3lB2V9kCa4SnOoEoonSh5IXLyXDl1oEBMGAa7eK1vaT4KCRLjnVTrY
ci51KzaHQPLym3U5a6NxFmIahC/SWbzMJLskPf8VDyUlCv+ruk22WUCBquthj9Pxlee8BQ5Y/Aig
wjsuCQhEjWNx/vnE6MHxow2HKBVHpcb8+5MtVTOZEkUubRxh+HMXGxjRYHvbYqwueIHzfR5zcm7Q
vPvrJAcF5y+XV9FS8267VfqSofElShA2V7at5EFzmI7jU3iV2vyRObIXR2fhuYUMha4hUGiniJKP
dgeND8c4Mrg9MFcSA0rYBV52AJkWOkZORmckvivTspol/1anxz3mBU09NiyXeeNE80qScssEvVdX
XxNH1H7Ow73Iw2H75ZYoI/KPu46AB8S0K2zy6FYV55nFQD78gJzr8DAwXvKwYNfa+kqxFgRGL2Hu
KuW8ILuQHKk6RZ+YE/RVm6nxO1rI30klespBqnuzwMOtc9ZLWqqBU31c4Qe45r0VtUuuk8RqM1xM
xOexHLGE8uYZa3ibb1XXcAKdXvVV3IwiHv/7wwkLzaxY1V/oF2Xdakvlp++bPjcNl8N2R+HciM+c
/XIA+b1x8tQ2GyGLQX0p+2QPJmITHt0WkdQV1vQB4Efl/Nqy/fcH2yg8tckq1d2cy5BHFainGCXj
OOGdAfhnr60vZQYdSkPNmDkGZeSCDRm3enONke2X9sIxKK2zpySLgx51EdKaoLdb4OtA0BVXxifI
OJEPGTTsCbuXgafot5SeEt4+uvGzNIhmBf+BxeONCPeX7xpEdLNYJTAzOAiSXe9gz7PMV6AXRCjd
/M4RG/EjIcOcFkMdihP0mgprca2LLXwoXvALqh7ezgUSPOyNOd8yUwn6hKdyGK+17RUOxh48+R5D
yPTI1uVq7WaBSl/IFz3RhwcDbmAxK0G2pSEIi1zLp0m65LK1uVnjc1OEgD6fWS5CzsFYSYiEWXQx
6s1c8dUOsRZJCtpII3ZDThJ1bBMkODpijAO5e04xAeGmkRZQjd+OASE9AAt1irfmZimtmdY5z/zd
rvOqSHxT7O5ud4YsUk1PUZFMqDVgZ1xnW9HOUhXaR8rlmNA21lO1Scppp9mMem+sGMQwdk2FY75R
RFxmgdy6PAGgxwffaw/ovAquxsTPpDiQIa6aPwTVSRUH1AhXChLN3VqLkqhjiaVgnzMVuqR5lpEA
DoIaawuVIMQFW5haGVERzcCLkApcpHnZlWELScAaytKV2+thEWFqJ7ZT4RMuiie1OCuOrYOyly92
uUVMx69M0Z/cc7XoYdTw7bF8ybrE91lHfYQdRMANl9LVlfGyKPv0kHW7VQ2UA+OEs8CjG9EfyiOZ
dVNc5jUJKMe8e7ujWNbu+1zAXOKzWaTqQMb9YxgehXZAdYVCMt809o4zjOaHzZE+1bCwvNvIlteD
tFuDFgnD1cB+FTFo5HiPLmcHRv2cy2JL+8sWVQQPY5HpwoO6pxwumC0hNdgVNsDOBBNggc6FyGeY
ko8YddtqLBRF7tQZw1tAGJsGVGk4jcNswf/hE7Tm+VYb3Z4AvletfO0n6wrVI4kSiZMrr6Lv0SB/
hxoNzI/6Yg1ZaCD+jqNprLavADnaaKE9OkG5UA02QfsLWhJd2dxWRSEDT6KWI98thWDRZ9/R/mL+
eaWSm1xu/3+I1iG99WhkDYRdYjszhE922K91wMcvqZ49+9ZF7AsiV6F+6r/0kCGaMZBLjaup6aVf
AB6C28ZZlXqAYovDAyZvDrp/LM3GEC7LXZmSCw7KFfj6Bae/9sZq49F7gvuViKhOaIUzLC8qoNsH
3SuelAQ9U+pRv8ZMdjPt0ShvgLqTnxq1xNGRyLkMuqxu+SCLfYA0rMtU+TpxmcJK69B0YSBW1qV/
NX33XC1BJu0F/NozMS9PMC7O+IuJpxfHkZYOtutS/MINGANTaFXHOrgqTdxdF8KAPMTcLe21iCtA
sPG27F1p4onCKdUVJRRXQB5qcaZnhaEbIS37q042mKOaysH9zRjWbTwipIDDyNxKuLmsOVOTL4jK
hZUvSjgVEXuzuOKQ/6B9I2hECiM5OCqPU6li0o0bw1kJgyU8qwHc0LzQt8TGE11/gc5DH/yD34i6
hkhvsBL8VQVTYd+082HTeRrFMTOQmWDCU1r3VMJ+GUh1SINEA3zQs8lh600eaVbRZOTPa9hwMKeE
H2Kse71BVQegfmke7fuLRSOTAQVVVk08cGky4rCG+V8CZRQLp9rgPJfqDJsff84TM3T17LlSovHm
q1x/6dV46Sx4+K5zl3fY7yDZa4wCKPvHTwmXFlcrjAON0/M2JTogRLZ7UTxcTG37E60vRGs37oFi
rG0JFMhBD3ZD/M64FjO1EJJBqz+ZLhcvRKO6pOyCVDPwUf3AupyltchXcqmGUAu+LJTQ3b0oGnQd
n8K0u84sEGDw8AJ2WBoLBQCPA1xN7nWDDjXIEueF3zgGc29hRHOkgeczXKnRAJIowLqwZp/6Jlgc
imYBmXqEpXjydKhIW+QSGB1rFG2y8T2B9ZPNBowRE+gXkX5AKz0kkNSL/j7eQI6EiaRluH/Uw2eM
EmOc5FSSxE/ut7bUtJoXw6ks86Vao33sNDPW18Xy72vLNeYG56oxnPlHz+UWmi/tIvu57ULA4XtN
alklDcrdDR6eJBbXbKmWcIKHqt4eXHd9hIwXw05Rj6DOu86uAkp58Avi/vtG7bEaAk1Qm31rLg5D
A5qMCfcobQyvGUwlv6Syf9svoMtFoFhTJ7TaH+bEG4tlhKe8J3WnLBZug9Yobvk4Sf7CynI1mkej
CBt2CsifFAAGwDLRNKTgMGk5OclS/9GDvuw/oiy08CE5388LJmwzR/YZStIT0joNpQ8hur4YveWT
Uw3VPrUP+gke8v8vHsEB4dmQntCQ0fisyUv4XDx40GOtdAiwhX0uxGBDJRSKcjGYbLtvyMdHgx5x
9I7p/awgsQbjN2ECIwNV44XG135CyF7Kpp8sN/5NF7ehb2KID6ZI0YAb7fpXdYSh7lzSmMByxfhG
6gilr5G7tVL/pDb35lX/X9JKSYaB/TJ5jl2rZMXI/XDwxKrJYRuGeLHtDifUYJhKBp5RG6BBHOiS
sH0zaH9HH63HIWHn2ODxivaUfQx9c7xUQ95Cz36RtaNhimEZL8cODHgp5uKsM9dLWIrhbu7RwEqY
JzukeLrFwhuBs9t6sP/BwNo28UL0WlVcgkhHo5vpKhPYcZer589i7+Rwei8Gu18sqiW5BuvuL5KF
pD2SgFOxTr1e80UXgV2LUcGWd1Yd6LaM3ikLlpeUGvmS+e+Ro2fpoKMu/AElypBtqwJtdVsscnJw
2ep/583wbKRuQMA9FZ6iB7lLK67M9rBtdqhgsUSAf84i4tzhISMFc1MxMjsA0y1h4dGvWF5NKHEA
AXMrNbdDhpszawUGN0OMzbDDm8Xnh8PNEG7X0RKem3HgPHmb6rneHQwWawmLhoI/dJtTC3eKff6a
O2vrJ028V4i0eYT7VsOfsitm/3hmJ6UFSYiW+ICHxBwqqeMrEzOaz/V4P+RTBD4wQhWbgWkFi08A
95HcJXJCU4ue/gnpQQzgn3nCk4EU8JLOB0Tr4t2bSQhzXdgESINjDAfJnOKNG4ueB23PB798S6AU
mvMCOm94udM3TyPHKvmaYALgz7w2Pa2L+HTtaQM68ag7wfoxTyzR4UpG91hVNw731BLT2Cjl1fDb
dBwnnzVS3yeB2jmN+1wtM5/lP5ddEUSuHWWumIYR5oySYEF9MaKVNGaDXCG2z5Nhs8EDeobqdMfj
guNKFF/UrvwRiVBSIFO1PcFbkHw5tA9JpBVz1cVaCxyYEqpA2P8cdpi8K/g0ONen7Ud/zwCVDwsu
v32zDDsNXptuvMLABxhp21jiPgRodbYcstTnvDHjq7WFan+iV5N1Yu66FreCvnAdHmaYLiAigczK
W9UkWHIPkfZuz3HpyJZavU6d42DBtxSGPtHtOc+yY8c3eDy+s7FsSpnoNd64sr4gz2fblk02WQqY
18nd9Z7DG7J+VyAdaLp4HeXh3daxig9ns0e6dwTwoTHwOVvLo8rhz0dbKZx7ksGsRe76X3gqLXMc
CuRLQgyTBFAiQ4NaccSlGkDTsos0bnZOLm28HQ1IdRfJcI435a6QDzJEdr5e41g55fbRPm+PKpBN
1D9p1fqcKa9wQ4pa4fAp2dAF46AZKbdHrANudrWb52B1+tIDS4iVLD8ILyx7mpS62ztrgwlWg9/U
ocZEUWEMnDSV9i40USz5aRxB9aKIveIX3fOd8auQzGP46nhlqUDhShwzW6xvhBpxX0S5vEn2aY0I
AB3+cGExv2/A9RTL7EqDYbmtYqUHD+UANGycC+a8DFIt2CSiXUMkS3PwQ1N3j/AGwpdjFf2PxPZD
7YRHKEq5AjA182k8zMXw/RdZIwz0E6DyO6o9sLF4+aUIWgP/L585P9Gt3HZBjw5LLYDYlypD9Ka4
jeCLV64Z/2+f+AyNcorsOYbu/XzxZ0g32E+AG4sgR9IONtBoKuJfZc1JyOJb+OzEGkSznDuYvWbw
+Y5XIdm3G0xBNInV+rQ4dXlOTF3HIAQoR9t/I0uJ/kFwfi0/nFVuSE3qurF2l3atGTPrl3PT5RXs
YFryrlKpZi+vsDAVl8fJJymXWcfq4FxWJWDm09yjCAfWFM/SMZvRZvxIqXIJ/zp2jFI127jXKIiX
Qa6EChAvowWTpwDkEC2tYCSqlhRkBD/uAlj1t84TmxcmNWMlL0YWZSFSAvimgtCvreDqNWNrpdn+
nN9gx8qm5gAVPrdLy0x/ky0mG6HrVO5Boga8HFAgmJg82PVjLaiTR6COC9NOFDCk07U5ItXnAXbn
bpETbOnN1ALLriIyI2DBOSQcuLtsz8HLuA6iyXTP3moFBckwmEP97pwTM6YM1ynl0hpMhiQKkVCC
MbUFiY4XjDve7RjUZZC7NQN7z1HnsrE60Oz15SM4Gn7wiAuMz2uUEVKukaRTQKhiDZUrftwlpgF7
pUIgympO/cPV0G+meqMmj449mDALr9D0tCXP2UtapPFgRHuKw9Gy78ClAA40bcklB4l2iPSG8Mta
RZDz5hQPDPfQWJBbFWVW3ATBvWBbZgKQ0h4Q4q0X4ZzHaZuduE046rsra9WfUfBgD12G2uH4d4GY
Nf+sA0LlZ94Onae0uiK/quXCv1UkKh5CAVFJBBc+JjgCloq26bAbGq8MY2VFhSacK4sEWxUfxq4N
6yPNaYb+hEay0QX6GkjjDQQw1pUX5idwDw8Sv4WbHMritDnT/Qw+eOQiEIyFaQ6oetJnSONsiW1j
H2lkqTnH33GJthm8Ec0hsQG7PEAEZGLezoUKavkbRtqOPwpqwTC7i2wswnoHaKKFZCdEvVgHlBVY
+yGCAsgSDlpIzSXbXwLJcwlZEpAVhNkN6mQdRaAMW0f8Zx1d5my68Kt/cHj4uxrve2KVZxzMtpRx
od9XEc/Wjwf+iRxmVF7Bvb8pejmN/2mjo/sQVSRcypaBHdZHy+6bY3efGowOd5OpywJbjtJVAn6l
gG1aXgl7oSYoY9Im1oP59uRtd2tBcBMvz5kBHKHzotyOeB/fVz02kMYPVZb9C1acLuz5pgWsYr4k
eFGhPXOYLUa9cWoT8z/Vbs7BbuDieaW/dyvNEnDyblTKb7ZJ37TTvDjd261fX5w6MwwoJZDoiYPK
0aaYQCz3McDApxOwwvBB1PEvojF2OVagwnANLgyKeDIMXbUYW4MxUG9CNxhClYun3GuELsqqBmd5
IowV/g4XKcqZyUJOmsAFRIF2NvytyHrYmMDb9muLyVxJh30omZA9pQbGbiMvXHlRxSbP4zPYtEZi
t86BoMseg7B4R0kp77iRLgaYHHJKRVZ3HOYaVTTTIptsvORke1z23nbROsetZi2Ec6VWX/vIl3C/
ee9cst/K/dXcPqMeNv6NyylvuXMXi5PnKjbcr8Ehbm0s3oHQpZdTK/jpip4JJpp+vH2uzZ64DmJM
NtHgUJZLxN15kQV71FdN2xXE9y2s7RFQ+VLJQs2MvQmmHH7ZV5BC/pH16SOBh7Fz4DG9RL4YGXxv
c0i4foCjUMwWUt0Jh/zCDGhrZf7j3tpuZmqaaruiGCgXPIuYTsKUi6XffeyU0j+QCYXPECUEGz8M
4sB9IYLVcyYlxHRHT5wwbUlFhNwp/lKStsKU+a/x0zrAgzoIu7q6p6Hqt3Z3b5NXRJ9++JEXSAd4
+3kyaAFJ8SL2lPhBmqzf0LqPE2KqydZD4n9TIc8CyIO5A155+ax44SQg0ggVMWjnqPiRvscn9LlF
OE947505Icj/edsqUtBNXCKcdVghtCbfhv4/hPL2T+uD4AyLKv06CYvAzMYbxMaZYCvciEOlybUp
lXsEZcItKHkaeM1KHamVnyo6agcjkKN+oieXUlI5HlnOY5DiN3KeYNV1Gs1919XotJvED1u17g3v
zCkmUFnq3T46mxU5XhsO3iBkaYr4I4weHHMFyDoQOvOxnmIxL9UHKXDSZR54SNQbQkbRRk69ikR2
piSmmBcFjXbdUsu0emP/5IjWHpeRJ3xx5RSOepk2ZTqgUkMl/KN3HtFMG0qaLQgyy8lU/gYzUv8g
1n7IDLMuKb1iY32skAbv+vHJfLr0b5H4bJ2cgEePYE4VXwixDQKljcBubrYy8pZv5XRhM3kDL0G3
NAgSO0DOXo6tgyUFORZlUV7b7HCsX3xnrLcI76R8BvpdngRhXNd6YgXboVZ4BJOunvmC7a5ZyTLy
X4KbtOHxaZ1dgq5DYrfmkpM3Q5scflR1LZutmil0F/fsUBpHDL36sNI6xwMlOi3RONyJD884TCZe
ywKMvRWb8iijD5gU7kSzG5IrczLA63Tj3PPtv2/f/bNJts4rbuUCLEJJsbjAA/c44vV1YNW/aOtJ
uwzXJdySMzZImrBv0Yt0FtobbdTLGbgnUAfu1QwiUFpUealv7pV8/1r1Z55nZOv6MUSNKTGaekC4
YCakGovT4FAzJCEaGPdcGWQlqKg9MeeURF+Ds3lqJM63G0PV3Zu2xWKj3DGzbbs8J3sPa1R2bFGX
aSsjQRaY0lnPGhqwfe41uf+4IjxTkbLUwzK3R37iaMrUXvEKiJLVLNvC192VcHHhdexI6Wtscy7Z
/NFkN0EaSot9YSlixo+r+IZvZ5CvlZJz1KKIWK7JQpC76M4tmi4whly24Q6hgj17uy0Pc4GG0z1U
bYIeJDgkK22X15ENuzVgnKzK1PJPl+BYMs3HkVlfFkDsx8BOAl8z3neOWZVJMMooAkYnmawUJ/K2
jpzOGWnwlQFF8tFVWItkmuUtIbec8XwQ6NEaM2j9PGe8bm2eErz27AZvji53PiKG4qS7NoORjhVE
onoggaDvKSucBlx2lZV7UdKbUnvQCmk87yvv+8feLzIQULn72uI4VraaCHlW6hws1kzTjjQSQ3P5
GrtPj7N67eG4alvzh+0/n+nzirCjvt9IA7U8an30BufDCg23N5MAU2lWPtTToMCGpj0B8yuK80D3
ddtN0YbfXguO2UnOASA6ZJZuu9xlaLUHOl0eLaWpRZ4gMvncCYIzSI8okY7nQsOUfslKW6Cdt0lr
8PornGIrGYFeXkyZ5HSRMq2N/GmCRwa4a7ZP32C2Of9t+SYP/To+U8qO58OPxRKYBJSXgr/uBJyE
BKmM4HP/KhlayLioplFplTwJKrC8JkTgTnbfZwXFnrrlNG6GYCnc8qYilycILnGBMEkpClbVYrHK
bX195wRo53Ee6gaBi5XKuA/RsawcHUyL7Yi3YwKxTTlm62oGpKYi+R8prCTukt7WVn2/LejZFbiF
uoJZ5pMEaUaQyGeYcEto9nyA9CRmrg9SAIdkZxvsLnsihJC4DNU9hoJ3OwBEGR5Mk8lexs4ykjnr
8rLFV53RCY6lEpxvcZ30KzNwMCz5LQNDGw+dnY27sYLCT/K6msPYl9/wL6SE3Lrk3JJ16oAT15EC
zT6sOZOBQqn/7TqzH/ByA847dXNEv82AeRPMTtXStGRnyVA2PFbnt1ysJc7XJQZI5onwAUtpL5H7
hLslFlpzUT2zGfNY2vNY8w3loBQKEHqolGbRmafaAFU3I3S8b1i3X6akgqscJoH1APABtyW2uKoQ
zEep1FYN1loplIIY0T1nmgpCLmnT4De1fdvPSfu/o5jdOZJQKCwD2Ir0mAaM6qryIHQhXCbcamjm
HubjOgrb2T2dvoioDpF90RXsKTkeaHeH1GMurS4eXvP+Xv5FLdrvbxNoz7fxLbXE9N/+IPLccBMb
5gG1LmrlUtqMHdLRNZj3JPwt1P2iA5n6rHUSgrxeWzVqXwXfqm8HbM/GWhfyzdjZ+LujDfZ/NTVq
/tfUZzRXIlg1RtnhvS/uFrJy9h3JksbROKm+XVCYDg0B2xSI4oq6JbweMarcCeqy4imonFPTUSfM
I/mlsu64Pgw3uxLQ174zqc7GwpKfpNIFi0bdQZOq09cqENGseFO7Dr8fUz2aXDEzVieGQy7co7Yp
8gCJ0glyzx3ggZyPVzaZrcDx88JXC4qjusjxd7Be1kEiDaTHfPVAoWaXSVeRqgsmcQBKKVWAJRij
xucKo4SaDn7ke+aPgmmL0G2J6gsdJ+mIZkSOYRsYFvyPeA1+nDdwNQNeU0OxPEp5xHKO7MlPMUf3
7XyrvkF3OvXW2hjtgsMj5PnhYRlQdXmwpOIZNJ2QY3PRrtOFGWfxAa3MWD4AuGc7r3bW7xNK7iX7
l/aAjuYOsWmDLbpfhnQROJdk8vT9B59HyvS0hQlnZwmLlC0nqqYonXidwtCnznMEVMEQ+qXmaFcB
+4pXrJxqlsyFfmpAxdlJ3JKmZfkPt7htQ3Gr9rr16HP72Q6iP/WstBnFNK+P0QvK9FVj1yU14X0S
bZ+AXhJqRkk47T8hHkIQkHBENvJV/TA8cKlEjVDKFiigywxF472F1Fw7BPPWY5QK80oQSlGxEMZE
W/AkcKMntDOiqNGrybmKIlC8NwMTmkV/141dp1KVgfAyD13symH3o2U325GkVXbb8UIP0/wman1G
k4A3UXkeXFR79ArOxLbACkZ89f7O0DODG/i9CbKsquRKeBpjvw6Iiorv7tP9+MdTgkS7tJZ4/4Jf
Ng4nL8U+XmDG6DEo1J98zsQcUB8R9+erdL+sCBk6YFQICoHQLYk5+nhb3Qjf/sMnzII1hxde12Sx
JiUzc2hW9sOiCc0B4iIJjE6nzch8qNcOvnn0+PobAsAMvS0OXU66vwETp28DUobbopC0sOLrnzmu
sy65GPIczRnDKfbsHVOQuz/dacrWRNXvX9Er+czT1yxy+p7ZXytkTu4dFQ/Rf/eazOlD4GGKVJn2
Vg0QuDQVClRcni/z89LHzU9eEs1ZiisNTzgwqfcCteXDTONJgLHPw187WH4Xof4VQ1ZONVFHxv9B
x2LEVv8eU1cqQ+wW3nxsrrcUJpRSXJn5n6Ai/eBMC1oSErCQFWS1XeWQqEs8CFlWfdOrKh0Cew9s
wyRVRDL8HgE84HsBbO3QHy/cBV3jHMy/ni5r8IoQs8pkgKq8kCfX2AO0k9aBIyGHpVFpqLVKkUvF
odqmdIx45emS/aV7L/rnsEMTl8bQ3wNWfsi5Ol09KAny7gAgWuT9lE+9r7/9gqiPjNWNGMxqAUuB
vY8//285e2PmHhEC/SMedUmdeMXRiKaoqZIxKIHA6r2vrYm5EBw6vgZ/taIqNJCvL19FVhcTkaWj
Iq4/fxl4+GMAtz5ItivDWD9ySlSssk6sjzIVhOh0UATZBwU2S24hlJC6mpxzDEZUs+2Zt6tP4f2m
toHw7ltgWhq+uX40svO9bQUJdE44zu7rlz2gj5awZ4LEhGwtl3b6yic9ZW8Pn6UsK+rm0xYWtkOI
HzGFusH46OgG+CeH8xIppUGNYs6X3HfPkHBNXn6qPQPglewIL1LI22bpFXkJKXZ0bibe9YbGK+tY
XqVVcjUv0i4k+/jsTYMNIQtyLJUz5T22N/O7WTJUoEv/DDk9yw7XNuoKL3qtVIxB2Kn1FU4YIBcy
COYV+ekkpVQcWiB4SxiLJTqpO6x8PfB8uScH+lheja8zYj5Xo4EQ1pYLnQYVydGWL+X3QhbrUjVS
xQiAiay1kYa6F7cTxW3OaSGs146CaUHrEgsnVJsNCU+Y/AAtPMPjM1t8jjciGt4Syu54eqlhMD+t
fFh8U4ukCi+iju0FNKGFZlb+JnQit/80QKzW1B4X3f79x9uzOfYO2XTtxEUVtC3gdNdqnvt4Y1gz
Vko6P3qSQzzyXWoEubjDd3Gg6YZ40hOmEjegfmSA2wgkDK2kQp3RYVLUScIkJ6eBFqyRabgNF1Dk
1GmV4HzCsEvRl3ib5/5VNVR8ulpoaMShR6swLyCmphALm5i5+koR9oHkrwNotUDEmhAYr5QvL78G
XaVYDdLpmw7wDPrLJF4AMh68dPrUvioGNQ1Oq0gPMDUz7wBvzfZ2DzpamPl3RpqEhEVdO+AT3r9y
0fkLSWN4dnE7Fgu8vtLzUzf2hl91RRmwP2Y/3pfPH7JYqRAvWYYJccD/JYl+DiQnaKg8dsllxvOL
hYqPx7g7SH88JhvMakpv70+9WVkIFwQBsq3lEIJt7377WO/XCQNZtwkTi+JVwfZVYHG8bSPkZRNm
mHbDehNbOIAqvwbbIjkaUtDihv9JuXb9V7Rg5hywwUykiKryW8p9jVMVgD3LWe3at4HRH6SUpXsd
YpUgq/Ntdked32VnNkNKI+SRHHW6bg3fFwIb9gGb96ijnQMqwtfwN4PQf+Mo4bLAAwypJymjnn5i
qfChnCYHoXJ0QHKUWUmUDuC9F16wY+FWSBpwMUSW2cXPAX8MBhxDKIkklwejqv2XSI5Z2k5gGM1Z
3t0zvVO7dazcwClMx5h7UdD2AhEmnrjKz0wEjzKATES/ngnzvhKjZ3ChwvQ39utK5Jp9DQQhpvcQ
TPMsnvfY6VDrFJpZaAfMIflWNzTyRh6Kc+7XcStmUnER/1hn+keFTmQyTJplPvrz1QUnkTejb5hj
kx4RBpoA+fTO430B7uqa65182th9FW+PIXtxeq4IAbtc4LxDAQq//Dcox/GMQuFea0kWljqS8sbp
J5cmAde9xM7UYtzuqHJZFQfU8paDE6sVQM5amAx32w/9aJfcAhoSqMLaiuoorNxJm35EPCiwR/Fd
nwszwO0cFymJkc4xxoxwEoKgxAAQCosiBc4/H/lFwPCfijbeNo7bVWzyLj9xGGGteQbllW6Si25I
lNHwq1HLILF7rpFPEvRQBqUWtQybdL9L6wa/ngcy4vbG27jPTtBOEkAt/oehU1tugiBHVGNs32Tb
YERKu8a95myWIKUSkF2Dqu6rh+8ypcWq3Gt6FyuqZi3kslucge7hoTjupwG6VUv0/mlEJP3UC/TX
xY2vdQhBaoW2wV/hzGnqca47FWp8r8UgJI7PfibjROKfHi51UUoQskNQk5qIYqd3MvqJHhqWlGLr
ya5WYJ0Qw4cNDRLLgluXjDMXtoGsY02LitGjKSs923rG996zIBkagU6BlL+xNDCUrImHjV7QW8Hf
TnDXZA84zK6NOV9nBd59BP7gs6liwvypREN1TxAgTwa0RrwuOQSleC/cYrTwh5VaAUwTFQA1d3Qn
s0rwZ+V3YrVmropjVq5CqW0CzID+ESQTfOYsXZAsbppLWILY7SwtnM2gnSw+/TSdVTqXy+oD6ioN
vgqafPk4g+9xFYaF8mU2KIUaXVSsq02h5i3NLt5zfHfRXKAhDL5VH87lCXLZkAyx+UDJjecODl7r
7tQySsnpIUZK5WTbbuFgsSMLirrMGxJA7oSjU3yekHCbosqDPEwbxumLXY6XStlxx71kHlL5z85g
SleZeiHQzmDM6ILkB629gof+ZhUMRcfsV1QjuuOzlrZYzDfmjbhKUQCbSoHyxaN/2n0PfLkoOtBV
tYFbbCBWnL8FhtJ5c5PwkyMEJSeGGN0EqPLWfZPvuwBQl74h0eb3OqQDpseu+Ch9vIFzXQcQNVEe
yCKzN0gLEQLIgoslpEwSXox1+h6Tu1X0bR16Tge5pN2AnzTA1Lh4tD6/dfr6z8gnl/3IvziacY+7
7hOb8db+E3N+vBS4pZqSQW7CED4S3Eh0g+OJ4m5glu3HrPxcpHP8xO19QDgHho/RlREeE+gKOoZf
m3R+j8MzkByc0gGUY49plI/jH78IuZGOlXcySw/dXwZqn8B1PMOYI7qcV/RV7ojeZRKP/WULcChj
ltyuGpzjUkGmwV3T9/Z+YV9jgI6/BJvbIXShkR+jvd1Tk4fkQ8xMnhwvMxd9jVbJhFIjm1hV4IV0
jV8AOFWhq7WP2Z8SNL29yTAq5aR6LmChAG/Km1NpXNmLtFr5I6V9HIIjCE9amJnsOhr85QOnwFgP
Rwp39UsctqdddWet2eBSmJQqAy6FS+g063fpjrQdqhZ+3Zi85TW/KcMb25F0xRLHyPZORSFipfLJ
Vl3k5z8zT3eVYD9CjJ6i8saK/MJGLRI9bdlMjdlhFZ1f4z/kMw/m3ODU/VzHCWuWbPpK2Ek4aUkH
5Pl0pMWdZcG8EUrSGLax4xtvuU8pHOTSoYpXd/JQ9xZm6poQq4HabKsA5q8MvVAv+E1NhNv1vKqS
dIHJ0Lj1fKg5V1vaHz9/oe7LRrdIZha+7q+3/JoANNXlSeTdPbWQnDmK4wIYeiHxAn52RPoiWR7K
xATPP2K/mpF2kGS3k6G7ikeJMDyu8FR/7M2GhicZDgLvBpnwIjxKp35d2pdgfyzlOzCrMkba4/Ue
cb51SXvdGoGAPrkOFXWAHcGOtXmGch9QByKSCCLS5Fcnlfilr2H13Ph9GPQbpVSEdp3GbSxKwDMc
rTd7YPsraAmFqdkHgAuDqs/26czjOrjf3UJME9GVJ9HrPZaizTNVr3RBwF1aWYUljL5wwN9AHo5W
6G4MepVsyfw6MdrcgSfkwuC0PZ7h19amjV7/Rzvm1xtZ2asOKA6fQP3EIpOoK0BD5a91NoIuWQhs
4xcQB0n6fjlBul2Um0PAhNclm/h9nccJ0AhI9CZEvNauYbiAeYyaA7a+wbjN5psjLDABviiTmIWR
pEQnUs0wv1s2rdYK4X+Lmd3UAO7kX0bNurpMK2RO0FLNVuKYeet6OgjgbNPNKVcf4HSIs11UnhBt
Es3wOna2UsA1qLoLvpUoU0DPym9R6ev/sTuT7Vv0h4rdi3TpZeH+cLTqPLRPuPecgN4iIZTM8sQ4
RZvVcKMnBnD/6VyWJvDKUoOLpRMsnl0kHa50GeRWx9yyVrMKZNPqqIkR6THOaEI7wj25KLSGIQXl
QYQVUX5qVKOi1GYUSeSTL0jgkbS1V8Nm8ctFtNocYtI+AUElR5oTA18gaty34rF5q+znMUWiVChf
cs4hQxhD1AYBE7JH5wu8oU+9UgNn794aHu2Cjkc4IXy58vM4eHrRA/Hl7McLTHH4SgSekZh4jNfH
J2QOLE15eRw4p8E1/h5KcJUIRwj4+pRlkIcDxwu5qN+jKVyIHFfZ3RNzg/3Y8zH1vGUqdnzIwL3p
xizaQ2m1Zp0yl7xsVTz8r2lgBbqL58Id4RF2giJ+z7k6paiWsXr5v6/dmADOc2pp78cuj951BNNd
44O0iIedO+atPCBOFvm7QGeUIkqAWn/bvlLYvn4ArYkLpLoZO8jP9SrquLxJr5P76KMKzrT/42BN
3VIg1IQdPKqKRMEmw9mSGvIxiEk3MLzduYRiFT/RHP1OSbtMFnUsXtXeBsxXhvdy9yx9J7dfy2+w
vZ7t3lOQrKMAe+bPUWyLVpu4WE2LXZKNOO76lgNiP79YaRwr/IrA3gxDi9su1Pp9bUmy+e/lRC3A
hiw7KWvb446WOWHew+XCQb8n94VaBewLZrDF4qvTPjH7iLgPqHjUij8gfvZBzArE1btCeQINHQ6G
sY5hv7F9NAauRE8BFU61uKPHDLzCQj9mPp+uRIg6fN8Rhcxcpx5e/OzDWGV/Gh4sRHYHSHTfVgLX
wjArkrshrdow1VCquABg0KnFLf0a9X9n4um0tr/UfFH0gitF6naZjZwjTDHmiKReOSz5jSCXjf8v
aMweeJV2LrtgV8P7kFwdioSspfeLKhhd429PWXvENrPSeqz9KZcbWLXCJEdxOTAIUzZB+d4oUNXA
IH/iJkvPXOJRk75PddsKQQOt6Y13aHlAQvycCH9JbDH9zkyeOCJskqvu0DkLXGFuasWvFs2tQpY+
kdfa/GP4JCPNQ8/57fU2V4am/+HANrA/+a8/KQ+R3UL5uvIfrp1r+ahIrXxUrRZDZlk3LQD8FbT6
7i4xMjUL3kP8mS1bsChMp9p2A3HIvEqCZ1k6apDU89bD/VMjmDUBDyYmJPF8btZrx+b0Ntm9ONjK
hFSiKS79c98Knc7TfqX5w2GazEKzMkxWHZbrb0NUr3MmJs1iR0dlxEj/wTvaM80IkGzAZdVYDL4f
+CF9kPORnnJPq8ltONtkpCSkl6YaLiyxhgRF2MugJerV0ET3zqO89ux0Rwsw8rUGFL04YMlyY1EC
9oGc99v/gqKTULco8sx8FfsXi7xgZzb/GLPAZJnHT9ow6bIKV+iu9WE5JEQRzvOlnlwCbYbAz5qS
tG8gKNiqtnk08JhUTl6o6fmor7G8o3C9ytKC4uaWz5AmjUMNctrsTfx71QJD4pvPEu4W6JBpTGMN
loJm/Jth7y3WRcaK+UE/F60Jrbmm4zb29e1HUumC1hzB7eH8hM/NTq2v8NDumHWIcArezbFThiN+
OheBSFUl8NpMbtVisOmTDvSmkg/1yPJkaoD6irs6OdFXLVH38M95NbsW7Ni9A6c+Xo4cB6Lo3+fb
FoeuYTtFOukzPr8j7zw+xWXSDo+Q0HYxEm+Z0SAbHwY9eqglACjNbYLZeAd02aEE67LNYsfKs7/X
K9f109r2UMUFxcjpbj4YNat+x+Jjmzo1sML2Z48DPbu77cm/Np9t7riOFJF3sAnm5VHfeWYQ936P
3/fiR0pdBaYZlGQUqU7vLDtEo5EsiI6BEWxZo6XnOB6oG2Q9JaGLyMqtd7sSk/pk5+X9oGJfPICs
x4ckn/n1SgBD1d3OiAk2QPSFfImnp0OU4MLmUEm+hvpOoQ+BhCHE1uwYGGM5lFbCy3UhCk74M/S+
E76zqyhxeenqRGZnmvm5oxiDTxHSUlIUuwmZv/0JLGMdsonfySqO0l/PBGHYxoyXZmKqOHEsCLaV
N9KCDh0gTGnQFdApHfahqpyTjrmXyQoVQVbodebVUy/930kKf9w9AcKkx0erjtppfPy6IgxqE0pw
5j542YRQUx+VaNxDev5fwpDbToLRPtzPlf6Hp4s1XpiqfZqVEs9Vwas2Xod6a5jd1US0w1T1W3Dn
w3GPxyu/yG9BAfOpMuodnPZ6GX4WT4+wzLwmzqIyQTK9EDObq+M6vfLwah+TUBD/rfGt8kFAOqr7
gxRIwOT+8TtjL1LaOKuHCYLN95Pz9v69nh2ZhSrd9frK6IT+c+0CB/k7bZ+gB3RddwYizi/4VPzm
GtnSo0HIz8iy2HrAqwIbH/V2+qh+rodN4Iq3FLmK3iqGjKCG0KVdF3Kk0gTRT989P7D5JVV7vZEw
YaFwt+aLKOIcZGr31DFduUjs07TR2895uzzIZ7JD349dx+1DrYzZovWIJcCa1xIht+C+4y7FlPaP
rKXN8uzSrB/eToD3H33aRbkrgeXUU6aZNTEOUUcn7y3+tJTgIcWGe21m1HcB4kZJK9YXCVqYEgsJ
qlT9tMcp8fsftOj+ua+47AB7N8q7lCDwSJUgy35XIx1nqiXaTd1fduaN8Stf8hhegKJmKwAe+N3U
/ruM8FoFlFjNsUtrE39PRC/07HBZpbr716GyJgHJoQcTc7lrRDM4hFSoKkvFpjgZH7xLZSPGXTA0
bsb6b8KrpAVMw/97/m56pACteCYXF3WVxKIOT4z9zQPM2TDI23LHy3IBbxliVI23E3nsWxt8qIMX
02Ud70P5WfofWk7xVYg7qU+xkW6lAoVX36TSXwbj+05D13yDURiEXyS3aL2Lju6HaNW04Yyy8NvQ
h/elUXxALpWzaMB4ttbdGktJbBMbr5F2HMsuzYvtL7BKY2kUTgbRAJ042OWi5wn8uYIlUUzckxD0
gJ3cY8zLYX8cgGdQ9K5oSTmLLr56gbT2Hc3CdRVItIOrkObIiRRwTgH7BsPZS8Yg/UD47IStZBpm
o0NaIQ83dMdmkERoH372tNdUSSTzSfbxWknOfm4rCJlkH2LpPhvhk4A27oOpQa5FsOrWSNbudg/X
9dTgmJLphm++rinmytvY1w7Aimm8iAlL4SmKhAPdttPCJXC95JCV9BOc61JEGJ51C5a7tqwSKtUj
fJTarEY9rXi/8L/gMUZlXX4EVe1InWEl4+8Y1/mPBvqCuE+fNIkr6ii/PpWmT7BhBZbiALAPEibs
XK3lOCCIjtw4jkoRTI6qnBlpyxaSvb/KzDJlMuAQ68hnJsS5KyTbuY1mCKb2ZZ5F9mO8qrCBcnAm
zRydKhigskWbQQ29y/le6Bv2GVc+ocpkgfqzd0Xce5Wl9WkuGbHPf6IXUOqusneKiQUE2Gi4LyUb
3rXCNP1o0XpnV60DnC+CWcid3irUeSSbi4EZZ+rK9/vaQxreC48y/3awOSHp/dFthMudjRWfaZ3N
QoLpPXtSrp/y2+d0bZocaGMROFgl25hLS3JBr3YTzk+BCWh6vhsMOGiChrRu9GYi60UbaORFEx9J
hPCQ+opKnJm0l0xqZhpUw2g1MpHlGUgUtwITVyqh41z19H2P9IC1rTIaDvEopfn0juP39kA2KZwD
GwA9anJTabCS9JVprVEmt9n01INqlXJs42Q3B9ZeDUyTOFUG2woLcBa5rJBYGCK2N2xgJGqWQFAV
O5w7UZ+eUTNjTIv/MCy+1JvL1LTkCppgA8luT1ffABt36AjnfRFndl5wzk9QKG+7/5PrOobw4361
R3p+07zX9Zaqls19nGgVRHTiQlrgF1eH/hfU5hF2vdDpfG6nvFI4KEnVfQBWZaQE/R8hZ+e7uHbO
kj/wptT/kDZllB7qMqioARuQ+N4CWs+EsZfox3xXQiYiUzV/Bry90sKob6o8j3p2Nu0MWkyTGJ36
Z83mCdRRKvQr/BdRshOYOA8bRj5NSViiFf2PQhKDmYiizptl2OIF6JpyATtSLG2M9qXQDbOe09bl
GHDKgOyrAFABpk9NdCO4WkdDXhOgW/YjEkAMM2m15nnWcFpDYF+tQwQvpoqVu3dxtIbv2zGJBGk0
EJetGZJR4sNPgNYI2zF5pM7G6/FGAR9cdb0hhHfpAipCXabXuHi0meZdfRig+8sEEGB1KVRipu+L
PY/WzMUBl8M+Bm8+JqBPe9eAmOfvj/TmP6ePzmzuARSV06AWoz7IR35VqZc7e2HqAiPU2oSAQ1Vh
bdK/WxFM9e/7ZUuKv17AHztD9EbKgzagJfz9ks8QKx0E37kitGc+GXHBJCeWWMDLNZigI1PQVqRA
HZx1yrGpy3fD8Nrw0vfBc4qzOKmfcSK72Bx387LKiaWSUUQULb4uMkJlJl10oQOQf2BS5hzzXM8o
o3Mffd+RGOH78k95BKJm5zR95Hg7S45ERzmFvJ5EmIy6BehdVcg8YZlpj6HIU+s0FFrQlwj80tAh
z1akRbzjl6+8596U/Eq9SalINDM0XrUm0EJWrj56O+BD7vj2RypP4CY67GDoRlGpWXmC8+4kvN0A
f+ykTRuU85c8scyxPSY7bA6gSsZXO1LK5vta9diLK94X2/WoWlPUsvjIT1fdfvBJ63StIF5XqjgO
hdhiD/vFfgbuyhiEedBiVy+npaqo+u6C65/Ui/oJ9F4skwkEElQ+Vv/wB3bYj1dXZxUbOrc+3COT
T2/zlSP24H8+6VxFi1MfuDenhJYnCref0I5AXs5J/13LsGySowRks3hG85Tp4da66BZaYAPp6doa
qZg3wy44sjip+13kAhmShE1rRoLf/fOfhWa7fgnn+bJRe2SULx8TONvy1HlOaBB9zGKhUGyhR08d
IzVgkmRSxux0FjJAhoWMPyTGz1xNCDCucFK/9njr0oKa9uzAKwPgUmBIYfrDDrJjOkFU8iq8jeii
xmt/7EZlECfOXuV//cgOQTudNoyUJ/cQYrovjJRwfKiys/cHTPgVTVeqnBYIgMsSI+TbtT0HlYtR
V1rrrW41hfvb1+TqGFnuyu6kXz6y2ScIoaY8zAZo0iMxfaK/8cY6RjOiUrR9Q9eoMFc0wTQlqwJf
gkXV/zb2pxttk3ZJHPfLh67ccGl64t2eQX+inJGTXCcvc96uScnfoNoMpfEQSM7NmKorMCGhK86n
uVmaTJqH6xFOmfxvf7sOiAJtUok3FOmfPrvx7YPcfmC2VS1aUN2/r0/WeTbJiBb7BceK3DsEjv1f
IPBaEKTCmXlyOz5rYPU4718hBzQe4nJcIYhBcw9a1Ej9MocB78ECE1aWb5Nosn98BmqwizM9dglc
5KnJ6waprEPUWjcar0GNfBL8EdO3oyr3qHS7YZFp1/yt+B9faUgOn6eJ1OI1/3LtnYIg39nb9Qtk
9ys8QpK9QhMCaDGZhtQotEb0GAoZaorrKXvOI7hbxrgCNG6EbDCrs65m5jotr/EV/kiv4ARfr/Y9
q21aLNhUuasS/Da+2/DMFjLZgokBReNZdHsCAfApd1QBDBqyZcCtd2uP4YDlp35/LC9kWQPYAz/o
DRagXJ44fFIEPtV7c7AB5MqQY5KlcyXFkI+kWUy/7aYA39TQQ0ybvnaNVS7BnhrSEjGWxMFI/2Ii
KNsd38mBp0WvN+97bkq5swULKeVXTgnU1mtkVKWH9vFKBalxpyZy+OhWU7WhqUKkIl1q3BSEKJFP
kCIIA5SFRehIFbvxx+7oAAK8UlepqFW8hOCzhjcKEn4pOox7omF8pISktROdTJ9IQpyZlfgwGF3D
jFptOTGyhc7HESm8+HXfP3SAC44uJ6KRnJagdj4KqguBQfnFrlzpYX5BdBhYaAraLpCSJt30MdyT
QjoB2tlqRGsoPsY5EDRkzxdW7bD0LTstXvr4iT78t7GWcfrIno/D5dOEsOyP9WLmTTRHNR7aKX9o
gP5vqsFiz24MaE2VMxcVfSLGT0Myk1AGfQC9GrluBx3HfzWvR311m0kA7vI/NZw14vMhSASL9/3D
TB6F7OuvGq8MaFTERRkadOV7OdjXstfL/J2xiSPn4XNjw3a2RtA61lG4fm8/YZx9jBNzio4t8eQI
n4Dxs0Op5n2acjcspV+nWe+jkS3OqUNMoS3c8WMjESZilTChE22ZAIv11H1SdbErRXaRoGvtiIjs
wDokOiJeqWrdgBPWQFsEewu7iJixtH8relJIMsZSKx+BxvwzR9P0eyOJgNcK7M4E6DgitJAO2AXx
DUoJNT6ZB7Vzez+85oTxHgzBghulPc9w/UDO2x4QfHKChipMDDiMSY0d4CvKF/NApdlqVhHZqZJI
f17m0cczFsDiZmyEaD+onYSLdEdEoLvyKW2zAXV2WFHyG5/eUQMpR5flbO7VqN2AnFlzPy04wlcI
Oc1D9NM8mrVLy2D6h1UvWWGRGYIY6bPOmmRzyWDG2GIG8AFPs8xHJelOxZW1VANPIzk6KBddY77s
xk8r7gmtIPXCQ0XwYzbDsbXCzo5CNDKwUcgUXoWvujTalqk3vEh/VIMWe56OIYy/eKVzWmaRswUn
BOuJbyqNF4QdWV1xLYlnarAdMsr09UbhQ4/LhnsusNDOdMArSWC6X6LSlz14fzfeQ71Ih6wzZsqF
H4hdYSBkheXYJeX7bhiKDEzg5sDZ+T8MqkI1p4TP3suON6f9tgRzinxTt215qWCxEDlVUBe+47DX
A8nE6zOVD+NVQP4915nqy7Amr7ZS38dOoqqY2wJ5FW/wMgQp1Yi0BaO8HV+iSllVbUzOS4gnPKjU
wPjmh+/gNmY+qC94cRu99yiyskl1uxhCn8bkeL4Kki0CGMRmS7pEePb/l6kT9E0nYnOwCD4qqLEK
ZL3IMpCHTyOLljwxhoNHDiAGQfSgEphLEoPdxlbjsONxBY2P7s7RiW5u4cVv67Qs2+fzqYo1/HkF
2jqL2VXkX9EdJhuK16/W889ClApH+1o8Qt+KlXTDu7/ne8kGO/hEPp8arbUkV4wOxmQwMRrslfSg
DwSfXDcGG3Qq/NTnfau6lUtuwVsyHMbR0RD3wm6UZtR7vXz+GmuGU0JbSCqLNNl6GPfbMw5oIuYR
c9EWgqmXEtF54Qzamrpxvgnfdn2MdQeh+XpXorr9dm6wFBHQfQPoBuMmKyaDhPxYJiFODZYF/kUu
HfbwonppW9YIM9+tbJxDfimuYcR/qKLt24JA6eDz/DRRz32+E4XYN78jk6DPUKa8UDR4xkyAT+67
xXbDqawjfvX+U8493f6n/kIx9Z04spK6n/m8c3zMmPg3PMew449FB029027Xt8dkYsHA8kkRqOYo
CV8Okvvx1JJMAxlAT/VeyQGhrdftBfisxRd0RRVEsuQbzODRMm63tAxxdpKQezWAlL/XqM8t2sWc
AQREX9ssTQfFGDKBZ9BPt96Wdsd+1BRu1pJnGXkRhDrfVWhi+S6R9YFCvCdfH9jHGYp8w6faOff7
b7um2dShKas+Hkj3CZGjqKLLzXrsLwi10YgKl37pVz8oertpZiUvFOGX6Qk77Oz6BS0G3LoXUeHv
41d4zZnxeifXVYT+iUKHvmxQj3dsEobQPiRWEiO2XjzK3TBKJ4XgrVr9Rn/YKfaowSi53e74s2AB
tsXTHCSKFiSppKaokzNO1jZgF5Kh7k0Z2Koiw7FSMYCd9NAkhWcEYxcXDtvHTjuFfD6ODgrrZlrJ
XY4GPconldQigl/2hWJvsmC2GsadAl/hJebhtJ07/XGOkCxb8yf/QSZcI7xiapRBCtMwB3zyrL8R
P/T/SNZN/9MLB7pbTcJtP2irxCZaXVGhuuUrNDSkhstezKX2G7Xmu0pjAJNar2TUC2IKSsc2Ly3X
AoSsrTtwoVDZdyIB2GK7+YV8oVXJ5y+etNXqJqEE1Fi6T+0uvrQm0Uo+oj947Z1x/JjpKBHhQi2+
yn5Z9AhNySA43MnsDgRaFyc6fpZCM4Vq4VuquRtEV/HXHKZ0Nn6vuZfaHn8m7/iZqi5JW+NvNSjI
400Qz9M0y5bSSzFcUZsWJGH/iWgk/yBkfx50FkL4caVwm9L2Y5FWkYb3erjVnnJTy2sk3FZuTT+M
I4rcqWnynA2XlSOgXCb/3DZ7SqZ5/uyCb3hRFBxfwZhIQbQQlHQVHlNbng+OMKz8cSIcYAAn9G6i
maUrw5GrUPkCof4/HofXrUw5OMGJsVfd/x/9xhhImZ4XTnpWWfVAU4WkVTzRz9GJ2wYD0cpTO3sQ
D1dq8fYPRnX21K4E6ypquMzlH8yZLNRHg6amVHUMqtelLmryyEz5Ql4nMW1uFsMjPMo/idPIv4Ho
YvJXRmbz1tkNbUJnblGaBetbYrWCbwGu0b9GHkRzTR0z42Jx8kesskD0T4gK/8/ZjXHan2+k5o/J
zCD2fUzg+Ub2SwJGJ3ZBm1qtWU8xvgZPmshalBgiIjCpZfpJTbnM1fHd1k2m9n4Hi/Nemg3M51mf
1DS6K7bKoO0rAupMqMSJ2cYyHGZcPseIr5VQxLW7tYZycJnyI7D/eo0J5ezANB91RbTVj56aFOs8
MPBaORpCTd5lz8wR6baOvWBNPAfkiO1PWa+5QbhJR9jk7Hh09u+F23RduL8Wr7BUoBIQA7FO/N0M
XIXTpYdu83s0oBc1PlOh+aZ8BhV85zldSpPB4/mfGbFQGih8ZumbgtrVdchLwQ01hwnsGWllyf9A
XdNy0mfkbeH4lQ/CXApWk1WoILximbZlhCsFygDdaWXE77GY+daTmWMtzUy+Pf3pukVSihsOhJHi
bdelsipXYVz58UlTw3qa9N3esr6bk9qqvFL7tLtg4PN8I7yZtqd120Q7B8uUm5984POdm1N8YFdv
sFyqtLenbg7r4M+1ktGAJv+q4cIim3JaJLd7697uAgcAwHVhM0ViL0SkM9ktOiP2T4B2RaWt1oYe
KmvUN/9qTsFUU9X3ftg99T6PewENWHA1uXj6PpL/fhJRTodwtmFn1kQKw3cM/9MtRod+dSe4Luyc
wBV/iw6IGBTDgjqRTt/YvmRByZvJmChLbByQM0Tqh13rwWknN9Yi5EqrKgAEomK6y9WZ+VJAH1jy
bLebVWTpSrhDw6EUcTD7r2uU+pjMPqSwy9B+IWtzs3Ljfw2xTC7yPC1qYj8lo0v73YCc++Gdh0oB
MVsANT27GtgiKf6oe/ojSGAW7IjsMLqq9ScD4OddGTkJ10JiVu3GYmJcbnzpNnIqCj+CfZ1gjcFk
I8/h/tfxzVyhgjodIBfelAZb8lZbvYAnqIYU2wOta6oNPprMrEZY7hJ3bKCnz3RFT8SAIZfZ8rQ3
APQ3FKzQoeXDUkRqx0asob/KnkzbnxvB2tWEagv9bUx156iv6mjW1W0UsoRIIzIqmLJHIOWqwj9d
AxwhhOSmyiu1YK3yv91ISy2c22P+zqEdc5kDCscF35ywI3JqcRDD005t78dJkxLWbVEVjP06ATkA
ofRhBO7+GuyyxfLWfV8HIQhi1robTbl2diRiD3bSKSUqvJcs7+zplSSWZ+7JQvC5rYArOTdlG0iB
Ga8ngVYptL07JaG82KzkNBC9uD+XrMz6o4dLJS4m71gzkMg1NB3v1fQAlG1zLewUaxnJRwsaj0oU
6LyQQ2qVLQ+sVnM9GBOleg7Mqwrx+s3ZVE79cGFUWbxofvtPqnF5z3SkHZ1AsmI6ASDItxCtRoWe
K8jL6fI5AmjMMlUIk7S0P3tKnHPwGlFiEkF9zGkdf3+mx1t2I2Nb1msQAmx42gvi5t+laAjxrzzZ
azdUnm68nBG/Sb8+aPhtVKyuCF9hwLOHydcQrPesKQEEA4OwPedZK8monHxKEiNk+ZbGgVLhEjX7
NqABdaaMXPbPCU7UDeXG1ZqhZ+abVnnMDgFAZba5WQNzPD05N1ZKx+kGwdRO3SFRKgeUwh2MgsBI
KMqOvOzEyRI5nlTvqSh5RkGhDN4hADZ6Uy4ZhWunxeMPjRCpUV2uu/1rMifXMPfwUGK9RuiIUOxv
QLFWHsO/YE+LdnYAIN1hh/Mmvb04KWElUM6Nom5wr+yk93TwELYyJX1CtVA7ZMhPt3uxHqdYF61o
e62zh53hoEHKq25GdTCo0DLMvXU9vft3gXdmKhhF19Mv/0Gw4jhsoJQWVYzTrXd+87rh2jWTttrL
UIQ/yIqkH8wEp4hSGihGcl82DKYEYv8bijoinPrCvuEYRSXTeV2ZzcGDtviipcmlVokQPiZc1mDq
KNszJNaRAOiDOrNBj23h87Th//jFco6g7V7QH6EIlRIU1zRht69cWY7zbDb15nl5a/wL16WKWPmd
YUz0M/jUealOM4E82mM1ZwAer0b6UXtNPPrWQKgudUKU4js4GIgwmaWPpTWHzUqlKyOccmvWt6lW
WsHvn87K5l3d/27TS1588hHDkB7CoYU+EBnTIzyMY7mLnxgzjviqGdJRmmYbnuRLopRPLGtx7j51
8A9L7Z33o+scPpFKWJIInD3AKToD6msiI3LWooXdzHI+L2Kvi0m/YQKxnoRz7M7eXNhCA/n84Gi9
ukPbCkFMqTnCE/5u76sbBPadGTySJvSOcT9dJU1UnJNOZ4P0ZXbbO/zrpvrUd8bsbFHVjhbQuxcz
49R4HNH+0sWIkCNYPUeYPCA0bN+PEu+ebYb9/EoFhiNibFTZ0y+oo+79TxYDE4MPksx8b3+o3Bs+
UnTD29cpsTgGABswr6bvY8h3p+Br0iC5nX5cqjTJdE/pjSQFXSQESSnqlhRJEmj8NALj7mQ1RDoj
5cU/57+xhMY7W8a0YAkyivg8vClN6oQ4RquiimPC50vA09JglH5ihnkFbFZqjcwOTRPHqLDRUPLH
M1msytfQTN2ZT3USQElRXM+reECYL9IUxR3HQIBRuWc5jMvKRMVkllz8l9kgRqWQydvTbRm02Crl
4jNCdm1pIKyHmamawzsOjikk+vZUnmjs0bglY0ylxb5JprbCFkIqHLhH8oKk1E6dXUlHuK1ScMX7
tnUexyxH71LrzVVssXZuMpAoxHE335XZhInhImQd25xkXJjL5j/xzBGbRKNtP04zAPQy12kiFxcC
CnOhQ62RS6B+wHyBoB1IQP4ATsroIOAc2aSpsaUBtLZFineG7ADqx9siR8v2eVkKi6F0EDE8Llin
NiyCChxe7Yj3z/yfxcnnGyKL5Kzm+eXiV1j1I7LIj+OoLmMSShsWhg8XDzfrJJzp1foiXxJxYwEP
VWen81w20C5gvBpUU1xJ36NXHnH3PvE9723/IdIGl8KHjYp7Sr1dK8B020QWvyuHr2unwLanOcpc
eUzhWYgVoYZEKZMFUm+IvpMXGO3BYEOErPrkUVjlNhlo1xlR/QIsCEI0aVno0UieiI6MM/VVX+td
UFifztvfrnSI5s2rItQYtYTlbyDYTx3FcCSdNiNAg2DhdNkwXP6QRe1QU5lUngwGB5Mgm9ipp+Ps
oUApyGcRxKxG1vBS+p3Y9vEqguxWQzrXcRvvqKcDYBZoNwcW++Sa0fyqGI3Ztp2TpxUo9hpkY5dO
a5FmDny03AblyrjERM6sBTT+it4t6FNRcR6dkigooEOhvg9ji9/xuRTcXVHpmv3hWH5dEveBIzzd
HYVOKs9jrWbCDXmgF9NKamq4E9GEs/8swgiuyFz2efZX13NXrNXKExy7bwpp6PvOol/ucfzE3itk
Rw6nPI8tpZdxbV3J1k2U1UiAGaGKrndV4UR9rQPW3hvsQcI5Cjs9XHhXeiDIhmJGbt3hiRqYzTZS
q4eLoeKHgVDvx5ul05ghrRr6O5xmvrBFne8jJGSzRuWaorfRWJkzf4nddNOLiqTA+XaKH4+PoXVu
JrauyoSJeI1TkDastTgphb5/5THGoSfyYxdmSWBVROUHFQ6nKgDszkE129ceiyth3mkTHybqWkuo
5wMX3RiIe3pSyg0++7e8LM0aRNkO6AA7WMfteSudxjOPYoUeDAjUtnqbHJWLapNIoEWpalsnDEtM
txdBfB2n9tk4YkdhkZ2mgk1oHFmWy0kyEBMjHvTfFMqzOMKjbWW5e6RzvgIpuOCKUFHd3DptuUUl
lahKCnibl9zUD2eKTcLwozQ4GAxIcE0VdAwEmHtHGrOeJt81m+6qMXANtRXpdrQjX88Xc00tZSHg
O4ciTT0pf4Xd14oO9ggdvmJt4yQyeA5TQaDjQT+43kxYGv3TFIrwmw7r7Y2YrDUK0Yp3UnmI73VI
dHRzPeD7Ipx4YBCOhpfGio/thXsmiiJjMbhoDbmgVp2Usgl+SfWi3v9cFOhXimXgTpbIwhpYNkIx
AA0qqB5mxwbAWVR1P7vMZ681BrIPcAce75tJnx18cGfJQYKLrCnjlJ0RDyVedq6O8fg7x0tcCD56
vdp5vDVTNeG0rt4YajiGvzRh2lnnwLYostRWhJhAYLlfrO1T0k560kbnF9XMJG5m5hkoqfl9F/27
AxHv4NJJYshH5WDuDkI7ZiJ+6Hc03MghHKkV4qw1ZnPFNTcr2KQJ4f8oaloDCeist8CIowTUt1L/
GkZYW/oFxmgoO9Qcr+MJ6GXKPLWDMQVaLjq5oHpenVn074Ys65RHgyZeRpHEtC8xDTNFgzDQ23IW
/j0n1qFCt3U3vg+iM5CjJj62HELNQUrhoxuZIriKl3bwANvg/HpjtcI4qCyWzwkrnGrd82NQkkhi
uoizRHlPpdJRW5BV6T7ckhtlt16D8FG3IGmhzfWsFdayOkZ6wgmj7hrMZYPtlHQNTyDDht7JXYrg
4K+1GqebBCz4eenTgxWDlUR28Aw+/NTSgw2DsfpiO2siLqhSlC/EKnkFHPm8QcK7yhF1rddR0GvP
yOvDlGgRhVjv6Do1JqnHcK1Mui8k5/UzYdwbVV1BzVjHQ0zvyKEZI3gkssOrW6n8/fM9Kwn1Ex9Y
e3s8QBLz3F+XmRB4Jb7yVYN+eMY492WNSt1sExmBcCfM+i2Rk6PP0MHWBMydc0m/PCA/N+QBurVZ
++4P+l7J1OH1LGB/y+LxK7A32Qu6gzWfsDuFmRuUR7Qk4x0v1+8Y3VoLe1/lWOWmgrok4u52nqSa
gJNjOc/yxTdOdn0AwE3rejtTFGMtKP6XdLh99DWC2immZDwzPwaspUProcr08imM4MyfS5gXaQyz
IC56JHb4NabRH5o6PdUP7/abGmVfaCjns61fD+t96gZjj+5jqlFVVEHVq/4Tuma4Ahf65eZsQ7i5
D+VIrP8X/gsQvmHrCK11SIF13peYNtje8emdmdl/t2tQcEDIWH1rwU+onB+hvNnv0lsHMKdST7zA
hE/wpIEYgJf+X36ponS5TUX4nQA3CkEguke6myCgV/4I2sTS5XoV0rP/4827A7+j2AH/hvTyGkyw
/KQVmaKdUxmbaae7UQreA39Wk1FEJgU5d64pCHcqMheIprOwuwe9j/5rpxf1nJo3q2SHBmrHswKi
esiDCnbG+XYQ6DbmjwWgqiC1zQwfstdFKh29oQEtICzBCvaYJUiAtwpGuTKnOtB3aE8+yuNUiEIi
8TJSnpPlQTl+F9vTo/XgMEdv1qWI0p3IWs6eUCWbprkoCHISGTe0LWNCPpvivlrzDcAUKdKSNRFe
v4emZOpIKizAiLDkLojsU3ZU7FgP/rS1lXwzuFCCTXFVzXuv7OT2k49srq4A4h0w00t+fgg90ya4
Wg7yhKh4ZDrO1vwxAP6/Okf+rivE5n6v8LKBv+KhhKv0QsE5kV6LZ3buHnji8WwAbvgWxXJFZ9GK
4C7No6y0p/zjXQrc+BmCgFCuIB7q8BVQan7jvrho6M1D8aCEqYleWG1dXJPyXQJcP8NFUZeRqhK7
q3FihEG4kVHKmWIRyplO1lO8wVIvam4n7fZAst8azX1+Tcs5/DWhOz0yggiQNbPc1BOJDodzlSSt
yXNkOaqhnG5TBnDn/g7U3R+ZCjNGYgZ7RcvHLO/yocTkFV8mQmCTFUz75FkbblPv1bD2HC28VXbV
L1Bj/DwXXz8bU5m525lXJNFr13vZIDMzuYZq+QqtEcg40hCDOfx5nuBuHIhEBAYoYIpJr662AMW6
WzfUGFxKQbdK1XKmFbSdXBkyZZTPT+rk6PHRQ4iakaxt2fh3mtI6gKJFi5TcyfOwj7+AseTRiswd
EwQvHtVCNWXC/zWCwWym3VdqgDXyQFz7B/hO44KZwgpRgJiNVzqUO5sYI25Ca7VJfzshd+ObZaVu
gbnjd8uwt4ZBjXnDy4ipxxVYLYlknW4pSUsCOL0ZNccs7fA/q1D0Tb247gZeBNQ4s/po+U8zL/Db
M/obRx2hROUcbbEDarFvVtzaYDxH5q2PgrenXVrjdkAY/bIdwtd5qiEozo19aMqGCjzUH03E4hic
Inugu41qYOJsjBbZetoZhgjI7bEm8eZaBYG0cYIWRyPXfK0PA6r8YpVrmaB0Utm8YWVQDfaL3K2G
Ou2X03ipqVOPVS6ocU22TnWiNng4aDUfE/KQ5P8MlBjYoDwRRvd7XeyD16kPBve5kUewsd8fUjmN
i3hVgXUcL5SJpqi2SFWT8Msh9PXe2JwP9Zh1IL3RbntBYlDoXhTMA9Y4oSwjITMFtSvxZpnjgcoJ
PV6Z4iHfqTl8lnCoShDf/I2GuSRrCoyJFkY+2udvpR91bV0zxZgrJA/u2S1oTql8nJxhta+OteYw
unYH7X1acGnSgwXmpbKsmlGXrRxRs+/K1ZVrygiPkMc6QaWXBJKOa01jHFJtV3O96yQhfXBuUz2X
QnFUf8rYQQPzuFjH6uWxUMDwQNHrdr32bpN/dDCzHJSgHXZ95bSnR5cK/sit0isp7FDOfbKOETVQ
CWnN/plj4G0Af64ARU2kq4qI01OutX2RrZggw9P9dmPBdElHOUuxNodqE9oDc7ivSf7gMP/IKyXm
CIbUiBlqgD5vOqJp4u25PnJHcpB3lCTmTR/L9DtcDL0BlNcMm96pb1bUpHIa4R3EWDkpGsIVY666
1h+CdoWwVg7My/ZtvRdJRrkzx29VHyxy43zVYp7FstbMFSo8YZluyYczVSxAqW3pkXJ49Q7tU+P3
T+lcbEpzeFPyoMqOtchHZHJK65zYQ9tDMG+AKNc9FCARZZJWbakYqJZVZ84CKGzeL5kZLJm9ec8z
fX+/SLK0qPtB8ELovQRyBd/b58qaqv9LNfQU0EEHBjhJepwLYdq2DTMPS59QOM1Dz9jYbBlSOEzX
r9DCT4qvj3cfjc7aCQLo3jBSOHNK5mcMNu7cB40vf7f4rM/Q/2kH9oi7yBjpVESCA8dGzBBUSzzH
HA22ZRLY9ZIHxWX03UWqSnmNTpzH0r4t8Vr09yguygLlN+9u+kU21qhQJrRtPE00cC0e6DypFQgC
EUB/lWo1WLrAMjI80J34lYw8q3D0Lj1T4sRrvAslheBrP9EzQHG8Q5vCK0WlfAtdo4b74xBgHzLX
mubrmQqd9tOf9kcW4jBNiKm/8tO8OMKn+Kgnit2Mbnjnk0j96z5lXc4Jd58bW8oyU6DBZiafTEjG
EMwwlDUL1BG1qZpunm0AkSspRYGpCZJkGKLqMuqRVfRA2w2uQnR6zEwdFuHkbv6OyEld3bTOXaBN
WyXN+0ISOTYt8asV0Civ6TMpwA5D+PAa/YhQmpMrSCLPFehQDF4v2IhTothesw8rMaEje2DTMMVj
fr53Rk1D7YDF/zGRRISrLbN2dIpEcRm/nQyXWEAzQYXhctXK4Ir1T+ERgMKfl+828MjxHZazBVxb
BfY85xAfEmTa13jYHkfR2P3zKSC2v+ojFGeTBh1c+LRLLb5rlBVP52ORh1uHKllbGJvl+da9g6/g
BoSkVW4ClaRNguV5CRP3hDsQBcRNLhu2PgnJQLwdzFebE26XnpNAlWoGSeCGo+VZjCzWFQXqRhMv
TaKjkSWT3pwrYA6a8CtdqPiUC9Q3hfwXL8/Y3/bj/SpMFEh9C1qddEZRzluBEgdmPzD03jS1IuSp
aTvh+OwpTVaB5TWaWXwEGBXZw8yZe7Zi1kjdc9PljVPQHdGvOB5x+5kR18GBshIqH0Q6xLzrFeU9
BhjmTvFXqDKEjWctKlGCXkzAgctTQMZvopudLujYli54R1rL+bKSXwfHVDj7gYj2kwNTUrIGNa1i
n/Absc9jhBnC1uQpIIOjLrmMVUBeJNu+F3EL4MLr5Ls4N/IlJ8ovZ4HieCqUEPDeq4FLNst8DUHi
r0/qbvlOXQ3CKogOa/7PApHbfHpnMRe0lYgR4ETATL7JAOSGmNpxrGGNl7ke0BsNoFrE5ledePuD
IJUGRAtD4ECQT0iYVlk+E83d1RWtNoa9+8qmCqcylwTzgFptsqrS33jm2JHM+mEk8vuTrcGP3eSN
wG45rKt6u7p1B0jJvyDfMzB85NrCfzfi+lzvpVAcCPV8jbo5JlVXn1KiboZSJMIQ8IJ5VFo0mLbL
R2aMSnt2QRSQumaHpRQf5xZNJ6BoR4eoSrDztns53/AKbB/B3JQX+7XSjdurd0kv9pIU4PDP3QBI
QC3pchYZgM3kpEbaY5LmwSK5iK1tuTy0+IUXpbfgdS/pz2GBJI7PSBUzJxRiIdcpzd3hyhXjB2pj
nG5bwwd5mRZWJWQtKaXdS8ZTEOWVNqD/V5vocY32voUBQH4F5Tf3j3XaZdHPfGhfMRrWhx8v8h+O
t2Cxtj2kAiooBNYkgw/upakpUvXISRFvEmzjQ3a2MQqjP4EfbRNClgrbUQ9MjrIrmhHdT73va7Jl
0WnIxIMZ2fT7lJgmGwK7k/wyEt7q+hq4gFH8tdFo/+spG/yD/6C6vtsCF6P3xAylLbDIrDtTD4mP
9qFRDR04bmvAACaMWqnHPlL/1uu6dzhKRSsN3UCCD1IOsExKS41yCoMQflJLNGiAVeBZaojnL/gH
CbLdYA0rYaG2KJF0bwnAh4+VG/d6rSUQLvXwTrT0/5QDbejv42F532JBGz19+d8zVwZgIW6FrHQ1
GqZHYTR9SV6U/EnDrHgNrYlz17NBVzw7QuEFo29IclmbtmYoFpu1Gqi0VuK/cJOmaumPgBQFywQR
fpAkW1ccg15XCwgBG25O/8J3z+f4XOCqj9Rw2pb0lOt2ebx1ofb7EK4/YSvNgwXjuZ2JRCAAmp3f
NpSKBbt+UpZbSkh8t3gF/JmYcsZ8+SeGiTNX1bR48s3vM8SE9NGr2NxvsVXrLFfAr1iPccwQ5aCX
DazUmU/PS+C3qyP4D1enkPoqFLEoAAkLbooxZGisGBS8Sm5DRh/qGz2Bb4u9GP8kUWI08MuXPi6/
GzNVZFh+MTxba0+ans0Fq+e5cGcwKtsL+gmJ2NG6RFBs0iZZhCn9lMqVEfSpyJyZ+/1sLG72RZUc
1fwML9NeorQzcsZ24St/7ZzvNebfgSHLdp4AkSq5LNALNkm+OcK/8g4Bp3MNhLhkRa4pDYSt8+SD
hjgAUHObI/2hJbAEVs1nYbwwc/DUHImieg+ZOZ/BCkZAsPn0fG1kz/BcjvulhIv8jSdNWB7Nw118
JO/BUC/vXswxxw0zfSVC0JDCkSU2AePwo9PjitcN81i1Bt0Y2LZWKhmUDziwgS/veyrPnWF5uveD
I3vIMv6ua8wx/irjqSeqXtPXERPpC4L6BUYAp0lg4PqnpSCeqPjqfbIGqhGoHGLtw+cQ4c473s3f
7ZV7jcj5+/EEMDLVOTwfpOFH5rPE3FJQCn12SZD7+dTU8KkWrvwNTy3cUZT5Vk7kq64BxXxACcuz
QOKZWk+shzMnwUF2uxM+G19TTrWF6YuT4xpSzWhsRjDUl8TI5nDyAi8dIXPtkXjaKLdo97+MhvEo
bmx4qiR8v5vUjiSJ7yPKpik0uucL25J/cHAQmt1Np3V/Y5tz5qYrZpc2TzVbhwhQvSKaSJliYTtu
tmGlhoDsbTpyZrnvSk9cwnZFr3p2we6v/zML/uylizbQXOi/7A8wGwrSdSNJhQv8OumS//HvrOuc
XbNya8fLOJljko3eFmxS06TWTv6lnBJZK7c3ljRM/mEEpYifJrahJM4wgjUnektEZVHriSACAjOP
ugGFdIlCeWrkYwA3HER/gNUGEn+4CY9a7bcSMoPPrrCGGqqiUH3SZOMQVh+YG26FAxi1CqDzXHaN
9OvMhKdVN8xan1agospf/q2IlUgkKaU81Gv4zeH2ZrPTRpt/NTNbFwaI5xOX+eUqgz/OEgfTyrd9
OGiLWwmMTN0RcbXV6a2eVXzUfpLKekqWRPGD8MyfoozBLHi/rsOnUUIo15Ei/TDc0mleOaUvM7Wm
yXUQFrhnKnf9vOKIP6e5OK65ZTK1Lm0RXrLiGSKiyukKgc2biX5a/Ljs+8vi2FrGDRvQ5nxrKJk7
A3LZ+uxiyCBMuPaH8k1v4m/Hexx85ea850DN51LunxqF9YnjhtcaHdZgff76Hbyl2jg9gCfQBiUZ
B9iWFfFCqKeJpWE+9OKzCTiLDZ+UtCtJZ6s3cupEGjgCy8OfnAqV8VKnJFHvQ4/As5dNZWB57JZx
uhz5E9wel9Mr+YTZVchH8fKTiHQPaRjeTTTr3g3FxjWHzxnwmpLGfA0joxB1nd1wlllJHs3+PRT7
hnwtEoEDxk3Chl8NBWNzxvgd4aX0r1CLMPFMSJT+kzx87JUwFauZahhs2kqb8NhpaYM60ujCkNJO
mWrR+rIo2XBDDbKbPEnjs9S4cyEKRfIchze0bxNd3fX1u+V/Wm6AIIQYgrSo+8bB+hvHSwLB+iW1
uTmfxXjUY1ij5BuTSPFWryGKx9y8XH8DwgxX3R2R2rlCwj0Jyuy8BAmeE8pE6G4RLe68iCfvF2PM
dmqYzGnAknGOnzIndjcq577701g7dsnTuPu5JcpuE7KAlcVevf/6OisGPe5XVMmcMJFBOqQY5gaD
NToL4oONpBatlnFJ9YqrEJm3lgZetoD4KF7vx61fkfmFVctTEv1GsA+BupMJREi/EYN8ZhXPnmMG
u69aIIpJJerXfYRsuUuMPQWIY6lQDCTRcdYNN6otFboQtc8UyhEbaiCP7xNWhVMzSKl7XmIGyyAs
hJl31H/FUChFP/wlAegAb20pCFaJ4wBZwLgFXbF85X3XaF7J7fS8aW8Fs+L3ZeyiVlfUNrUu2Qo5
61zXNeXqCQVQMNipNK+jzpGgUDAoiIJmZe6waghqnW8KlcT0wKBXkY+MtptfyVNJhBm6WxL4PkBl
cXwjZp8RfKko/2JSvIEdzEFgvC2rwjFGsKmWMK9C7OnBRfpiHCmbrBdgLd8jTx0/HknmHfVxMuBy
ChLB4yAjKoKfNqxZCo58U/fGXFlmg7dHN+TXd5lVgnFktW+x774yxfuf5Dj2HsVFKUpK3I5FDNkO
Htis1Ahni+b1bfCT/uiwSiSD0AOEzyfE5Zc+cjCciHjdgkglbg6oX92vBgC8KxDeQN7RrpUrURc4
u4PEMNAcEUHH4zwGCGVp5RcXR15kPEKqp9JpgXXHZUzz7XWhKi6PGAHlsdF4EnVROmqxiZlOCLa+
xxf6zMx5gWUdeeZxRQ8cHEbdEcG5rgg/kXWy0+AdF9K0DHoDaOC3Cz1o9HyJ3+muPCPJpDiPsaYM
J5KW8pWwWBDRQFS+RVT1kiDr/I74RQU2Z4trddtkC1ETi0XVzIxw4vq08KbNKHJGv+BRC5BxsqXX
i5kbxPCI9T+ScC6nxdSuyYmydkmVOMhl78/YdZ85BeGwk5R8gU26XN/YvGvyY7xpOmx0Pud45a+5
aIttxQj0S9aQrnWE7Ln7ijonc28ZXT4DpzSwS3oMndFXpYiE+cGpSL5xk3767s3AqB9EqnzQPwPf
ANNI5bFdVEjMPLFhF2NB/12TU8Ijcy4xFKa0q0YGz+h8PPAW7oWbvYzBa+GTUndtW/BkdsKgJ7GG
o6muFlJO7NK3IDM4Fu/HDFdpG1nKX7o4yzj7Viu4kTs9wH+RItMpDcyZmVr1j/6p9hg12yNcuCe6
uMcCij4sPvbCYqRJv8ePxHQEMgbnXN0Bn/Uw6DFYQm/lpZEOJtpyc6RTDe+JuLxBdZCfXG4Intrk
pRpMuLrSVQpOO2Lb9exl1qpC3uKwIGNi+Y8+AN94OiN3IZC4twnHPzV4xvwzXkDNMV8RcfP9TGZa
Mcz3vCdkqRH6qzmmdfa40ihc4D1vRbo7ScruVRoQbkd7fyskWXdTf0/mx6+BYekCCoFVy42ybeXH
19MM5pXBNsPp5SHCfRKR1Cgs6DVKtjmYEwo8XFtVi+DyvgYIBqbVrQTU0ksgipXNVBPT6KMsmDyd
ju1Alhf+ygt287pwzvbxTICcrd71USiCz+aBj8MaWc3udRmvDgSl42iIV6GyM08Kb9VBQTfRpYKO
yvShqnZ5KSQ5/DLc2oEC5qUxJdeYBtnV79IGNnbqXXSEhUe+4uGbW6ZlKcJMUkPyKUuaak1wWH2E
JFGmC+LrLy0+4+tPH2JYmtUcf0BG6j4+D6QthOkpl8Hahyw0UCDUXfLoIH2V/xGHIv5CkDVtRzbq
veBzkEg/cbgmtii+fv6xl+D8zS3U+XDSJm8hie/1LQG0s1B4ik/kO2T0QnKus2bCENYNF93ERZ41
gmd1uYpGUbvL+89ZmB74FxAK9nXPnU4rmYxN22Qa7VND97FlirpGUhhgwQVfjyh5g5/L7ZgfU55x
HuDT2rGYlDg/4Mi/j7GpBZk/fcWhTDUrdod57ADGXRPaPqJBvuM6DIdq65JJDjrSPlck/V6u1JtD
PNzJpGUQ9N3RKQWyDRMeDK1OYTmuhRiAyYmT7ViCcnmCYQI5phO1Z/4s++A3hZancqarNttOWfY4
NYGS6LlamBcWp51x4cje65/hNhl+y89d3Uyx+qHln7aB2g4p8HAhGwf4zmQSj62MQRwZvPShL1nX
reUqPY8q+cxaLxsf1r/7TgJGhDD4Dk4fSYPm0X7m0E1XNTibZ0ABxN+6nx9RMQJsmDk05kRWN2ex
qmdpyvaSF9YyAPBfMVlxAKs1kJn8kzemqWDVIpE2elfR5Ywigzsu+4zFnwTElUGvUFUcyOl9CuG5
OaxvYS0X2pWp2HvVDdgFzgna3kHnyKTcOQ0L/Hi0j/SzjNkZZKud+wg7w1HzjydYGb9tZUVY28IU
NqlAFAHjw8UJ61Y6jPtbYpKLxAW7z76l+rWK6o6lQUtyR6FvG1E65TfT8t5p2bf/GIOLu24tGiNL
5tDWmto7Oi6GEesDY1PJU1i8y/uCUUZYvRKeHADKU0AhpyxIyhqSuBXcZ1Q6RPVwJw+By6cfSBYW
Sdrk7LLIM5kRx5kb96tPsjv7YiA27hnnd7///h/pP2JGs/i4B7N18w9IMJGe9w/Fl1XayBtF3Uic
n0p+C5W9uokwQ0HzJ3MyrTXoTtXeqPOStuEAQbou2qo80DHI2pRAygjluLAJ20L5fZxxNviyB5xA
D29sJW0YpkcnSuk7w5D8RU9gqpaTz4iVQACKOWHP4C2EB2jbEX2IZbRRa/s33IdrYhv1yqkYCjlT
kXVp74HpkNaDnzpy8KgyhCM3JtcifEYtt81023sQf/o1FeiI1MKZX8odn98nejREm4TJ41zCLJDn
xKhNynwmtZRHhwxEgp+SYwfY8/nuH+rSKZ+96DAn5CbiG+jMBTl1xOZe81UQeSjV1NuLvOfcTb5p
F8wVJ/deaOMO3CdeSLOvWi1xdtee3X4Ho9w14wUmRTabtnzevKpBCdGGXBpREchqF+Ji6UcLb9gK
i9zia7e86YBos7uIfz6SBXzV4HeVe4a7yRb3L2iCQByDUgfxad7vGNFcUaNXn5BmqnzVkPPmdm6T
VjhuPjqPg8R2PzOe4Lvr0Mknr/nsJnyDWQXe2m71WHR+QFoyvZcNIJUDMUmEYD8i3LxbUehWxu8c
FGXTB4C1ZHhBw0BJGVoARf3fgQLcXWDnQqvqQjqsUlySiRWfKO0y2JJy5Q/HS40vpvSZwTvIdZZM
+LmqWpA4RtYnF1YMHyWL5OTSRzeikwLxmu29ymFy8XKWQC1m1eJsR+D8BTuL3F6Xwtv/bJRbVI6y
t6APx7kmsgx2+EYx7Z9g5rA9NNDK1YuXXICw4GHIStUL06lG6OS3xoGri8IFtMh1QCHdGqfgTshC
l9aEavwxED4Kgu63+i9qERfhq+VYzo5BH/cP2nBIj8jxKF/YLlTia9i5Q4FuMu64IRH1nhi+7781
rmsTODDoXM/b2Hz1gxx6OLdI5H2uNX0WlArMXP/2+IZlVRICm8YeUOs3i9cd85snG2itJQCFd7dt
AcVL076R9wCvvSImwrQzkTz0V3QbE6kJ20Ng5t1gJMAp7qNdyCCEE6FJs+Sqs4J35y4E4P38/OlG
9UCwHeXaM49y4QhxV6fb0tRYSQvfR37rU8JGeIo5AcnutwlIukR0JjrjsRezR8lgcwA5DtgI/i9A
A/Xg7EGpCXScvvj1XidgGjatjbED+WkgdV0Jp04xpGrkg4FffXe+RIy9Tlm0egc5j2mRBaLsb6TB
NOiTa/6k8882DbgUqX7gKfr5ewg69Ot3DJR/tobqjgEYhxu2viIy7vRjEFejFCHWjA8xjpsJLN+w
XH9wP8yG7j0rdmWjiHQ3ZTt62fD5scK3dzhXaIHD/kJB4XjL81DfiQagpUH/4NT7NidGmx5pAEAu
Dv4kgyQ8Yphak9t0ENCuYJNFQCOrPzmp1ymrIZw8L6mW1UNiBREeBfJRRJ8zou1NEVR4OZEhpBzo
4Wy8KxqwWS9zDhdJOfBtjbCA/iZsI75bZ3xPFNmtWm4LwcqOLYkCHIE5km6eKmlWeqIY/dSskIkv
LV4sDQKpwNMTQJG0YIB9ZLknMsZutiK3JfqaCDxXwYxlp/X0XRh5W3Bzs6PiykoW9argkwYQDrH9
XK3xkCXtwHLJesaaaplCQhi1pvZgW/5b8XnlhIXc/MLwl0fDnKcmSLmveIJzVWxgyF28mqr0SYKi
lBbzMI6NGdtSI+FBvQ9i4z9e5iIbL1CEEFtb+rbEN3UysoLnMW7fHEwO5OjrpFK35Z6hbt9xgdER
LF0X7liUnNFDupCsyr04cPgesHcCc/x7hNe6o+oGfaFM0lkdCz2xP3R+5OHAYSR5HevJM6ocGgSi
pk68shtJzJLPJWRvJyiVYZWwka0AuX1AalCzTLstbyLswKz0ln6FTcIPS4akWPlvsZ9FgJEK+9nk
z2IGFgmUQIgjuD9ZWHX8MHiUuq4aFhsN1rMavoqutnDJLTkIN4KtUmO3Xy0m+Z3+0V5UgyRjjhZm
1BwRnQiOAs/MjrWBX5umUwxVdc3WkAcxYGG+VdkG43FVgkn4+WOVJdt2cEvedRpbjAeMCF0/srzp
zFar3WvpXu0dHO+/Y2kImqBsphEVkYGVuWGTUUEx21LT6rawrpOZZNfvv6i8U3dilBIOuMcg/4F1
eeXQTNMf1RM1QlfFPHIza3Whu2v0MwEBA7I1DZ50MGbxoLWYR9T2iL196Xy3M0bmVYDYQ0rIEFrZ
2f6vu++Ql9o9rWHMpds3oa4d/q4A6K/xRjjRUNrcfhEswRNBovZaHTUL3doqmb6NPRKDoQegWJ5U
TZ1Ew44ofjOdi4jR9MTP1tPJcciECjbt31UxKckmYakiVaSInrDPIh3B15gIN1hwx4kZgsPKMjuw
Uj8oO7B2ka1pQiYDi9zfqxy2qS6x7SBQ5f4Pofgi+zqaPHYjdPxN6TeNvxNkXGrQiUMG9oXv+WNG
0DQ0X8vLp+0saQ2QzUpCtFTk6IFR3e4RtBBi0/RAjGLEII+xJxL24Ag1AIKoJZaXYJRI426357An
uU5WNRcMr+zPbBe075/q6HDOZekUI5UR3u2f7jxUeQyhNxxTRn5gMSqdx9AYRHaT1XsOzuouCxQE
+RR6sAxxqoGlYP20itEeVJS52R42J8RX3mYTLrxcOStFqh1Nq5lEkliXk5b2pt4b3gOzc22aht/L
3qiEItsqHB5T7g3QWukmAeohMVYQh9ggcuQQwftQqUNzFfc7ixhNcC1gMncyUC6PrIxnQ32pgE7a
7zUlmVz8UuevlqIK6Pyly5Ewgm6yo7AG17mPApVeMp9MHTSngc7QVRGiqRugOmIYzY9H3nMtRMKm
ds9mpWPzjIqjRvQMYnMiDEOerdAx0gK+V6q6tLA9JNArvYF9t7/CLOWZoDMJVgGCou5ufcso8N03
DdIOkvmxm6VczWenRpvuHAOnlkf1u6f/gpTsx66q1oOk0nQh4ei/H/YBmKLJDNn6Zi1cHHmlIwto
rCm9WnRAE63y2iNnHiEhkGOb4MiAqaCgbhktfR1m3Qrg+/QbwvWzmLyeubSLMAISRWljO8hhagiK
Cp7lOBb8Vc946s2/yqRuKRz6Z/8hvUaFQbiMu5bQJns4iFChT5cIJSraVdh9aqbRIcqe2Y6liafv
bNSKNpDkL35V7Np64gGPPLmE1eFdlzAZUkH+Edcn0NRV1Q5YHf3kQhJPj2P69+ZHjUTlrVLLcvdj
F3PVIbNkw6VT9WdNhQLVR8z4TDOxunuLByTBTe/72rB6M0FcE+9cmkhjf3UoLb3bfIuYkI6dErM9
XVlTMYVakAoWV/V0HKwjU+I6pFt3eiy1Pz86T06ivvNqj+jLM6jlOPb2nSngKY09u0rI6HFBkaO+
KM2ksfWYOW9Gi2mVZbwCfKWgRz/XXEp6ELAos9oc7Z/chUDCVtTsr9H9oWAGY8lBGWRaflzipmnd
+t4QY7JHYCuRFRvQxR45CO/a87XpXSr4oWEO9/wq7mqm1HL9oJynNilciFxI/NiWtrIOV8GZCqTp
B0+b1znmgNieR0XQOSejzoMQS4owgwu/ywURxx9qPmTNpzcPPDqIR0WY9mk4j9BzhoeN7Kb2/Ufx
Hk+9Aaskx+zk92aEKLHc6R44RGUbhpZQCSRqVq3Togj8z/vlIF/C+Tjb+qI9tg9AUL+SZWARBRt1
GaK/4OllNeXejeDbPU5eu03iBki+MSd8w81CAaQ5jFf+kWQO1Q2ZxTmEQWXJvVzo4R4txiiWCdUc
do1QitYriCeMBa8W7tq6rqE8/qPyhgR2fY9qIthtbcVPH6h/KoKJTWZjvIMBkydJMeMCGW8Ctc9j
lxRrVgVJ2CKG6LT2qJRS1RaCgcLJg7hmWFw2GxsB7de/B84oVrj4aZeodb48L3JwpbNf5LjYbdcw
eWbAJWo5HMr3oL4Rj5aErwEEoPJFtDewTfg3/32ybOtWGST4TiMo7Wwu3cQTCJ6g77gp/ZjD9+hM
Re3gVFvUP8wwkPaSDbUEVJimmupXS8++FrX+0rpSRxuMosK3FkPr1UpKeokNmj4SiQn7O9pcAALD
YWibBNp7G1bYbHSbvDfpdTg7fF7caZN+ROIkGYWZRpKpNfGR/XSzpyH/nyCqmfIYMey9tGCl1hpn
6Lg+uvHodP5rJqzPNGR8tDefsXlpKPdpbAqdGuu/ltSq46ztrqVsooUrHtOlsb3qJqvgs4Dw87BM
Kpev7FsP77rTeGBhQLGCsmmItheATTv4zwE15Cxo+H5ArsdR0ChQq9deeIC18BRKcaM/b8NTcNJq
Kq8f0LQ1wH//N759dziBqklc1fwLAegzCdFObIL8lKoiguQpMlB1e51T5umf1Jb/unMeEX6Vmy7o
OSnVouu1CtQAWL+vzMhcIAME7DBWCdBygQoaucx5BtYEoGARR6CkVHNLcrctjvKtnnSUnGDhcRZw
uPn0/9Fx4Aw8R/8HVQJmf0o1j6YCkFar9q1JNrNgZgoWiSSI1zmutVyPlkLPiP4E2AH/PDlRbxp4
XmEByG+0OOtN6b8C00Vvn5zIoyzIeL/qtBrSfTMrPkXsBtygaOwBpQvz48tT0rRYt7LKsi9JJi2/
Fi1856wR3ZmOTB6Un6HVtEqGmLLZCM1M+5GUHoa7uIxCbn9WI5ftQGTO4oPVgbl1tTWjl5e9VS7/
TJg0CAoVFp71C8KVMRAvqYeoQ5FrPc8dK9Jfm3OpvCBOQJoXTuPw5wCAJ99QqXcr5959I9GX3sSb
entKItcXetixSAO230ucHRc+qsT3/GPzeZvOuARh8YspZf9rbzAuokdnwBg5iNSgfX/xu5lzwSgu
3ykV89tmAl96OZdIZwjgkWprje4ovhBkT416/NRxb24UjDrfr7oGSUDSDydoE/911dzG1MnM8zfS
IrOQNuqkTEpy0GGglrTLPoxDzEd3vmtz2ZpSunZRVJ84ISBRA3nmov9MbbkendQs7tOeQ/+CkPy+
ucMVUB4PbB3rrQZ2dbILvyvcDi2Tc+VnATFEi2GIJCsFCfROYj8pkjhvEcNwiRY7nnWqyqF/kloO
y7pGqfeWaeF/6CduS96fj1ulI98SeUpk1eR0SLKGA0p3E50mkKoSS9/Ntl3yNtJhL8Z2q+2tBf43
/sZVNKH1c5rD1ncap5NvFUJM1yGL5iISn6s6+YoLcl8AL4HW4fb2UgRbsuIx+LT9B0J+J5j5Iejz
RZGCt4/T0DAB52sjbnWFlnQLNK6z3EtQ0LMgiPi4HWgZDCj9f4FFQMdGy8/RxV4oIRJBdkFS86Gi
uUNmDaIdu1emb1q28hwI7uOwhyBOHwEp8gzOQq+cgcNPvsVzoW/nGopGdYHF63jynBqFhlT+zYZk
iqf/PRZ0lZPOGSKJHQzZUVsTjwIPMt1w4fUX7s51QFTB+cc3ABE9/1AJ6pHobA+OCB8XyxHiotot
PZ35oQeX3dMWe6QzBtUEiXTB3/bYczw4afQwHISGIDQ1/lDyXx2kZRI9BmgJiUq8rlGVQeOzV4Im
MjVcVwl1m8ENnz2EJx6CHY419LicXw6/serj+sxZHNw+tAG0GQKVW/qAFG/v84jnVmCbRhaTO4Wr
8OlahRJg13kzz9QZLv7MUoGjRBNi4UqCJjtZKTxO0JDVyYaCQ/IBvTo9jyZTpISWR77a7U+hzkuS
8PNeX65d04+sVouhL/3WztquAqj0ValCBo1mKeSG7IyOSkntfoRenFZqhRuh/Qoo54cgYBR/Xmti
rIvdEBNCD2G7yvurXCprJwHvG5ahA1vOHHeCV+mQLPquotJKSN03Dcqtyu1eEOygbRQrX/mgcN48
WhzAvEETuBsmyz1yBaL1jxaPARs4pR2AxlAtNSxzZQeCcJw6r5D6lvi+WOPHBSi39XEAkG2lXN8+
qKoPpGJl9nsR8r7EAooyOCriYzgqO32olqRrsH6/6jh/qFrUOAwGVgnJooXRXdTM+hrSFG/CjfZH
yEsRHDZedN6l6DKEB2HsmcwctOCKPZkYMcO8Q0gOoqQ70WzH2Vvec7aCLrmnv2U82yYYJxLpI1Lm
5vi6Xmaiwo3fisBnjmtuVqPw9vmjt0jfQRCu9YC806cieXNXbyzjkrOxfShdbImZ6ryE0LKo8dEM
xMhTVVKk0dKXoD4MMebtXHL92URKItfl2kFgeMxSVKqZxeL8/SApFUeWkftYxoVqfPVe4K+/YdSF
6huJHwKBYfY1B/Mq5xbJaVRj+I2aILFbQ/Iutr8odcwT2bslMS6a/Nq6bEdKqwg3KAVkaqgr28XJ
8khyfLsCmL3vAaphL6GXPj/yAHm8qZkEfoVk5U8AeqSD2VMFKfRcwPS5hwX631CLhzyzABvXVNeM
uaQCyG7ODMaLP8N8wCFg9/rqJwX7qB1wmJnBI9CBAwo60VaLwPqnyKspX/jhg1wdLqKOVuqMoQ25
xAcRVepkDlAUXjswOq6uN01wrR3hQ7GQ2FxkxiCHeX2KxM0MaKwnbXAGIFpKReAAPZrFt8YvAZn5
/IF6HRwnG7gMA0SAJQM6f0n/506ua5XvDzUBjSxOROvPNm+TH2vCM8XANKwnCSrRaz9GiiCYgyWs
hOSdb9UqMHoYQbg0EyNTJNfeuWSYdbxeAxzUukYL3jdKB0mI2cveEuqzGHwxjGmwC3xQzlLvtzO8
4ll4g6wA82Jbsph+y0ukFTvogWyINcjDYbEJyDdB5oRVQvvtygkHgCiyZ7VMY6l553nBw+fe2MVb
jwhl5U/6PzXdr3Ajyul0IHMguqTryzfMletzgHUf3RtYoQTJ9P6AlEhPkdBcm6kH0hy3oxYx4W/a
SPurcXO1rE9PFKExgnh72EHkw1iWRQ0Mc685zu9gIAWwO1mkNL0DrJrZPEwFnDPBISAmXukUC511
ugKDamwKzKnYr0EkyAV4hkMRRMMivpzGcvm0tlbZwAgKXLMxx9XkgroWzrGemIAn3UJzS5jWBPE6
75R+EsFQs0OEQdN5hlKwo8Ms4XejprGp2ESV3WpYwLTRp8S57SRKkJieFjsRubOvsDi9thVRPs++
TXIeojJ/zzD8qQCqCoaCzLNFUwBLGVvFSEyRVTwdNhqBvLfz2ve9uGMiLZaFb6/w3UXSvTvn+9BH
zeT0tVo2dky7jkJASsdUj0pd0eQPwcX9Cx7z0BtFsN6ylwLw2YYIjxSkW8rADt6yOBhwHJXkBo16
wfqLcM3Z/0hjIl2gbF0caFmY20I1aa8mzqHYHGfDJP7cIFP5riDsV7i4Y+i6qJeG9M/1XMXPG1iL
wHBwdySpBTJhuCdAXu4jeVk1+AUOpHEeiHEaBKxeZsT3Rz9WrDzo65Yzj02qNlykZW596np7I2uZ
jQ+vfx+HvYsH2QcUwb9Fkm+gH54urlIHzerkYiB47DfAJ0JFV6ebXaOL2inkMKLAYfKaXrVVa7cC
Hd2eIkKu093QiSvZeJLEmIay2WKNqyjMaTsvHM6zY1bvxIHmUnzttsjjyCrTnjjbDdPz/xZrZ9m0
g7vk8/pjRZWB+hsv2y/ozQCb0fB/vDTrEmRx3MQ9xJOM90Y/eqVF5m9ejTJLVb99y7pjt2ov0r91
Yi+DT9OEHVLMgBb5k4y0SeomV2iHUlmaGItRz6FSQPVPhyOflw1wUgvQX4flYGr/IBw+7Zx7PTKg
Jln6/bGqzcPFGT3n/q8snetSTVA0ontbiTmH011W8k8X5Vzlu5DvgkN0jWbJDdNL2/8fzPVN6ust
P9MEl9Uz6PFK3gx9ZD6UG5PqL4Gk4kGXVvqZR80r56pc5jLAz8Pt4E5Z4JcP3fgXK6+ENAemR6F5
iQQWX53xzAFfFw0csqcB/Dg2o80VCQhyVikT+lK9lBj8ZS+bhh9AjJJiV9vAYD9KVDiabXj189DU
YoC+Vwq7UtTuMVRRVpVKDhiLEnkEIXQpHxPLBzbFugtPwyzB4uOe5q74UjJ667Ob+7gDBZ9CliYU
PE5WXEt+QdoR7ru1aZ3gsGVtHfZfj0k8jvFzA/4zhfqCcQkik+shD198bJGO3W2UNXH5M9WHh8mt
K9qzbohZ2HIs3GnK0TWo6CJPiYba2QWOhd5Yhq/wcRaJ3nr4gvGOA2lWnV6O2Q535k++68CKLvsN
Wj22iQDmkz5KAg1E3hMPlDxW8GCpt23LmGJW3tjvmBsonFnjrMSSkeXy4xynJzDfY8bNpQ+I4+ru
B82uX2J4tDTm9aUK7UmHduhn3LA5LqnXDDaRjdnocLTjJRFYsrXLEaC7vw0kvON39whNwMXsumwx
XFoWjaUcJCi6HgUMyA4Cxjl1DFDUeQXCfr9xWl5Ksbi1UETfI3kSCWX8LyvOaL/ypIbOIhN51zBP
adYO22+sZZCKhIfTC0P6B+L23rukcC05Vp4knRpXLgAyWfkh+0+CyUerVQrCHJkLKPvkenjsckaI
xcq9jEJmEsBeaTwevvHHPm+cjyOYLvaFmB8lr8Pz4qtgHGbg4y+TCvQPlyCePpBQ8Sd58bJhHFRW
yWUsgBuYvYzXUkYFBWcLhqfW9CwtH1gR+GYDGzncrhr5wQB3DG7nGl+kdAbORE4QCzcybf8xD0/n
2N1UrhUUFPjAODLLnqZur/jEFM12z/SKBzPnbCZWLNuM5FPCLQeVKClgHY5nHuIxBCK4+w8nby7b
G2oKKTyB+u1seeWSsGvZdgTPOxlATJVG7SjGmPZb+XBnzmbpA1apm03r8gRoQXBvAVJog/6tsfS9
xHhhv7w35eZpI8ALXJhwJNFNoySaHYQehSOQ64jkPfeAReilyGLY7i+wJDoYsz1Q+zTKBWjI5g5o
9KqeRnt7s/N+xPUItd5Iy/4Yw+ie40MS4lLc1Wq9/XAJLZCy+34mldAu8hfcGI7S6dsvyLZWJGab
2l3sefpIWUeVzFFHMCGqtB2M4CDXjxWgLcA12BDw23XZKMlN+2TNsEoieKij7pbbTAhr6GoATVSv
di31xvhWiZLW19GuHghsFweZpEKHnB0Xyb1blOjlxh+C0bWbUdze5fgXE2dx3y8n1F8b1st6UBcH
msuyHK+CXSQ7hUc4H/J9WivGQmrO1WkUdYjVixZITeK8Rlw46J3vQsljrhhf8ZojxA9EgL2P230M
FGUF4RrwShXORUkzLHZOtgd+HBU4jy44yG79w5krblm8CP5q/mpVSYBkiS94o0q2ZKzkZ6rB7hL8
BhtquLCbKmA28QPZAWh4Ed7M5apUrMHVvfaSWm7/OJu6b8C5K9AXsOYCO+JHoXkYdevTSoSOHymc
1UcFySUvj1KHaV/5cOvEipvBCmU+PY8JvgyaoVi38uLiTgvBAobekKdwByqj8P5OZNfz58EyXYEm
kVm93iBAWXT1SxQO21Xf0Xo1jFf8yQ2kJNVRUSOQ6v6dexgjiZAV0fa5+TvrSpLo3xOObF1WY6qU
LlQokORsyWjHUgSr1qxBTsGBTMw6vJtE+HG9wQ4tCrp9SDuH4Ancqj3NFZssfvm+plLXEfFn881K
3z6Z5zdfM9byQHkyrVLZZfiKcoM8ROswIDl0uz4+pyXxCSa+9xF+f5jkQDxrJPgUb5uEX3j1vpdI
SCYj7eZetEqiowxzzPVuMT64MYXYzpm4A7COexjehdkJCYYPRF/hXsRAMDNhi8tAWlqDL8QE+oeW
HwburUv/VAGnDpFcGxMBf+WYoErQIOE8bk6/ydnX236PHzYKBL/T9lckitB5zz8sU+IAO5lYYxvY
SpMP+J1Tvaf2BJ7s8rxKj2E11ec4SmWMtXZp4F3juQKjXpHy2kjJfJ8P3IA/dHwapLVkpu7yjF2Y
n7uF+kYgDGrE5d9r7ZM1xBy7HkIdvy/5cKr6lgvHieM+xjQc9qtkuSpksnWqqKGq2qKt/jiRFAg5
fR0oQNeQm8w3uGS4ku75gtJwnxf5pQ6sZMf/irn+pIasCMwmsc8sE4RypCwXQ6+VOZ7qHnOwrL3u
BcBtJ8PvpUS2964w6Mt9T7TrSWDSwRYpLlrEbyKIfY4Z7ogSIWy1UcyoaN9kzpcbHHLjmwC/FL1F
lnbwIMgabAc19miys8JcYpDJpeiVhGkDlrFvbBeUZcAA9tkUDL2EGYKQ4w8ZpUm/XOywJMYOUhXB
IPGWV822HB+BpUjwW4ZR2p9EcfzmhQer+HkNXyFh/qc2zmGoi+rMZ1gYyxZS1ceP5yEbHpbO8b++
Xbo8hVPIFbZrMQ7UATKq2UOoZLiD9CfU+b0cE2hAkBfrktGhlSgcLgyzPAT3FTH8VOsO70NFjbHw
sx30G4lKP1OPgWhs3t+9VvxzDLpcYYs4IXclHQoZfZAsKTUAqeeOLrLIXs7IAAQybcjMWSOxEggo
lRWBdHdlVeLlr1Z7FhZ0K8rWz/K84P5OhEcqmeWKF3pP4Z0k7A6W2IScBOUfqrfXWk4opJa7k7Gl
T1Wzv5yZZlqgM91KfP2ma8IiIpGvIgZXbGrJUaVZlqnLCaT/IWw/elpSal18/k8VNabq2ZrNEXr9
Joyp5lxHuncXmYm4mdt5lKj/2jPq5KonMwROmODapZhGc4GHb0TZJkML1+bqL5RpfDMKfRqaM4FA
DbhFblIxegGBNSLGsnV+9mloS+AKC83J3PvSSOXWPTpIjFoJJ9WmexnRTWX0gcNjSo14vHG2lDi3
CP/PHY3+KweGGO7tkxHu3CuVlsUuGR6gSPZ/gnyQnzfb+xgKc9zDgrmN92kFbjGe0DD2toiQqLNM
NbULrxQvxPuRD745pbph3CpNU2vrbAUnvKyiemEsi5NLWCrxkJY59NeWSJoJlNws4RmBnA/fUSMq
Rf/oqbux4AXFUXIJfyfds50HT4WEbdVJ2ORGLHc8ePuSWcj+S6c60gc7SlZRCsfX1DxcYeW/PhQk
s7lW0K6qUEokfenM35+YyAEiCzcvVCRkY/x8ulaGV6UO3LxMrxSnqPDGPz0wO1oDrBcNKmdXI1gz
Y4Bpv76QcQNGlNsydaPPczXGMsk187ouyyOY5vXbw+2ZOejPCOhkZ8XR8HEblCm3Mal1ASQo+ni8
EXUAZE6/QTnUPOr3Hy/ulMFnlyX8vPyUVwdJuv7k6pzdgdsBV7DqiGtmgLBgVLsXxt7q1NdLdAbm
k1sGxS1cLbLHHBBCqpJRVGQC2JEPrsSWQpNXQzEcerBLMj5GqlejQZLNmQqovOug2PSxvTdflqVy
dW6YuXp3bhMFc4j1j30ahuTImRqSXLsgpFS9XphU9TngxOBZ2Z5ouAQZxitwO1w6cv1Fj38YDcU7
r+AclOulPwetM0KGmqL+80iNyEb1o0IYFT9yqBi/fQOf/J9nuTelSs+/798FvotLraD9msV8jsiE
Bz0ppZsR3am9jlhl/uBEy2XnOjrJS2UlT+PBzMGUFMytXvmFVYj15vi0SLeFLw5wmVw9AfZJrVFw
YycvVPgRA6aPgLXryUfpbA57GwFqrge9a26ATSEKo71NrjW5gDakym4qdFddZrLQ/hUgXUct+tsU
h76YaKETjcTezByHsuqze1brdbXT1TcPAT/xI/TaKvUitUirjoLj5AGNkuvabbG5OkpLuNmWFZmU
tdo+Gjz2Wli3+FfdCamk8xxlvuVz/JSAJA7W2UbTpqmUmPP+8dZ9B2sQyl8eJihwWue1qd/OVDY5
FFDFzAPa3BkNDMeatVRWtVIDXUmNgZvSa167ZKwnbUuiPhGFii0ZdKNjFSM23yl/TBw0Cze1O1ow
77i1tq8T20tBNVdG/P4y+fmjm+dYXtxZGn0uB8iv9tQsrU9AuJmfBuoQAGaYIzGcxHn0qlDpiAun
y3srC02H7vKpDoxf4Q4TFPgo2nm5smINe7/BOgoY1NvpOoUSdDzRpKDwilFrWaIOFALfYmA5tTv+
Kegn0e9yVALatqVeHgQwG0NDa5Uhk+cmlRDTyN+mKgTnxgC2dTbQweuV+xQzAd01DSh6QXtPO4ez
HCojDJ14ZSfCNsSCHc/VllgSm6sT0S/DqhfTb2daUoGE5pFSBtT0Z3m7lsv1yy7ciOuSD0B0Cbjo
BlRjTRBE9tskfy7qDiLeiGce7u1tEf8wxHZ2Fcr6WIifXNn4VL+sdofZteUMfuK4Fklufzbw2I6z
nohOqO6IWnDN67D54QNjDG3CtjjQ66H13iESSqzrAUYLDV/fo8K7Eln4KU0UshStecc92Hnz+VYn
QQwTEBInKgj8nsd+NM1EF0ghLsy9PWFJ5tlbstIugOWUrRNQOcXm398xQsmC6kIbkh2nZUEl4Apx
1DX99Qq21eNjVdmeHZkYs4VGZm7MLZFEgpFw8Q4lFycP1kPNWpB9Yzn9AU8DPJ9YGj3lsbTdjbSa
uY8CIX9Z6sUFwjPxP9DVVWRFwB4mH4JHnT5ouwWRRHuYzMhSWWsNUn3ieDuneoTG77FQ8QJsVvqU
1G5nmmPsWdeTA38n+jY3NucHntA9nA0jCo7sudZt/eEf/BgOUKftWgHlmpJsNEIlLuoiSQlY8+K3
cSOdBSVzlPgeVTjEPTa9XqhvRafiEbZDAFW5YHIexYnt8D5vZPjj1dP+uzMc1lNrRKhUN4wrG2hW
3BqFv4TdbmTSNgHdtH4opDtYgm5KU3l3ROcOYYbMpBk7slnl591YKUXWypTndNCk8neIW9WL4Xom
MHJv59E25YHOsc3mRdCuB7aZuBwMFDgWqZTl2H+esPZ/6hK/nuMXsgHYkA6ukB8moeVsmnmZiuZp
7uQwFnehy/fiAGDnb4mzURD6MNW8K3yT3DO+mCg3C6xvf8yzhhCao2Q+8VRW1di0ruKo6zI0ZFdb
47+Bbeqj0MbtpW6sSaZLpUSRYMH9LlBZ+IszVIw56OWNi+l4JathY/hEv6OSARgbw8YCpAbBnkTt
FdmPtxKIiImmWqnUDyRdArBOBP8E4XrU8LUxKv7voHQz02mNNd+YFFNG4lRhc6edVrXMYDL16weg
bB+Wpp/Oc5wvRKj6rKiFt+ruHmFORxy/wKb6zwR4NoN2o5SY7cEUdeNADpa9VE1zodb7C0+N8DW7
MupVWbCttjPwPh5eUqBBBcRJ8SpIdnewIqVteBCzgFNzmcWs2Rx86GWJp3l/CRfvoTZ1uI4rClzS
0NgAXPvheE4rQXhLJxMcMOo1NvoV8oS9Jztcu9ZySHLhUxaSIauNWVVZpYzftMmT8ZKT/gR/mrLk
rNmMnLLMNQSBTjuvpNgbiskv+VeoabB5wiwcTKbRTkxATih7DQUX0NpXvLIgYTpQTnw/46qDnV+S
Rh8QI4SYVhxzmB1sBODtO3mlBB7Iybes9MI2pgyeE62PTZMzS8d09wedEHYeN84/OqqmOGA6MKEM
awgrDJ/N8KMrxpvXjDbU9vpIYcPU8YcoIJtZgyih0F4JdsX5LVuqs1PuAm2Y6WRWFVy6JWqcxJQ+
iRe/z5/6rZRgbq9h7ENzw7SKmWJzlq04uGEKmPp9wEovHYFN9/uOVx+4+wKRbphn4V+PWZak2YeK
KdUCybkc/NVk0y/iG/AtgDIr7/16he2SRUiylR5e6C0MeSUcQFV/8MmU52XusBIszODtVa58yQrQ
OZAtL+LBHcsKm6YYHX5JQQTKAbRB2fZV3SNNKKqVfnt0vYob2Nr2xS6Um+twtLtsft2OChLc/7mI
74MXvYjVCehaPlzciG7ujFewkJuF325xN/RufuWIXSmAJdp7OWPr1pXcyV+m3GvJjxLrV5Lb/2zT
WixKRTtK0SPrkm4sRU9XSc7o87yMpt+xsVT3jT9+rAvkIsA4X/DHzEQsyAbCxwHOJ5F8L5RlrnvD
P9lbQLxovLq9c2djy5IXWhmXXFuLxgKwGwoL6rdiXhbnpWX6iWwtW/TzfbBpWAkveTTpb9+nEVVc
kB3DvILEQZBkr5R1siQ77NOllSgjQW8SIKuZorXkeAmw1uUFJIdvLcbhhTCyzmMr/+F0ts+SKjaM
yNdmwCRjkK37xXzHgoWPW0fGzo3fErAfONUTWZHLMDIXo0kyF7eVgnVdWwtTFhNzq0lsD5LzO6NL
FPOBIFDEIxK3vyp/V3SpJtscgh6eAbzCy+lKcucktwzMlX6nCscwtUG+GKATzJepzi2rYzB70mCl
kpt44RAuS5rEkHfbSJnzw7aaVvLkmCEBw4TXAw8N7nL9t38CXr5NOJr2Hj8KJJHDEQULRGHZ4Q7n
Gl5StVeGVLlHU2pB5GvMnG3kYQ/6zL4DIPUIa5qP+L7zg/9vP/e3SqHg3+0LlqCOqKZJsZgcs4IV
+xej5HvUC7C2ryo6rlMvVSq9rgptvMUUA4SPBAO4eIn0VxVvwla1/pPkJqqDd4JhmYFLEcY3W6nm
XyrCjy+iEWmXwXTvOx3Mn6gBHkZnHGixU7H1UavdRq9Z5m3/ll1NUeGd+Q0BZUJBmR11koSf4Yle
kbCo6x0SdcY8oWd1hLXs9LAwkQI+JcfjC+GVNLs5kIy5IE2IZlYAJoltvdj2nPgRpEXbNBJJUsuA
41oL6YWenp9PzsOz6GF0/U0CzVS4wW3AaUIKea8AUZVdnUq4GHq1rxGycNsOAY9DiA6vXMv6PXlV
mCbpTWH1Rg9VsfmXvofadhzwCsHU0wwEjetI2rPQo7w0bYGPU9N+jagmztkrioyunBxPjKuYEOAk
f2m54pHc4ALV3w18Yc9YDYvZxlVO2M8lM4GT0dzqgO87DFvdWRpSxMs7CdJq5aD6+7Y6ILaM7dd7
Y+g2AFu+R+GVn5W1jR+j2M1In2LfKsw4pX6FVnQTHZtndgsgNWtdqVDq70uQS35ff+kviCZqtunH
C0rudGJflbEbeFXwMOeez5q+ZzVR56QkFeDytR8v7QxVL9wvBHm7VeqrUk+ari9whUeOVnfU55D1
Lev4gZcsxc9gM0Zp7wcEOO872VqbbDgsrcMrUar6znVdY+1hg7fx1Mjxj8b4MWEo4tIsMcsluYum
L/7F5R7QEpBaj7rI2PqH1AjmMGqiqC4CRnCcf0AddzrKwTraODY3zjISjr8CnzSu41LP9skwMy8u
/VqOdzPjWIg9HU0IZeybdV7oGMcYDi4DJkQ0YrlVvSqo5Ct8MYwaWeTZn3J3tWisX4ZY9p84v0r5
fM6ZMxHHmmTJ1go9k4YTIkddW3wLfdDdvX/5XazTAT6kBlSP6Z2yfO77iwRFU3KOml0hYcSf1VOM
UGpzHSAtcxVGd93cg2mEFqLmv85jbGdnqAfg4rKEsnjaAGSwluY4dACnlOs92hW82LambMGJmMX9
IO8pkNkyzXczBIQ+iXa5FLRKMadspTwlTJJEQy3Z/BaRI3m8yIJycAF/dCkzTc7iXuY7SPHSUSs1
KSKoIin1nLQrsSoplrUMG+iZmYS4EFz8Tp/fxgqBDq3cBZL4oljylU6im8zi0V7h6GAxNcvHfyEP
jzas4mUrgE33wN55EzJo081ycfGoqArWrylCiIW+IV1RVFXMayWTRMstLj7Iu9TwhQQkYCr9xgV+
C1D4L8NIT/fw7+zjVLMPJ1ZUd7kcFBPMCW6Hs0cTe8XjniR9ALmSZ41gu8BSyGwQgi3jSgiDSdAL
Ny6+2d5Qk5hOuU8jPqHNEn7f5gCZZPA2qxc1wZddhjMWtS8AJ7LU2zurpDBcIXhrvFHUZYB8bIsD
9JwbiUMQZ7+tB+Jc+G6aa57+jSUXxFDhBYwr0GF4zJdVQtt0zMbq1ZGe9vjRFlkTIM2BiWhTM1Qm
8M0noa6MFFtchnmacSsWpDG/iMc3mMUNUZlW9s7X9CoHt7V2VTC0fDEqSTyC/WK/p59MpadxaHP4
uuJfn0NGYM1F9v/T2Rr9GlYsD7ka0blF4SquYgG7edNCJI9aaaTYEp3BKA0YdBnTWBHDLfRc6CLR
w+23w+1hAWawIuwAMHgFtE7cEW1SXc37yDnOzl5a3fzs7ErRc5hx3XhMm8jxXvulExd2od9z+3vg
4gnc2H5GD7DVwEFNs6BtIABIXuBY6bzAWhOYYPFrw1Euyi/6S7F2fvWT5z4EzDWTQntZyFCS3/s3
gqXJxZ4kmSEKc6NXoBFOmUKkcNn5AMfmgfizYjULrn1RROWjaIgYyP1wiZpR2HiM6A/YLM7bK9+2
xyq8VaGVxrSckGKA/9b7kdLKJVAOU4i1hkdUoBxkVIGhH8LtTZ/rDMYjDpON9cOg8TNGemWyxaoq
TJ81DTkp+eMzD23CoeBvc3TxKu0juMczEQK5PUi8A9O7oU8rtcp92Y7NuIrJWVTEerIb5pi7j/pE
XHCyryI3xvSGUt9EwDpTsdOXEF2RM9cnER1abPChBYsvHgfA2T7DU4Yt9AUeravWu8o/Qd9HdSZ7
lDfgOIXr6pqAZ59mumvwdwbgvI3LNwB8G8JVNFD8d2Vr/l0hpTunknhsHab17Y0wdLNaLRRISs/C
oTssZAs1Ni6KNXDpQirRNSH6dWvFxZqqTvZ4J0s+EYYaomhwoRFZilhhF//LK839KU4jPrkVGLU+
JxbEfqzrKpCbFO3+mhAtdX+zN2pHymzhh6VdHdSD4pD9OybXk4e/Ok9Qb27zBSjIxTIuR286tqTO
4JElVIsi1/L17f3Pg+LsqvE0ph/pDnI5RetU5pZogaWMk9aSLXqle8NdBP8vfkpMzyVQWkp7gZRI
MODRHVjxImklpyUJHbWwFt61YsEiiDKyQ6475O3Kurfh3XHDjjUUsJSE4x/RkmEkObkUQs9syUxW
+CVYxcS0m2k46zLpQVv8dvh2D8jnjLXPqAo9j5pLv760RnV/3x4yG/rJ/cTXq5/G9jCdXNkXazRB
1VsVr7rRHjBUt+HFyIKVTmnRSCdAfrjzsIumKgtaitD7R+f8zKHXACU+P8joWuF6Fom965IYye9Y
qUTdwSvm+RSV1aWEdGu3pVgSAiFNjjyZPDmYAioBtikg6Q7x6FO5LdIMDc+3ApkGyXAMVviqDVNu
uRpL6BdfIBbd1QTDiFFCOuZHOW3JVvUGta262mrsHwnJRqgQ09944+VAn/F5VtrCG4p+c47T/+nj
xRN+NOoaLykhpnVvqaJuVlXtYjrhUHzwpXwR5akXpSSByKFXoydEWehJerubhTi3FDkbo8/Dr7s9
AQZmjIb08kzjorii+STgyDK5UB3o1bdT5LCnE3oDRCv1Tu7ly11jwYLGTpbbtafPVAO2IrCujZey
XdwCZeVl+staeMlSAp9tOn+P7ziKMd8taDPxFkfkePvcVGRNZkIiO9QNKq4zt6+sdskIoq5jQBh5
DXK0GOGwAQTF75pp1LnoELEfcR820eyaqYDHqLmsATcP8tg7OpDx03ttU04bMosdrJ7fkHjpAkO1
z6S+YSYghDqq5AD+kkeKZyGVqfW7GnSCEqfyq0pIQWe6EHPehH29OIH+NFTNrEYagzxIVfM3KAm1
mdUumPFQo/0eZb1OIaq9oSTPUA1kHANfHt57iaZ21rgSQjES241GkG9zYWIGBwr8m3oKG1f0C//9
FXDBPM7FgF/5+retfLIwLxpaepPHOjx03wX5wWwWn1qos0gslBA7L2JTzmhPvCAMX+7nUXVGkujL
cs/33Kml5dLyy/8VEghpi/aLWyFHE92cfE1ZAJbfDf9ggIhOLRinF9JoplWQO3LvyrHwTsjFjr/K
N2g8rL+k2zgIZDoRrgydnCpehubyPwj94+CJACatE3b8oK7TfHx9/YMb/iq8r5N23oz5azcZu8/d
Kx+RGB5FWTVnONwhaxmKARUTQaBl6gH3k2n7Wwa1YWiNi+xdCeLMObxeC6ghPLqXdBectj+mmXHg
cupNTX8LVm0VbEYD46zg0JKM6LDiePszsNShouVXONH8D1V2jwT+tixBzKuNwcgNSOirhYQLbYrk
bLkERcOTXi0jyiKQLiyazYs89joQXtDkY+MdLiYEPbGIEWFJ5BJBklVJsQVD4UG6uOSLcX9l1eHf
8Pe65Yuvg0gbWjJoY9jBYjXFld+vaB5zKShnuh+b2K7vst0AzoJ4dou2ns68vpFvYBhu+fH8Ouka
PPAjFFAas+BoysjnIF8EvsSYvG7HuJgTim7VFqCSbW1L3cI/MIsm0Rc9s5j2E2xL5l+47txnE+NU
SdtCtWXVnIQPU/RV8v5oTlagw4tPu8j39R13UHBEOMHIeQjXyEEtozTWXwGR1QbDaAD31u+ID8nR
xlQG81sZy4hsaZu+N51VO+TUOvJdwVHzNfa/VzejEGFcZpi9/N3/srh85om0we7RqgqLb4yPSktC
9cRlXhZV/27nmiKmnBHcDoEMAF3e3hlvv8u3SE+xCPniX7ujHKPVPnIDCG2MLTtb/h8cAPbDTccw
m9WwBtnnIDdDKF7WCAOm09urtnRXyCzvnbSxB9bNFX1GABsteZVmAjA9K4sCfaKP3/RnZFQcUCSJ
NFPo8hw8M0cNEW1hwxf4f0g5yiBhVmUfvzV4oPoA4EdeFAhIMTORistkCtYVzwz1KOznFbxEe3ua
INayOupaMuWHvPqAZOqEgL1paDQajcfeFazIFKzgN2Y9NIzoD1lQAwuk6fe82nhZUBPhZgv3Z6e5
Rs+g6Rx/f8E8gCbsNAGnWxyHOzVtA2VSo6w561voVkaNnQBnlP93nSaqe2zUmv4/PLs+DFMhcwjb
8MDiMO5eg5wKLiUsbsmMQa9Qq0UMT6RdL7i4ogKxUm+U6mGp8IoESAeHG2jeYxPLX/IJyylMzLRN
yLbf1BJm/5cIoW7F0lxEur0Nf3StA7OaZaMxnEkfjjtG+LszHoDArJhftrXh3/slxMnleo2roVtX
tinpT98k7K7ZUCMq8dCyf4rmBLyV7zgFUBRHEzxzolNRBSJeXxYgKUoc/c4dhSC7SXNR6BQxCWq2
2GjthEVk8hL9XEs7P6KtLHuUz9w4wKr2i1xeGGVrReZH9gpeWPPy7UPtiOrKasSvwC2nvTKiyn79
/alnp7yDb4AK9AdiOIGta3lJprOBUUXkq6/APrczXbcx3qkQYTkW89EgPRFtwM8c8SoJ3zBHCtph
tEAMXEwuAVflCBg+Ckn8ONx12lyHgviUIMEJBXc2cyO/CZ/Onqz7dj3SAliuSZqeebYq8vm4D1sj
Aog0wU9ZvvvRoHv94Bk7n54qlGY2/aHTgE/7fJPnMMLc4CpRPbMBo1amzYttTuzspzCFNUgmx3+d
49S+D6c+Bc0EkrrGRtrnf9Hna2Hy0RMr7dNJZaAyNFELm0SXZSKgYxWUXmSo2yz/Am+XZl8BN+3N
3/RllpuZV/K591X6UhJ1DlLW53h3rnHTO83QhSsmDkSGhlhH1bZOfFpHLBm9aEgFQXJI9g6EJQlP
gCmv67UK09EjDluWZMTNhqTbhzbttcIRtQPmmRB8gYUiaRq0hpq/L3JkDEATYIlBLeYA1ubtx8IR
cKfZwMRm9zxGtTbDdU9uni7sjlHbM4yVdwc6h1yUAkZAEKyusC1Bg+cv0h5/Mzyoysit68rkO/ln
hlUBMoTo1Ke3DnafPNXUFnmV/let00ovYRG96c2wrA2YWHycLDOr5wtg8+v7qVcE7rKZnddSDwuJ
kYzHRzmaIe4ln/uY35wdQ8Q8kKkli6Rk4GmRosnPDO0BsIb+q+ZBPG55AqYmZP5/ts7J2TY9Yw8p
g/42l9pB6RvACZCSX9WDsMSCq9cGjs7jcBN0P27cqlk11tpJiXcwiEURFbw2EquzzUoVkayNQZda
HQyaFIsoQPoUZwcP7cjOGKHFdnNFEE1M7yUo5iqRXH6Amah7ZUJcHFY/rTr8NymnPdqWCUeLfoP1
gERmrW7STeH6vsbfFnhI4bCzC5cw6OEi6vgBq7hUL1OmPAZqKceAdfpaIC6w8ha1HnRps4VpTZ7V
h0CpgZPSzbj0s/L/FU0FsjgWmi3vCfwrirgugxIVHkOQuuA2hvnRf0akbzr5MB/jdaH/DqtwPDli
jB7/YGd2tKT7DYKf4l5WBYJr6/Lvj4FurKEAqiJ4q1z/lfGxhBVMnGZCfkdADYbgatzBu0JmhyqT
NBq2+yJtXaMyRqdOEgQhCO6RgVJVAvTjLIBNG7Uypy0ve6Gd2J41zDfq1Dhqsn6DZzwXIYpzdYMN
BD4EwDUqUG6H27wU7SjTWfVilrGiLbG10WFcvnT7VB/XAiX5QOlEgfHmtbcl6nc6I1fPqZzfCtSw
X8RnXoW9fyFJEyTMNzHDE5kfrIPuSi3F7BHLd/dCwPj79JI+GJLlk7IRDLBz55nIzQkppI2E4WPD
CbblsWrK3i5+KgaSCiyCDbqhqtkna+QCVChS49QmF/DrbPWukZ1enkfxQDfD/Gi1hNKm/jSG70Iz
GjNDNRYf559PgMvyO2+l3BeVYjDIQRZvx8u05hTyaRu/ZK7P70Nkd44+4VN9sK4CfI6D6ZfSt42A
Mwc7z8pwHHu5PXCyK1zm2MA6/iHJkdQsjb3AQfeJZuvnC1MK2s1UvEd1tKWuwxhL8X/il10+0H6P
JvfMuEoWkWotzqZeHWdzSnGYfZr6BHxxBF7RKvwdFaVsLXJEGgfiqd1p79I7pu2FA1QDtnNfqy+b
I+2eDEwf227CUYgjcp7ZJsucZYJiqeOGEA6BIc5e3ZjZL3guNbevijHZm0pj11P2C/GJWUC/+tbQ
GZUPlpbf9eEmBwtDA6G/JckxVaG9ZT85tZZYMefRlqjeSLg7FhLf64be59a+ld3aia1JwuyuU7by
dMdB9vM0OPIWqBDg+C/IyVF5mx58vIfY6Qhhit93nLA9AUObe7W8yHULB2H74qb3U76XmcHX4XzZ
uatykx+Zah+7CRd5PXVmGE12aGvkzw6D7JQSuX8AiUtceFv3L0PevmMMqSzKid5+na8wTUuvTIH3
51bIXtclflMqbbiVbmxwRSKSVbgDjBhcwNgWN4zSeyTJOmwjH92VQexfOO2hEx05IpQ5n94vvDtk
pskkkf2+eADwNyTrRlda9pPjzyFZRd0iwKgFYvQwrPxPqN/0aaQKuMTL/+u1KQnGy1AzEqwVjxC5
zgZ8Ardyz4C6el8jwrxdnSLEb1U3fNrJoo4UmglWa4gZyzIiELKkA6wJGMmZ75qxX3Ne5lZRfBr8
C6EIzjEuSiBiFZ3s5wQLj7ZNKr4Puby2fAQzFK0xRGob6ZAhXusPyLRkHvQKoTF4dYM1fkP+sMsp
FMOO6VYHCnHtBLWc35x9IUh7cJdKe1STidE2kDg65eJVWyOit2efj2tcEU+Gxycwbqn58hoh7efC
NHvdbXisiqk9Yy8NqpjtUOu7JR/G1if0btsVepD54aNgym6YfIQUTTZnQcH/igK9AVPdDvATw4PA
YPEt71nZhQYSz6fPY5nHfHRdBYAnoIWXFs63Sxv4dvnfWdU+AVggcYS/iZl3LvnlY1MJ8oTPHQKm
bU5gUTU3UnSf3k2Li3A0a/5J8Tv3ZM7H9xFt4GapaXVNXIjnejfjUaa7X+LPYRRLtTEWH8yNcJyU
TMLE3gSWJt1oZBmFRd8ZPRiZPib9Jsop8fZyxTfUsXHpGCLSUnkh+TcvN4Rh190MGTdNPaK9O/RZ
UI1t4AhwX2oPWy6keS27imy2EKY0ZO6s0Xeb3TztolqKLEzZgWr6+deb7zae8/pIwx/FXVAldXA9
9LTzCmSdaGAHlNVsIpNar/b4xM1pgq4JFNC5EZLMlwjB23sgHCBeTZPg+ayNChLMsfcQG4+6Ht/P
HJ2oDOzvRGbCioJR1Qmu+qH2jrdiSkNwkj6Qn/QSlyAxWgou0tDils7VzUiX3BeKtqrPyU4t1oKS
tlV9dZEJMvccgojgeGq3dUjNHIiDgssklnjAbS4Dag2VdZz3CCEw2MLSAR/kmvVBc3mjDQ5GvOt8
yU6jH33e+qUt0uJBlXltNnaS4DPO0tmp4hjkfJB9gkiVBqGkE3l0i1fNRnN0zjqknC6LUxNSXFbL
aYTsZpctsxT3MuwCphkbyjLxriGuz8I6yubmV2CZkDAPJEu+7QlCDrrkkPoFSlylDsyUiPROr6eU
ojZ47cBAY0VWsjns9r9gM+hqp0qIZvKz+2ANknRu/KGr5YczB4klocMz4nz1jo+pXYmKZHajZSy8
QNUrEoQDC7a9UHwFjrscSAMd1VLZkQcysR6fPdAyQ9lDtFeyL+LfG1GoDdSfl+APxYkwatcca3pk
pw8UnW23CRxVOMHV4+jnIZk+zXCAeLFVo0tFwBgFE/t2JXTBVH0PDU/peOSgnAA3Z6TEGntiAA3h
i38hteUrpb50/iwscdY+/PwonxpfxR9NUCEjI9QaZ3vjcfSRdrMHRCvg7YfhSFEaCHRRCFouNHxx
DFPjIT8K3zGGuINAiDu7c3JWPV8g9eSHj0D5GkygAOeIEVg2ZihJlPbSXyE0/GihC0j/jDlW3g1Z
SbBY9IFqNJd19sc+MiSLTNwvtGBpb/HKBuxmquza4+Ugwv28qs/06hQhjiI4pwx0lRdv2L9VO0Bw
cmUCKKirno71CgwEWJRg+v+5d/3rzpy2JBpG/fsJcsqj0IWMuECo4epEi4wVbx6hBD1wudS2T7cK
wsBvRFrfN0USZ3Z37e9sXdwcYmSGICFQ4bqqY3/wjOTPSiF4i2cGh8vFm6JTe/o6HvNj+lDH2prL
jv2oyli3J9g4i8jRxXPWvlTVp4SXNcDBZqke41RNikDP7hchSRmiusNzlgPBasl3cBa4zGmO1tbD
y4uzgReBC812JfHco51wMl/p0g5hX2fZQrUS3HA8GQuhB1/MCug67y//Grgj+vnnib8Kamg7UcRx
vCywOcFCpDp596VpquBTtBuWm4sAlXinmtzjt6EZ7SHHPt8/CBtbialdZf1QjVYFqsxzqchkKwgV
awL55O4peIk0wGrXnRg0oikvK0liyNQArv3Az7gyzrlIy4T9EXqNUnVXLkl0O/f1Obp7cDTeYqks
VQLeANLnA1W/+O1h7y12rTyT/hJgO1lDNo8koZl+lzxLtqOTj+49vHaajPG16hyKkuntzhYLfYf9
Yj5vgmC0CyrgCeoxvDD7nwJrPBS0e4QjsvYo35/ZJeQDZpZNA7oT/epKiHMCrxom0mSlZl34+c3b
n2/QQ/ooojQIsNxxxPLAKnzj+9DRUhQYHllGshy5EDF51+dF4qQwkK+IUt/oUVpWnIIYHTFMfk58
MMS9uqpWvdrigrS39ZsS3IJN74kYb4uBZNP/cwRUFvcbJzGZYjHnwKTj48jsa6ZEKvxcHM+EfrYk
tf1Bak+a6M6O51IN9hBulhlhxd9Oea72LQjLx4DmgeNa6AS0saaWPNhU82hsoNTYIzSeVIaSaVED
tSi1rMd5tttS7YKlxR+ne0v+AhdFpyDROHwlO7wLpoC3S3dNkb0Ysde+34OMLNIKoyWu+O9SROof
xVeqOJsphyeklJ1hdvl/ha8dEFaLtk4vy15RAch/8w9cYATgfsRL1WhFWbasZKEz+2S06qGv3ISq
kphMDFeQiAsP2DnNoko6hMdFKWkQ7OqW6G5hSPqgt38Iyqorf2S0kJuYIzTCsZph2ANFsr8KZLT0
sp1K723TSj/YQLQf/EIZuTwrsZaEexH8BDKhfp9286MLbUO44qik0zJPpFrGQJf5IEWdOFSJCLdR
Z6wv4hdLZIELc+RSxoV9jSwu7zXpOj8nhMX0XnJHidjf9jiHESE5Gyg5C55ZvPN7HN0vFWDwB0u7
l8zV4Pj/osGX/J3TPLHujW/gD7Brhb89188VicQB6ck84YI5uKSZnMt6a919WDWGndQOHDM02ae7
xWo9g0m/idlkiYCH0k7DJfxNclI3T0aYZFzr9QEW51NSS/s4goocpPjlnqoWjABmmSaKK0x5aDNZ
eTg37uODt9O8tF+QMn8KMpELKgKFM8T7J0bNMMm+bGuNVGS6Y2fD196a5XRc0YVcgBnnWBHQNfL2
mL+fPKyPbAcUz/Q6slX74wBygjIVsh18Za56jJnX3+tTbEXvWmpJZRWmO4ariTdhyLg4EPc1UUoJ
GUu1WnCy9WRajn1CK0sthWUtcxmqGN4wAOl8s4btwFFFBpYJYnoGcPTcIiSwzqjtrNpE/znijChX
1bn3ZO7UFQFnQj1EBiUvtCwJ5xML8sSPkI28mWevIDWk8Q7CXhL3Oor5GiDFrGajLVjL8JCPY+yQ
agYrA8g7+EkzN2NsanqrTT1zM+XfGk3USRX5aGwCQnZ2Q5+r9PmJCyla8bQ5PJAObhJ6LdEaoCvR
oHt7z7jm3g2WCqalhkAu+ExC8Sc7ZwGHY2+7cC/pmHqN4fOjCdoILDVY2J0YMHbKmjIMopZC+b4Z
3L+w5YFk0NKQAh2lxZ2TZPQz/vr1yKoimopuvYc4pSUBagrKtJvCD+1LsZJQAea5mX22YrSplUmf
9Ku1uMUY50TC/8Peeoqd/dpaLp1iqKbwoDPc4KmLkTNLnxxaKZskMxeIewEPv04KGfxbrUhddSVQ
nULBiwTknpHtc+WCKHBTyjf47jwRiwWx0he/BgM4hFautcp2txvVF3mw4+63Wdx6iAxekqzT7FCV
IDSJzL+5E4XJDGUmdyPL+Yay/738OWd9dOsRthuIWDtJ4nliA92U9BFbe2A6MFQUUhB9sAbbdA8P
J2xGT2D3MI1N/xV1DfMJVO5ntfehFVNT+JtgkefAmv/AMeyE9xE0xtFaFWyYBSWdQKuWOMqbmkuh
xZWMgdrQEEjMb8Sl3ldKXCuYaPD/tGADDytOCilqsy9yDlLtIZAzmTOKYh/DnTUYjAwYcqO9tIOL
0zWTfZwv6CSUA6P9SoKuwZO5/86JrA8hy0fM1PwcXyo4gyvRl+YZj5UYSnXsRL+OIp2bP3z4B053
q6jlrDyR4JyVRes+6my1gQnTZQCXcfGgC49n/xEaX8+2pCv354icEPH06fu30xR0m/o8kkXc8+3A
MtRZvJYts7o6fGiMPvF3bw+JIOlATOHAJReHiX0jxUGaNlD43bLRYz+2Ya50boqTrHshrDw8yu7k
GeEDkrjVrRfbRqh6U6URKBQZg76bP38N9TehcASWIqNGSdLcrLRQvRo7GtZXOaiTGYo0Z/O5Lte+
AQIR+xrRSOMKjnBCoJo9H87Fao5Z/RN4z21zj2hYW2izsPDiYGj+2qnZd4JwHzsIS/g2kdBcQuA9
NUFurMk7/51OmuASne6aAgXMRRFwY/Du7gmxvdnqOGUKaAoSPb9Kok5VtgRrJ65Z7eco3FpKz2F/
iVCkPiak/AyFZxqOWwnRcox3cjzPhmtJ4+fVb++fN58SN/vvc7p5aqq12dis7UD9NOXM8wqtfbXm
KuGrfXQFh5BOwXWDnmNWAkJE9DCSB+rOoy0dnYxEQL/AupAGuZ5lO/wzys5BDaH4HY1iUD+63aCA
X573NrNC++pEHqDquhzZLf7IsNrMR0TUTRnjsLZ2PbyfnKv6dCUqfnk+JFkv4YwC3BXonyxJXfrZ
bXaJbG9hdIrnVsHS97HCAKYU4/FUbkPH2XvfaRn46dpbeM5yrsix0txPCwtgrj5K0V1zh0DN7fhp
eU4su7ru31puueoIDuYi2KOXkuGRWHLa8Em0XK8MkqFKi8K1gMQxRCJzBFqiPmScxqc6kY7YCdd/
S6kEK88ir0kJDQ6xaCZu3GOZ4qoftC00Zc3ITdcJWUOqoZnqSSkB8uvl+QYtz5IjG9oSum3XYPAJ
NzTYUZDXyrn4BUN9zPK5VsLjwP2pz7Nnb5HrBthIqRNlPCF7W0lmntKGFdd4aruKJzj3mt9FlVHj
SPEk02b41mcGd0FWFnmbbJ0/OC5M2r0ffNVEiVBNslEDKhhtoC39Mi4UHj5++O8gomRRDBFLX7zX
sxk+HAO4/KrjGaQjI6rRFe05uGRYa9328sgJEuKUQTkgbYjvQ9BOJuhYjWkU+9X1FwtK2U/8L8wR
VxTQ89FbjznCPO0oSxGdmRkWMLJWpRV4xM/AAtIFTwUT/yNcrARkRs/vpJJKp2DSyWCe75vuQQnZ
oo/Cq03+Xwtql6T4hzjecdRtf4VLn0eo4urh8MSB5/yZhmTyLhDoWFomS29bqavSMuf1buqT1+bU
4maJT4ZG6+Pwx0VEPtUMVd8alZ9tRTS5keV5hCW0IVi2SIygIZ1K+vVy5FGd0GGSDZvGtrL0wwCn
fgK7u9NCouyJJDWyPOvukzm7tW22vOAicuvshX9xLLvmJTjCx6CMfb8M9VtLgwJQGI+HnzCtT5ij
fNec3oQv4VMkaIiGK9V9EKI01LuN7K7zjyFsM5X4Z4bOEsIYVc51CaOPjSs7ArvWECF1oZJ02LN+
bNb+rx1i/hOEj+i7EoMGmdP6Y42GWjt+HPzrvVc/PL2+Pz8ywXPdFUY2DuuiSx5EOKUSP+Moazpe
HKlHY9i74A5GWBsEoS4mz7Cmm2D1k/K44jUGR+YJEjQ2iRDfByHk80zC6SwgiXS68ve+a/afGdxg
3RMUzxDyUZNYVE5it68qq//wQH04i3PNFWRqofpIEnKTEgtC8UGs2KQlfPLNfsMvYlxXqDcMuipc
wAcUX5cTkK96ub4RvlBFX7qcKJ4X0M6MiGrK8F90RXgpTn+u2PxgNrUjYWnPAvf6wF7DfbfpgF3Q
oEgoQIj+r2w1g3gVhAoOGBq5me6Dn/AmKGRX3CJdLmgAs7NLfBDkKq9wWw8UQwDHrdbtg59ZnY44
a4twN2heDpPQmwd3tlzAJpVGjIgI+DWOnwE/+fUR5w4t1P0364azYiyELLyLNQwOw2kJDe5Onrdk
5IPd0pNHTa6BBOLXJdVz7mS3VlRnmr7wNfAInloOsCR9VAQqWWuVmvTDbjwpMtoT0Wi1sJip0vFL
Fb5qAnmeMjlZI0gYujtSctDCLXQUwPwVKIlFB2FCGc6hIqmC+9kVSNPgLS0wEtFVQ+0+tCIYdc+8
+Fou9wf8fWu+nZS1d6C0q9+KRrIk0A4DSd/5Q7NU7OuEDHOSfbt/YZIgjYqePFC1SOrNuVQrhenW
asITqO/wY6YMkwFVLpd/IMa/oALK3s4xGwKa8AgJhcOnOB6byeQuxge8fax0EfzfVhpwE0DqZCFU
vZAiYpg8mNe9qte/lMrPi9w2gyTs6XqFOxLzEGQvZrQ3Hsvtqsjb7Tuyhk4f8r6ncqgDcNaIvUmn
a1tbxykFx0gYs91vJ4V4ofmFUw2g0lw3123VMvHmrFhuu5TpXVFDnIPE4G+IZrX6Ck2iXfL1bENT
LiOM25y02JNVPbi6C3QucraeXGuvCz5QbEX4qgubuOtC5UMUcy2/vmOBSvPhQ5wYih1z4dxtQohp
ni7teLrD3HR+FNg4TYCNuuFoWLHPfek23m4gxWCoDv7Q3z8QEVD+dU7sN1M0AqfvLj1s/N3s0L+8
EXj1Va1nuc9D+ZSMi7Z4it95VtyrVY7NtNWE4a2xwzMxqQH+qsV8iFbn+RZ0mxqb3GXQJxkl7JWt
oNZ/0/f+QPwIazcKUMu5zWVBvukCjLX7am9shigf3QxSKlVdWJGw+sTf4y0FQzA/Yf/dz/uhX1wh
MTr58R/+jDtnRS3AmAwPuoF8Rbt6DF22+nED6f7sHZuumkjAwtZqOVsGtApB65XIPSiBJdLP2suQ
L8jgPksVLB4EHZbMSjN9bpYxr1zt35dHI0Qvt3D4SwtOi0xyx4o2wgXTCI16FV6+PQspPbefJIN2
08qoA7KxzYm6ZxBR+ewjq+d/TyV++npA1IkMZ1DAxTXUkKycybFezbuR8fdeBEBTESXc2AR4MOWd
b5BbddOOgZxj2hXCLYuhvqDf7yosqcmBG8uuuw/NopyG29RTkxEL+H0WNcV1bJf3x9N9KQvjUY2D
Y8TnafEIsvc5/C+jZOIy/VRtnA/yJTQUEdHA39y6YN0vh+bRS7dlup0Jt3WzCOh+FO0NIjO5ZN/z
+qGE+f2Z+wVnqRQv9XvBUaizbGF+9D9PETCHahBLQkX+ObWS7l3HNeVroojE2OPn9oyDNvg9Oqv5
Zq5fA2tRv/TKqgo4m1BFmOsvHzXsrXZatuvxi4zyqITuErKG3gUKbXxHYjwaLBMrPPbXYowu5Rhf
ob0pAK26d7YIuwzLLrOdq0YdyEV1/q86Jcjm4wUYVV/LtYyB08rdIAvWTqA7d2wpH+MNphJ2ooew
R8260E4kzkSey+67fejq+umhtvW0sCgw+yv5A2nZ3IbZ9mUdauNKizBYcGcv9SbgTB2cEXBroimN
+jwUiDSqUuRRvZF0z8nLU0Hu6atg0PqLYRdIT/tF8FTAWqLtyAwhZwI9fbDJgW1H/kQybLbMT+gF
gBDmOt3mdBbAKj9dtmc6PERZcp9nEMQrSz+bHcoo7Les6dEajmgve5W3GtslrhHsVDy2YnJdZyKE
I7E29J6G0LTDqpOEpjuEVsB32/6IydBJdxF1IW4P9Ok8mfN/jN6R4TjBPWmdGkuMPoUGytRRZ6QU
UDhHghLPFPC8FUbWg6UsVZokXnxFUfybvaFutv0IIAXKyfgagucf0WuO8lvy/RK9YqYrF7Z6oRlW
f8qhmq3vK2MyrvWJYz7sCtzNBSS3eng8AySdwoYmN6eWwHJjQRZXVihgWBXv96X6ysrA8/iL4Igv
OfyFy4/6R4QV3FrX6wij9GjkDE6mRmGgJejxflmEa7O2LQpO8w+P6pI2MIOzwXGmk20QLjnnRFxo
V2ywC4Ainx4yXzy530cMjgDko+mIVJYMz/M133VNioxeBQtKrfMCZuMHB6H3boA7YxBXBKmHgM1l
TBjPtigIG+NRjUd0/hK4q7SzrsRU4J5E8ivaD6bHw0cRpiJCPlaS+d26KHDYekX+XI+jq9de2/8x
Wsd56GnrOUSN3cwOS51rOyaq0q4SzaV6xXC0Xxmw07AWgSUPKTwwRDcyyrT7CsskLaCKJZF08Qpl
WZSVJ8M/N/aP9/X9RFZWK0u4kPmcN1ta+T1kuLtkgKClXQbDOVW0MJqAKilK6XC3S3dFviH2Y3KN
tBdnt9Dj3u964NI/KchGHTTVyhvcCfhxG5viCz6UQexWSFzLxApXP4LYjXAsb3omHu5LXLHvYjR9
faTV/NxSd/PAGtylWIX39jfKImWchGb+3maLp6PanZ8vSLJYB03r6Q+DRloQAvz8sC10D/rhaLdn
KkmuuL6Vldl7+UXQF1z/J4ERqjb/Zn+iWtJxpMypG1fbZ4f1beFoo42PU4TEKO7r+EATwllw6hDm
UNlWtHbp5BAR2QBMBiGyBr5uaAkodT/oBXRxf05SfsnsGXrcdQgu8/Phce5iygKoPTg8tbVGKgWS
WbtKZtJ5vF7fprGlj3k0+XtLXJG3Eiu/Fh2IckCVmRunpD0GVwwjFeN/qbitfMq/6J883X5AFyud
4yQFveOJ/7jNLgtxikMkFUet61x6ycAhc0EVbuFG1nva2Iovope0dHlyoaroIqF67vYWeFQxSWRZ
oHpKpIVJBnaD8V3OCmZCxgQxLAXPKpQPP3esoySvYMV0ArtHopV3Iy+co6zNP3LaZOo1zQmv04EJ
ekzn+UZyK/4Lh+04TYH/phPDMMsRmK7l6a5CBhOBLh8W4Dk/QQo+s8mexzI1HwWAwUlbsftVok8R
Wx2TNeAamvSkEiMfBm4CXZCCDgF/RjZcxp6aZqSGTaIkDPqLQXR2GHDXLlKScv5z1lTOvWB9Z0Ya
10SXtc2mPrfAtJm2JLySuB9+2d/JrkryScv+2bATOuTN0FJmgrTu9klzXV/jJT15FKUjaH4wth9A
Fnl6RLk/MbAJZ08ygq+U0S5Qpzn40NlxRWjjwWWdfoQit/gZeOgv436uoYDuIFabBTkU1VA35tWR
AXTyDpE8+fpBGfYPh9QkAi27dPXs/IW6pXE3+RIzduw6YwUgDD9vYHvRbRr39EXfPKarpoeG5Z+S
087chQ/z1gg+Icpv5/RAE5XOEv3NXAYRvG2B5PBPcLAbMFSQcntlTQa+nPSHVAZZO0R97m45KEkZ
wMzsA7eeRjsS5OOAnziSd8xjPXmbg/1LSvN494UHpu/VWPQjBGizBJgAGF6URcxAxQcJVgPBB/72
s8Lm8buwS1xAY+f91fswoaSfIaf44PVKSCfIHfMw6Z3IhdOJI/yEuCwAqWCaEkxmS8pFYuJ1Y3Wj
hmp2oZhIA9LObyFcTJq4gY3TM15CfHVFlLwQ4BuDKu9UBkyPm2hII8yHiz4uuWyktRJgp1rjoNqR
oXL/NzluPk3rJsmQdLKezEDLoht5I0IDdyHnFdLZjHoglVY59Q7FAjEtvj0RH+xo6ENsBxdMdIA5
xABdWvucWkbBrg2Hr1lDtJN9g/RllzulQQs4yyxKUCGI43HKK16HJVF8moYS+LVSlM2CmqE9HYR2
1BX1ZbuKHF3CDu2kPEm1RUJwDymF20n5OL+M1Q90ZX/XFj3BnHwFNIuWccqhnMWJYwOZGa+GhEAm
VfI06aFoki3TrCny50q2vjoaCRNZ4DacHzr2LPRvYHjEFBWcIleCpacXssvOn1SbUdQlAcfJj1b6
w8+D/YrcBsMbV89OcGJ2LupxNXfOH4t+66lYbzixZY9cJCTy8FQ15dskFvN0Vzb2rT8sgSD3nXa7
Df0kmY63U14J5rnd7hyw82WvbeejhhkHjdalcOCKw2SoMaXpREu8Q6kYbzBblckg/ynBI59ayNin
64u8iNRU5bkcQiVc5S2UwBdNyE5aTj+B/RzBVwdt/vBLRjbgzMlSntzUDgVYTLk4/BIm5i7I5dT/
VVzdPlQ9oYYLEMh7lhTMeXiy2GCOJxpRLzTlAFF0dC0+6L8i1ok+sWE7NHIuYDS/Y7G6bv9vr/YT
YL8+vNmtw2zOG2TN89jlLGoGettfm3dXh8F10stt3aSlPGJiF0wkt8U1TNlA43Cce4SGemijkNc2
Mg/WXMb2BTECf5msd6YT/t/w6jTT47Z6JoZl5n4N/+FpYLHnXS+N93I5FGaQOFnvf4hyCKW1bdC2
XG5mung8IbyxIdSleMrGLvdNY2EmS2PH5r9D2JeCBVPl3KAIy2u4k+nZNvbRx/NlqTvsOltfyXkc
dMfOlJ9UVrDcOztr2NpEo8rcFhLqzoFGNK2qVVLNSB/2WQmHbNms2q0QkiIqf6My3amervgj0kmb
hC4RtfqgRWm0nYo3lB0MgshHQi6Anlu2Estd23dGmP3zIOEHPsTNL/8ISit/68z2iRsDFHQr5Nle
dhY/8is6uCjO6MtP+n2y8B8iRjUcNnvN117E1lvQsV4Z9+dvS0vglFcgc14iz6WTAqyH6jDsYwtv
zN/cbTQ2CIURzdbDyw8sSKNEpbaPJcUl6/6itpf6N5zg5Zf/aARN+Ni8vYV6OMm1XYNHlEj9lLV5
WEWmsilWz5X0czND846NAwODSayiQn08dFjMLRWH4FPkgFRALSuIOjYU9OFYUn+VE/1vSCFg1j/h
IFma2wRQrQHJBK+DHgQ7fuGDtWnm841CXfePwduLYmb7e1LgM96l5SMK9Tg1xLQrAuS8O4MmMfKJ
uRKLKfc0JITaFkG7bpwPuPX5DEH9pFlaQrJoFxanXM4RCO7jq/ZtHHdxMANd7/V43+g1n+/WeD6S
clM1vprQNDxYyT5TagtlV3eWVTl8+KSpXjHMJuejBoPt9DmLZCkoGscKj+4syr4zuXBUHmETZoPT
yARBpTbcUo2g4IGFd21/PnTg/I0DZ9jT9Knl0QapVC0IVlU19OsqlUzhMdfo67kdIXB7B7an+NS2
r8ZRk2e247AfC9QhDwIInim/2iuwdmhA7xK9zbmxC1Wy6X7PI0dwXHAw4OGq5E0EWkiYZZAC8GOu
yymzpm4sEP5i8QwrX3r7vqTwbmC4eJgZVjzXb1+HdNUJx87KsBQE2QxNGE3SO3OhEyOnixE2BWQv
sZdlquVLMv3KK7wLbUCo70N1JRu6nPZyXDMd0bCoNGl21Aasx3zCYwBHpZJPLyMf6wi1ZOzbiSZG
fCWihiUYA7vEMqkZiArYWy+V1ngllXc7lTCJI4Bow0m2dVHz2Zgryl8Mitud55PdmV+NR1IMw5Yq
Nz4Hs0oh0jZVrRUB5L9LX2DjJ7M7R6ae0E9iJjKNXew4WWuxZUOrJmPQLh2l0of9BxjEIOgWe6Ua
fIxYI+HzUBpy3JvN1esYNzDcrGVD6a8tEv8i63MU4rqvn6ar0aDuEX4Z3ZOC/HuvQWvlO3SajeOu
YGihzcMSdht7uD5au3714TZNinZs+Ca3/y3cjg14GNBmGGvSGGikqS53K2S1G926ooP+5liwUIiD
M9KYDWM0QpDMv8/ZrfyuQF0eqWSYjZ4MiiNYOiW7pKxft0T9G6sew6yyISGIKCVwpeFfeVRIrrJC
T40UUhvTRr4SFWOiojp+eKS5037aj8iHX1vofccJdBnwCbfSIJ6N+96PpGyitd1/IYHnBQZYy85c
VE7zMLSew57V6x+Y5jX89e1OlTp8UODz3gGNuZuRO0UWDW+ogUMQxil0EPK0syqQN0kAcjE3kM6/
fE/A3BqFCIYE7IzKhk3AUv3T2tK2JdraMf3VpXXXOgfVfAwbclyrBsPiawORWwAS0vvXLy7rb8ua
094Wu90/JtbOp7OYs4tGrqpYJFfrZb+AQv908LNsf+9E0K0nd+MVeALLR9nONCL4Zy7+PVBYjf5v
NZaXn0Cs8XYubIErMvATELwilRU6fIHTM1vwkGxB2DLbHjcmWOS7KCr0sOGIrIkt3G/Y6Lz9XLUj
vHiGX8s2HPKeATPO/x9+XAc0jNE+JULAly0h0sipVXrGEQ4X980JWPhyBZGPYGAIPAk9LImwtwb7
w+nk5kRyczCPXpQwPvopHEK2x1SUYW5Woj+OFYWso9OeULxS3GVWpDbLuydriHGQegS13QBIh0+Q
recSpDYOVhKXTEEAab6XVAaPhdMw+dLaQgcwdBOOKudf9kmWBR/Z32NswsgXAn+giaLIUPIioaJv
OolImVbnDosuYr1zrOxGSGw0ek1ap4nXBSFD//45Ttm2rSGrboro2Q8rjmjXfGEsH4PzGysQFI3U
5p/hbRGptThb8mdO2C7vDYWBHvMQ48EGXVSy/V1zq43x62vrGGYmoXf3stBmmqeeov5VLrSmtjEj
aCrGOSE6GmPn/EENmURfMepb9arNVXNWF2q/uYy6cpX9rSACBlxP3JIyrHPFjsvvS24X0GieRJ2N
OxmlXXXWrRyciPsx2ASn/Ha25whwAzL7do5b0ZCHPZQYmBEtdqPpOA1D3dgDyKmrcS7EmOPbprwn
3OJ2ZiLh+0XOiI2JU2LBivO4vwhTlMUBu0/LtLrTSzKiIdpdTYQ8RacmCUMBryAidqG4g6qqYLRs
Hw0l2T9WRXBXWEqQJ5fgqOQodnByHGHUiBnDLTuq0AMLpb0kNBjT2Yndo0hSpNKClRzgNuWxPVgA
BKDXLcbMeoO5c24c7i+DxrVqLlAryh04DDuViahOjs3BGU1rksx61BsYgEKex6tCmSuTBvPKKFLM
WWOCHxG2LSIByl/24+68O00vu3J47IF5KLTioS5L+bz1ffzEeO9MxJn54a8sbVnMJK1lxWb/jxLB
7VslCfq+jFL9RqelkPZfWCyisuo8lRzQDx88XC7jIM/awK0JRza4if+w4ltbPdeyMCm2pPvb4Rfh
fcjtynbYSW9PX0IY1fe2sPRUB/EtauJ972sQ9c5uUX7barUqoYkAqb6/gO6Ymeo6DaZg2ysKJ35P
9mSmspQ+IsBaii2oQXqYj2tA29r/6pil+Iju8UnwZGmKw3R5V5G8ExNSz7oJtV3+7WnjBDZyL9Rx
E9c0u6P8oJ2DD0o6AuxnLQ63/5h4lNM7hLZkmC0YOjpIFtwN8kFpig+1zKme3RiIWJ0SEOYcZUDM
Q1QjsBPcNEzEgLKF218OvBsxpuAF9mrJ8godwrPm5pJDMRbGv6UYr49OYI93w0tcuEmtianPGpUq
xu/+7ijigK4YWi/brIf1/R0hLLlZc/zwLK+ddVMvvOKlFTxBCxonAAb7WHNLD5Dss4A+tCVOJxFI
TBTXoqrIC3tzgLoIwSz6rYARaJqggzCNNzFQVOqap/G7vtLknUDCOHvQ6MFw3nrGCbBkp/5UxGST
SL+LZODTyB7c30hY5fQaCaDu6GYROSwpwrilKelOfdUHQ1/3smaVD4+3UI66wh31Aj5/fFM3T4vo
wanx+yKfb1qfAihIlUG3LzKRM+aL6k9o7zhhMeb3+5X7k4qmwh98EqNNV/4oyM/EuYLgvCXZlAhr
o4nlQIEmfaqC74IRGqbYD1Fj4sc4p6JshpXlC5G9WecpokDDJ3YQRZLUOmsMIT77SnoNIS/27Y8E
85R0qHZHHAVG2aFasJ1WgiQ2tZ/v9OjZbPyOI7GC8IzojyZ/MVOaabl8jBD80Bg7cE8nLfc104nb
Xk1g2WOqy4QJEMA4DvcY6nTELsVUL09JfbXKjmSCLJWwEgMc2j3yB/rJmIkJZEjbtfkWCz9pRtR7
MZDt7cuRUR62FowdHPlc2e6L6pbBW3R8lRNekScWpEr6esJzdbMtD5EgpV3pg4i7b+yy/q0n6jr2
f2cBmrzol0fmyk7okAP/k3wf4ibNYhZ4ZGhdJGG++CAyzXfp65mz5b5v28Fe0GLAeAuYZWsEvKQv
xYkF7hbkmOHj6GX8V8X6iuq48f292oRoPcdMScp/Aa86w9oz3/v4IC3e/Y+lS5ecjk6IKfu4fvDn
beQK2r8cp2znJW2p6DVNx9nJ8YVEUr/Rw8T1n1HFSlKdCO41Pf3ifuxAO9MBRJZOJci6j4+fVL/+
uXNJMXqtJJ3xhkkq1hUm9TYRcNO5rrcVVP4zQmHthpGqrDCkrg6w8imoujfvETOJjz2r6lrxH2hF
N+gXg3XuzcUGb2S9cA7Xmr216Kd8zhBJe2JvHjxLXttp/E05Jt/eFrLWopaC0VYwija8tUe/YFUU
HaPws5hfdhdUl87l6700uKfhwU8mOkief5lsYS7d4fsSDDZRltnoyRJt3nKG/Un6LeZpilwWuM3c
F6sq9wj1P/O+utO8GiNjuQRjX8rJwFbxwEs7z1j5pL4bPYqiRg/Qs9ui993m8Zv4Y3TSIxU+pkgH
Ggh9DwRPZQXDiOgCk7xCHLz/kc+unmnM7slM36+ed9bW9x3AtKGSqpehYIo8SLBC/7W5uAZaA9hm
UleY5CXAgcCdYXwV+Er1QdvhkBA7qXZOYOx3WtnjRHSJGwvxipaTnSUzL9Exh+DGewo1TTxYYi1A
UxaIaXKGU2cALntDC8XWQwl6Cb3GSz+AsTo1pewdOWmxjIzKQtIpJiov9ywU9k8JgPrPx8TlBNM/
BCgtrwT9wWqZYceWBaO+lIecUZXXpPJQQAzxuc8yPkAcUBnfZQWsUDXN/k9WjY08OEjPr3SYVX9w
aGe5Z71ONGyZAGn010YlRRkWMVSmhBlgsC5cDVNOGRQSN9HlXNEdkoDAog/IM4Vc/DKPxLaHvLCB
uo/L/leJL5+NGCVrAQwWR4gnYxd0f0nR4sHFf40Iw0Dr1h5xoQkHHWmyJ1fyqNU6lQJW5MIyMOaE
cQQMJOwv8U7AXBr1ODXTqy0kSDbIDm8j+GTffLM23jm8eGoX9TzEE186/R957wF5PGPQyzls6iPp
WuzGOBIGpAVLW+fRL7E52A89OZb/se1RuRvaSdaSaSTbkVbF6Cz9HhdC/1fFWqa88xmk24Ir7eH1
2sTektvDOV2fuu72gjwtRmfIN59lEhT9izHvo04Q7CudVZgAlTpuLx0GFSks3XyhnFtPwU54Ig2m
E4h/+VI9d5irJ1s8VTSeZWKIkMoq2ysDFCFkWEFH3CwDxI6AzXuUMs5nwF3RkNuD95mrvc2t1Meg
qe3/HVxb2gdqXC7MsO9GidTt9X9kk/Z0/t1yTZsfXBfSvq812iI5hTqnR/vzTKAk3sBJe+Tkt84g
AK4nDaGLcc9CBAfwcdY0R9iPYVrZ8Ohhb/WLCH/EEwh0B+8HL8I5/sGy49IwuoLRmbzZ5kD54Fys
J/oOSvXeQxFvkTbnbvlCpt2tYck/Xg7rmY9Ew7to5jnOSurjX2KVsM/Kl9i44uidu6xQczlRFwSa
56Y+YgItnX0fA5SVcQDlmYa6N6egvsZNKiCHaa3gs7kKIbgE9gHBuICHYCPGcNvkJC3rQ3KvmiJ8
HoJOaSg8IOjBMlfiZ50uN51V2WCzQ7nXXzvst5kX9JYmHO086u2ovnsuT23Vb2x8SUsxdWj1uOrj
SRE8KIMSsj3RDGFw6PlvZ98IXik5meuSVVG7GsTK6ZTnfxBj5KcAx0w4VNkU5zRPhVbNtN64KiQ0
O0MQUPQVyPNcAU31zRBubNeW4q69OeTt/15IfH9f7yDLB9snHj/YpOtbnBP9jsyF8/H3VBCoSCsa
go63moVNcoSmu/75KHXTvrSFz0up+pXzu40mDP0rhc3NlDYjlxUY6P3Cm6ZTK1LBFHVHyenWI7IC
h65FGALt1gPf9ZhtuYrujeqVLTgK9xKb+48pD4W11xsCR9iS4ZWFRvD6RljZa+BpXg0UPpgdoyr/
KMxy2KizjQXg+mnKJoJMVIsPKXDosveR3nd0IwRN8IHW7jCDIACI2+hW+HP0lJuyaTYUXM98dN8j
YQiTmmLQ6DJefvWsNgHqQYOQyPMmzDgOYHWSi1C4s/IifG7cs9ScEmx/fS/1bDaoXAzCkeq6xVz8
BJhBzCKGeVtyLfl4aV4aT+02uc34xI17jnUYtwHADkN9hpJp0N5m/OX+7W7VrKQsa+lW8F4IeX/m
7OO3ypjwE07iTNQIQzVuvIYMhbil9qRrY+uUCmblk1X5sIrcGILDBoTc2uvuVCsDMGgvLlgOH43C
XtHAzgmh9ytaqDcR06txPbHMUxcr0Tgp0BJlXa9yBIN6dxLg7m2DdeIS4Cp/sk6w667MzwPgUmW7
/3Pj0SqXyCrBpKcGJP3khz+TZPNqiVjKy5Xygm21GTzcuxS5iszTwRwaZfr44xyG3yMrWeCqLGQq
48S4CZudqC8oTsP70GHCe9di9bBA4za7XN4bpqUNsmm6/1kDqk4nFM5px/ohFOvO/txy+qjglZEX
VTl2NAmjriwnhMjxVzcDFhcTngajdhbIhd055UkC0jSbyC3joq/kn29OjLvndTcooxWSTx+ri7fF
U4c8UcmhX6BR+4Gi5wTNCDwgPa8wzvY7O22iLtBIQGvwwbMspItUqc/xlhq4+WCbVGJU7tlm4p/H
A2lGlcSuujgwrZT9u4+e4Vmh0HUg9SEXszYxc7HInn1nIcRuP3Cr1h0okVtVFxZ2qSFPHi9Zw3EY
02KzC7zyvhenlLmIrIDxzJZC4EOySmQLrY244UbenSFNEYzeCyqAjJtZ2+/fBQeRK+DLeDffkZL3
eDEyGCVzla5ferINcOA59XdnAR8YVaDUpmCAGyKi2gFYiDuBm3oaqHjj+UlGibnv0cbYOcCmNPp5
MZVEwnyIlhxytbWTywWjb8TtGmTCebYATt5MAf0T1eQXuqF3dVFwLy/IuePfisyh3yELgP0u+yBv
i0y2LCwMBj+gvPgohTNXosn2uw9/C8pOKYvUNVS2yngnfvFE1a90twgb0Eq4Bk1U9MZuDsv9mF/W
t4aRI25ELg3ZlvlS/2b0sN0XV2anWTSEVjVlbqhPto2TUfAQ4exDWgqquoWAhwmv/4EkZSHFgxqm
y+ZEE3iI0KyMm2wviwYHDepWAgMzCj3Fv+NdwzrUtMHhQlOnbIaVEDrd0EhI3TEZ+96YUuSvxBWS
6CU8t4ASKimRCiVACpZGrsBTh0ddz9gOT6MHlmaM8oS3oyk4ZEUHYMs7bXocE0k1wDUU4aDTYYFt
P66s6DAekr+nxvn/axjbfCtl8X49qmh7TvzU6pJ2W8KhNAzI5nx9IycRll/Jtrb3xuNd83xkZ13Z
9ljoQFbavGojaVH9STXNwNYizBB1D05jt0/GcF4AhXvNWepWaLaPPmaWy/HS4376nlB36uJGI4dg
EGQ/PpODvi/k+nPHMUNCrWeQCVYHIwmdQqTf609RTyNaLIgdeJx5dE8NXRD76M2K9MJZ9ptMPko9
GqWrfncAKQIOoGp4A48snAel0X3j2atUFjN0IC6YxT/v3Ka0yvTVW/uyqbFNMHBi01LqbWo6zO+6
KMsPbxf54yppWw3dXWk5JGE6KshKGjOBNS/9tIbBXYr9gElD45b+c1uoww1TOzbCV1XUiS7EXuYW
i8XmiJAMPkTbz1TlB5phIdq+dDeXxugn06ZnRFGJYYIEOANv6DHQdobjVopWR+ebQgWvZgIxLsNX
pusF9trg2jPE+YzRLSHUaj+cRSG9W/FFQ3Rl0ezaLGQugEH814vcgvKfSFJQI/lj/HP52uedunIM
dS+mgCkEH/1mC3+y28xklqLZHuT1JApui7Wzi8doNm4zowmw9cRCMY47qWwnI9PrAiCXhChc2oSV
bqfnt6VHuNu2zB5kgWhtCspz4RDWrbZojCqsFaj3CQb4qrviMyuXtcLVzUdq+fcGmItpdVYv2wq7
PvU10pd2F4t1+1OPwIcOXkodfcz/qoM22XVnZeW6QYshHOt0tAPhvGuSh5FskFVxVSWtEQRrfBBZ
oLw0iCZrx6JRNwWAUfBtD9kh7BfGMKVUujeGOfpRl8kvMiFeho2f6FOGLLAm1LeEGxbaBlF5kVxg
MRZ6Lv/DnzpUeIb9mSrnVQsVVuw3rsztdR85fQY3Rlb0n1kYanQwJNXx7dMnyXen8MHk9v7vN6gz
LfbDM+6T29tVZNTNDG9Vk0nrtrKvBDQ8Zynu+pHS5y6L8ERUfPlCnNi714ZZbhRaCO0iYJnoUy37
1VcAvZxjkkA7MvVezIbZDJiQ9iifCn4mNcOuE+18jgquowTtXRz27Ai7+rW1w+Qr7+Cx/OkJ628L
7s1lUeMp83CwLHjDczFREpexDPf1loHLk4FMhvXcdBKS4WwYMUwyOCYcyW5ewdsGakC6SCHWoeDQ
LKQuYP3IFtv7RJjMR+ZtsOIvjYOv7spKdyCx21QLh+OlLJtuMKPyp54le8fCP/P9+M0tv9dgkTAL
j3uKiA1kIzko2XCN6LnL4aXDdNMfnxGB1C7DQcgDlNjT54+j103PeSf9uwcTIrt3W4o4u9Xg6IXe
ve6F3Wqabe2em1GYKgMTC25AhZQ8xjptLl2xPThrl72Q55zcPvTAEpy1lMsIn9Kexsf7g/4W0/mv
Ovyjs2BGolYUapPqcJs99WPL4bZZB0MD7dHqu/1PPZxyXM4jCTcxq64R4h/Oi21opEUHP65k8tXv
TPMS/7NomEjUZvMX/pA6kbJZUOeOXRaa0gp91sADuI95LGWkJvQ9eMW0s4TEJuhqYukQ3QbdB3WZ
j113Uyw8ay+QKwxNrcbnOBX7U3jc1EE8M3WfGfFqx9PtzwBPl1m+h9XC1WkuD84lrIdDbYBfBwYm
nuKB8sj1LPT67qNfUIrF9/6iE13bKc24EtrCssvzzxU/IPl/m6IEX6GtENEdML1b9ogSIAZ1KHZ8
3XgxeoMByXceoNuSQgj80pU4soUnvhj63G0q60lndntP65Vzp3lX7EskRxvayhlL43GIhmeZR4nV
Bmlk/4cq8kBV7MrDZAMShoXZipFrkEMJsW0raFpMlpwvQ2ZpkS/S77IeHtCr4dVDRYa9VxOS+hSF
Lov0THz6pge44Guk7RtxUEb74vqVwVy1c/nOxqS18AcHd4yT5r5ikkH9Q8zfYo2V+xiQiomn7u+5
01jRGNNnEQnSNdXvuzMmJJOE5VJ6mGQ1Fm2HBVImG+zoMfX2jB0O1z3e+F2IK+GhJFWMsdbyTCUK
SHYH1cOp3NYvMqnSvZ485r5p0EqPuwoNMe12NvFu5A44TbocxtdD/IN5b2pzGUi2+dkIGXP6oiFg
aGpeZ1P1rOVbXWK8gyPlRmKwOuX4pNEHLDchMWnIbxJKe4wNFI5dSVvrdF/WSfvSBp5ijW6XMYsV
cyXT9r4CS07SWPxVNu34c8E2R9d+pPjzBGuwuYX73kyl6Vb/EByTM3C3FSc5PdBDMXRVCCaIAhgS
nf+8GcFOeG6IMlmhm8xq9VPCKe2i/Q0iS6mgGxNoKezbHqpMojATa5YhgKmDEtHAVWI89MxXzrLm
6/iOpKa8Sx7LCC1kSiw53iKEE0UmIkVQvfk1AujHbr2DY71/JdoPdUqHpgYp7aSsTVWMskwRIDJH
DHCwbAWDO2y5+j81ZwvDH/Kabdh+B5l8FxFn18ky9+mwt6BfZqcEGJsoab9WHKsiKD5tIcZMmEZI
oXdvtvauhhdYa7stlXhs89cga1dQp62K24e8TSLEmTunjojWR+eIPme6KMg52a0Q2NedpjuU1qMe
+7HSrpxptsFOOxshD2kH1wI/jk5CCXLdWok1jiHVKzkShXpSpJHVV5IFdq/A1wrFRR8roRAUi/TW
NzrqFxIIopWQR6OEFcFlvi5Ti0RlKrVZFWk7K/NgmdhGqb1uHZa03k4leqLubaOmmF5J6KMDWGIc
wlSF64xx/2IzSfuqKhhaTdgn7RbbCjv6p2AdcN+tZJ4dpew/mFlSV3cn92PgFl91ZgJP2TaW9N+S
9VmfwhYv3fRVRbMrBeJXroc2tleH6yOySvEfPsGazUEL3OrtFfx5kDpi1F7h5lLS5ohOja+5fSwO
oQkSWdNpi7FGSPuB9xf13oii8yxjBzdrWzEf7+P/beTJHRfrcAxVGyxbUIdWIH8nQ4s9VsgqHf7k
oTnQdRIpGwc8HLHjXWyqzT8+G4AIcfKvzQJ7it9TFdxAo0XLHhSS/Ln89P9tI2fLCwgeoR2X8dPC
ySmo0MOhQP8/CV0mkpv5qRyW3yM+xyCgbdASL49yeY3V25AgsgqTBc4Pp3jzpJLBhiaD0HDmHYJx
xHhl/IBE06RIVpyPjAPJ+vDDGC3iTuL+MvNnEb9elHZR+2hHhH01ZjT84YV2LZBOvMGovz/95yof
lqJQeArMu9ZbQSg1WYMKoCE23HLTt0J0GVpd6h3QINATV9kAlzxJnQaruXa5QozPnBZdRubOapSg
RlTWZXRu4J1danj3CVfEyEGO0V/IjcfoMQzdIpq/P9+f4Mzc0HrCBOhnCM1OoTV6BMn3kH1Dy30b
5tWoJ19i5O1CR5eX7w4mt8RFgpJCPO+gQzbhaCHCEDrDewHOmijJCttfSio21vPdVaVENYPqiACr
i0WuZULTwJvJ3FYng2W122Zv+JboRn7ry8/hV6zDWr5RNXmKZkBrhWlkxkZTR/TLycY/8Omf/6uS
2vX06jY0sZ6Bdgh3oJit18S+2phY22Ft8F4DBJA7h8EyTpcbTixhZ0qRO55PdMKKqcT+T/gYQeOQ
DT5aIRiP8HEYKMZlMpv3Ok111+w33zgrHKAPVTChfz1pbE3H93NAe34ZcurK+ssjjspPO+knlzYW
iOTky9V+vh7xCrrhbcukQTqjRN0M2nnJghw33qYl0mMzcywsqZcQrZs1yDVQv1j4HkSg3VjgkUB5
dTcC1cE0buGMSOcAuD0RBeeMLBH6JeCrxk9RNJRE0/mNBQmnhw9ebTgIkjXxa0b8+LoGMPgtKXbr
e2EpXgssysg2x/NSf2Us3Dvp+9kgROc+YvnGdJdYYGIqL9P4ErgMCd4clHxQKtutTfc47c9qVo+e
RbNqVSlgvZkEwA3TSPiuqaB3Fj7kEcY+znQS07OGcgASRVo2IA0AsO8O02qdnCcrirQW901mSsNm
tBYZmiecuycfd8Byt+jA/TJp2JHNWbqCSHXbE5Gk4U2LCrh0im3yNQidh4564phu3JPhLX118FaV
K/S4DxAM1SnBbtnavTrd/Wty699VzjcHZ6E784xL7P/F4uoYFCR0ftw+bWjO+FI32gL7fiYrlwGc
TjaExhnC7UJSQlect16ePnEmzPQMJXiiQ04ur3DoO79UwGFuxQHkePJYD42ads1i8KeK5RTUEhfN
rLUQ4nXyuQqXHItXrFRmaCdg84jOUxvuT0hc/4/o4T2SfDHn6rlnTfXKlFEtW+OvDanqlPVUMxXq
8e6rLCtvCg2DWxVIa0s6aM4FmBFSNzppDw8nogI1LuRWtTliojdvhMZ7LXbnIAD9HVBvBw4CG8Ze
pzPJSje/VWMz3VYkp63E4RcYztu+aN72IT8tXAQKMLQ3GqPkKaC+o1WkIFXyNsW5b0+qNbNvtDZT
aLmkbUoe6UKMpCekalCaWl5bfSyjWDswG6p6zEHwndJssMN3DyHcPvKsBBR+mTkpoNP76DpSV3cO
R8L20b4QUMEZERJ5seu8k2oFqVait6mxn8mZsSCT793TgnN+j0bKDULHLMBCHb7WXrhgLhS3TeCQ
xbCr0RjkvJg0ujtCwEtOArZtS/Kjca2HTcu4AYD0LcXcp606Fv7419UE8XctMaFJWHhSrqIrWpUe
zRcmZDQOcCWEIT4m5OGmITwimetRgQDNgXfMGowfQRiv6mZyepkjeQ0zyW1G1XL0wMMoW3lWBrMy
q/mbzZ6b/73DE0cLvbd+708fAuRaDZpR4YAmPaE/y7gF4DQjc3R68nFYJbewjlxeS09Liqo5HQL7
x5wgIwzizqp/RdeIvdrlUuL8EEOqBlal+dZ+cNKqopNErLHQb2umldMzS70VmZpLZOj5ommzGmP3
Xe5zq/+g4a2sek3ndEPMQcuOPdc8+HaszwlK3utbNj4+TgKEir3AnIaM51HzB93Qv05MSP7Ghdzb
w/wh2xyjzqFpF+Jwptvx3al14f6VenajRMVqpeGLFzaeeJPt7pyTotn1cC00BfAYuslhJq7MF+jr
CUtWpG6ErjG5EZQbnNN4tRw+A+gY5e1btWq6SGHu+ND34CpaumZqT13RUDulEgUN6zlvv2o6mUnc
0f9vQxTN/VA2eyeghdmKDhmtc2cWCJtjf35VTl0rBkAR51KCxWf9SqqC1IEJG2C1Pz5I4rVjt2JZ
Xe0UjZusCCZEMqZqV3AGkqyIPHAp3kmXz2BHfNAk/YUsPjVAYlTZbFgkELBCWK+2vdJ1ZVYHAMuY
50sHdtaPPVHuhwMrLDhiHiB/pB0bH4WC4Alvrqu51b0h9wR9UKJificfLi8QokVmYVSieivfXArE
VR0wRIRnOnKD2X3/LQCs+uVDAw/Rl9WCsb/6qOzBmSe+oazYXqroO0IXkQe/vcGisjWqFCdDoeGV
jeBx45v632ve5IJnAS+1jEvKXQbBm/g4uwU+lzHFsXlO3weTcNpQNGBh163j3S3Aurmqz4PVg0Mk
xjFqG9Ve8+ZwYAwmML5+p9p1qI/XpvJF+zJqiBYXR0c9PPgD8R/USVyABcVzBTI2PdnfADiKxUwL
2xUC66mTtOMD4IiACX9LRqXfBlH5SMiuhAjiz3FF6vuE05Xq0YMQUm8dSL8HhafSFoVNF2/ILRh2
uDhTge1YQadBBapo45rl8+iqjebEJ7WSzwBiAWgJ/iygKkFHqtVwTeh+nquFY1PTKKCTf5i8J9Zh
VcqtCNTpACCIPRaGd/sNZ0tQrDVGZxp284dQHAYJ7qqW87CLUN1Z7vL07ZdGaBZhkeyT65NT8vh8
x5qrKvyI2mmXS4HJ0Hk2edolbnYfOvMDF47cC26Eisz4pG/7xsg5j4kW36bd1RPI/xr6j4Av8Flj
iiqSFDa8dwgAGiG604d0HZ3NNOssFYiF747Rskahq68o0NyswRbrL/6By9wbrkwyd9kIcUvNFb4R
Vlef1QZMNoy7nVUTaupYvHBs5M87HPgsyGcEX2RMYjLwkVgHy1zUCKY2lxq2bV8AGKTmW1Ac9S7U
uXD2L2uufgIu4VdF6kz2SgOwSJmI8VkeNH+X1tvscZsgoZCXM4c8mM/aOyDia34Ql1cZgTZJbYbl
e8MkcBm9Zj1h+3kJnH0P9SVZTpwv6l91ke02wv+mDlKKbalemAvI7OvNcNASWz/MaupYiumb4kjU
Sk+KH4tR3BChBY28O1jbZrOBEzZpj4RV5SWEPyrNANa/AmzqtTT+0ss52hPUFl1iEJfe4XD4JfwA
XUWXEmAXjwfONlbXCasP5AiwVzIxMlojIdiljbYAvlTpZeShUCmLnz7rGq2uN+4iMbZyg4JVmZU1
RtzLoGj8wTtYUzdsGiHNioF4ZLn4DnhWKTXwJVeVu1qD055O98LbC9c1hpkVRpyCDVp6FhDC1O2u
kTvq1xXLpjR8G85TrmNQjP4wt9Z4V8Nxc8fk2uOCP/iBSl9RxX3srxT3ecV1wjEHaGvbcXJbWEdU
uSGl4eW4bXYh4C9+RPHFovTzGA5PMtdPmRlXkU4kE78h54MWIRY2nZx0miSNgwUDCieR090ZVCm8
4dCwgiFOP+bEZZbMVWKJZYY2kgO97rjLQo4NvUym+nZ3KrqPRSw24/6XmppwChrkReEML9PY5V8m
J4bCj3VjRc4NBJoqthCVGiSLXJ3bpi5fDNjxymNiHorfvudzZHWPe2Tw5QmCTdE4moxWkaBghIed
6yDLoBLhLXEKwlRn0wtE+dl+3k0EWGDH8fWAWtIu9Ryb+zIQP1MbAQC0tXhi6pOLowwU20HcJrf7
CEzDi3HuljSpG7NJpTOHfKDYXraBVGj5OJnMGg4CvrSdncNWSWD7DUbcqd3GlMzWgFHMtBHYBduS
iFB8Kj5HD78gNZAGA3ll3orpN+2TCeoNCcXwlk2HP47Y9rnFAvinnTPIVA6lNuVc+f6je9ozbuc8
484JU5aAK3pWcWxMVPfLlyXqZdC898g92RdCwgY2jvvQcmzVMYiBSNakYWxQz8Sqp5ba6+32kAzr
RPd41kvVTUrvLHcpRy5cEJ4twqkUC6yS/0cc/2BkIA1PzBuYvSrkPhZPsThTnwLHqOprinI/sVtW
EhFYguPxVhAnxAu9nM490ms0NtVJvlP1IpTt781cjp9bsm3HfgOVXyFOyEajMssh8liiXHUJarRc
u2ELBcI49g3RMdhlLCURYDy02YwSeT2+c4ycMJ/FwJZTBrmAQ4SiQR5waMmcthKcTqLcxyTsfpHY
KhJqrtcgBgE/3vJeiH1dYU180vBhoCGVtDEbht5n4yvWBV8gE3VPy6GYORRKDaKlZtif7uBV+O17
tctFyEQaHsYVV894V4Quqj2aFh67hSZk0WG724D6xbUp/RVPtqCX66fxmCrLiRqKwqTSkynngjBS
EuF6hVj58hZrEAsHKj/vT9/T1liYtbKQ3Ty4kd68HNYJBAzUvQvLeKRROQFFLmQkMXKWylgEAprU
iOcWL5MmO8muKotHJNhwl4hs+LkXqFsiFDpTJWE1r9DGt+dNgrihZwb4Xm5EhH2dfWWpHKSg+s/k
L/Z4OZZnG6ySnDpOXu0gXIuLDoKEGpOvnXeBxHhCil+KK90NEheRPbSg/h5PodfQSaV4kDfmfmNW
5WzOZlffCW3ajBCX5d9EKFDszyXYSdpPIGizkR6iY8/0QtOZ4DmVHjcMBWq1JA+RdFClLs/quK5M
QZqtX8LXyZgLkKl13qW10GSTHHUclO15c+Mjp6qUiqCn8xVdbRqnTkGT7Z36ZHuMU+/NNlf+03JH
FXmtoOGVDXhV+XwySg/DUZk4G7Wx/vjCh7jDrzHfnJ5LiLwgpUTWjbIGCRL3dBOYsI0Ngbx8YOe2
MmpdiVsfQo9LWnSeHw3LfEwe1inPhgdH1tyx4vb1pIEOsbfeiCglGQq+SHy22LxqGyHpSs5UspUp
7zy2JjIVFUzqelKwHDGX0rIGHUSYd4YJBKUIbBAHw0bIk8ovMpBPkFwPxOajIuV+0LxpsCB3V4Yy
iqP21c56407ULDE7Iw20bYJEOQPZZgGbj/cZfdi0nGybf1uTJqHL+idqrCBgOZiyVuP3IWbj/71P
0XAJgREmUPI3pLiZHpE92GB2+Yus1tmFHFFEtXMePjR6xWhc119xYZveZguOAhlq/NMUO/OajLAr
pHZvXhepDUwY+oqcX+bkRCpwm+yUs6NkiVsAOcQ5CzPsVjp9JpPAK2DXkdJD3AFnN2OqVDovOseR
94jcpWPSBVzap8cYq0xTX0SujDVviQE3cKhwwDhgotTw2HWX18yZuV5jQl3ANaZqT7EMGVE5on9K
KI5vGRzuAg9lCW6xaIytGzG/QdT40Q/Me9/2HFZO4b6jgVyG6YKBSyrrGD4JDcX9aB+ig6qBqahU
i8Z9I21mioOEHn5ws/gZK1SdFilKpd787Wf6SkxlXCK4hvZYUjZ3SuLRz7xiYb/d294HYVMaF5DY
WAl1Ojd20Tmnj5Xylg86+PQpjU+DnWsGhtD0/3bGxEDrHmb7k1RCIfeNFb0zsZ+bHk+tZJQoHgkg
KZO/337dDHRgug0nAD+6UPxrAPqlJyo0ja/z4evDMsm6yyj2YpXJOxxq8HNExnBjS1Q/el3/Y7p8
S1EEPeBrDmU644nkoetnbhDb4MbDVs5ZWZ1X6hVOlDsReLBog4+QMNrQ4WSZQYHUnV3wqaqwF8E6
DlqaWMSDGwr0w5sWnmRpANAtIsGa3azCGxZIEkhwvECH80BG563wgB4tMU0CzRBMFBgylUsCpXu1
kEyPW2lUHi+ODDlBq6ae+2TdsoqGfM6p19kgMIbb0DxRUwJbB0A0gmnG+VF7XjWNFSrinq/1Ikuk
SGRZTsT1oYalqUv3crvNBpJSyg3QaDBjqyo9x0N1SC3Mz728C3wpcBruxwDeaPQbhYAXxmncxUOK
UnS9kd4wPZH+JmV/ZEDacZqqLPV42bMoDsg/hr7gLm2I+7AQDAkOdk7lBNamYI5MtHCsdudtD0gY
jsQHWiA0APTZ7ABunmEH8nHEuDrjDxf9iMVFCVOQzzh5AkyMaVLYQycFAFReP+QHlMIqOpY0mnl8
szmjVcvCRoBiunkmk1ttllBpjO07rH/U4mMTuF2XcV7HJjznIKug9K08LBUYGBf3FBTktPxj3qs0
ufs9f4nReMLXF2F1GD1b68o3NKVfbgprmh6oJekcNEIq/G6/KzwUfrvRarmfldJ6pvm0MM/KORy+
YCxzSumrDTGdsa0sQ5Fx3jx0gbil52/DY6E+juwH/+41uv9KOZDMWaFWJPWHzEnWmsovQ6ccTY3X
uhMrzFWAvWi9xdFHhLmbzHDRcGTEk5hZqSRJPuoazw5vMrQ62SRpldfISMX0z/bCVyzu42LpoMN2
eG3pXxMiDivX1g4wNNIWoyCs5HCUNNSaaiZr7TxPQFmTZSNkc/JsGDiwa2e8cG1f/YGDimY2Tkgg
Ji2+STcJXurPOCE4jmQtZSZJgMh2cUCqriB0eiIBg3w7xHw9ZiwMQLQf9uGepiARx00Q1DEvwSdo
tdV/0JDbxQkJ+KjmNpKfo+PDmd1llyhLlsizqcfqYfPWZHWqxY5IVqfBmlIbnMN8peb61BDDK2vj
TDovw2TfelNTVNRBVCH7wRZdzozuKcHAY1Q25tB55FcqaIQLbxmWUrmQO+JL4UyfRvaIyff+gmHZ
+gf8ZAr6Oib4pQkNupTP9oY5Qm7jKQfW1oPtSOTwYJd13mWFcxjb2HsYpmXaFdh7VYfXF4eqWuAX
HwPkWRH3k4IJ/q0legt/FTQ05erZjVc+bOPA0NlO2R1fy9GfoH9oltkIl3wbHVkD2g5TQAHd9bFY
x4MzAaK7x2qfsvRrwUuMtDa3HNbdNLHBE9d519nd5m4RgrlO/wMwToS8ulE4Zy7lAn/mQ3dYPBHp
I8cSvgs4myTtiqy3heXDmr0ufHY+9CPuFuQmkmm+6dyheTQx+Ufw33Eq4wZI8Fst9LRnXg0xa+EP
N5wnyHZb3oCq9zsWSbl1wQmV/9+bAPByllkDaJhpEl2UOvP1G24rvf3gxB3mFoqWigTumGC4zDry
0wHAxCg94ku5l6Cux7OjQ0VipCGHxdBAo1AL6mWtcnD5NgoERnCJv5k7fvvyAE2jTdpwnyW/mynA
pbHrrI+8PYNU8+y3QilkFPvgccV8sLs3LeVh2oDfhzP+UtKXa+XNhCk2Og3m4jUyvbYQU+7VtbUA
F8D3jI9bmiwNv6quVbdbC0XEQNBN6WxmR3x5f+coomsWmdF/nMIj+IumZS36iafm9tf4ZbRta6H2
xwGYQb2Oc6BFfaaokpYhptmR9A099uZLMhY/WkXmv1qO/MUEbuJu8V6wF29pobBYD85wA5Z9+ZfA
oFT6Wxf+6hY8yz+zguZnMybnoa5ukR/MLKtl9ehLM3bmp3J7pt0jdhJ7ywRyBWx9u3Bw5dyx8Apa
hrZwx0ceOUrZjM9OjFsQVbGD8yLoFAEge59c8OgX6GlHu0+SFZVa6QKRvNZxGwlKNjDU1PeaS3JE
CNvBmGIcIUTFUokTlBCf9gujZjmqtr3/E9/yL8DRZPyW2V3psBmnDsDWrQs3oLJMS/9u0YEe1FJ1
hGss3GpY/6acf/ayI19lDXl2Bjg0r4O6cGezuth1yCACf5eY9p/WqrpuV9UBwl/FZIApi7m2OiHN
qrnbNlunyKYC7kEAdcbjqycoYr+BlmtXLasspj10NCK6AdLGUIkPBqzTkOxxkD5MsY2I6Kt0MgJv
5cW01NvohSf7StL3HW/fWbhlGMDUtIw2qhZ6q0QN8/F7Dp78nAVOjwAvfjr0eS06+br0/v+pgmrL
P6Vyx+vr4XahXKtWVOi+FXsZBHz0NaQrcXYfqaFYHYwH0wky11btW/hv6DhMmeF5TCqSV3fAOZF/
Xn2Bfgx+y/LXuWVOBC5YK7U9/zwaJyZblKc6dMwD4q4MraJNlQyqJmY8z2AtCBcm68tHce8MsmMq
GtbE5vEgxw9TpMvYrPUfHJi1XVsEm1O7sSgrCgbhV+aQuKe4Sl7zme4AvQ96Y4fZSllGqzj0dpCj
u1L9jUelRJ31KR3AAXouiLuKyMQnY3SXstpiFJ/0brAYfjYIaHTqCVOn0zJPOm7Z53ZPTvYE576J
PvvfseAOKiAy0kQpdexM5w6LP56ACH2Qb0mvtR8aBya/zOK9f8BxT4bO+e8IGs2NWUG2SHgS0uSM
Q0JR3YWTCBE0kqmhgajpTqkQragYqDQ/EhU903esNlcdd00EWNE9fmBOKm2af/JYuUdPk31UCd38
zNVAbPW7B5gOHWq9kTTMyvSx4q1c46fZin59O4BOcAzj28SmkUEpqK96eJZk3Jv1C2K+eDCu0EWq
04vnZZS7FBYztI3YLRAMbGqcUJueJvuHSZILHon59/t/BX+8AicgLnA7YHWgDlJx1NDssKtBS3Bx
C3ZqbGFBeFHrwdKTkCiMndyg3LErK2wjNz6HO/v2KxBy+U3Lx2p0+SFBk1JQmfIlyfaYSEoARo9j
jpVJEmWtZ4bM1javVevuL6phEZFOV73RsfPLAVkn3PvZXjzisqq1NLIYaAqEpXjEdB+UK1aGeYy8
cKPa/aaR78dzOWPON5GLpEeWX/wBtAJfYwH3oLHahbd0PId72NJpikWR7qoyk0LFZjmnM1CILLry
PA7COm+j/Uk4pQKz5tnj6dXHO/aQQtAyAeEH2PLS+zdkpwVEdHlWKYKBSshC43Q/wCuIz2hWQC7d
XMhf0wBrRizTsX1xabmURquLMNyi53pHX/Tfs2KT++i4tEiRJIyfifkFCrxbg4XwvOx+N4y6umIP
qrl8TXHPTBfmXq6SP43LUiWmoSd/VL82zSqLHwAPvp8QnFfG10xLrzNtE+wdZCHzkXkS+1z8hLVX
7WySP2TsNV5SfiDlOfGTgdAEQ+MccMjnbHWYnEjLKbhjdjaSwVh2bTNIr2ddfGKFuhzaRNsF7hk2
jakh+ZgO5gsj1sfrhoCLGRUlLxctUlZnSixP7Sq1QZdclBHDbcr3H0JJuXyxB5F0PsZDhYvKLmuK
EqhLumt10fZ70s/3WXuCwqi6AyFKRJtwtn00GlE+wI+LCmlvJKj8YxUTdC/6iOXJdYdesbaUIv9f
fYKw+LLfMG8E26ENlOd07BGKv6sKA9bIGzCJuMr0DdYGyX99JLhYOSDARtXh/GIopQMKTL6V3Hb4
diPZMftqqXBehFYuhx7YCzTUTHn+qLCEfFaayGgH/4PbMvcXYmdC9GCFiAhzSrWcDndbHnXAzecr
ppyCcaxh3bHkGBzDZ5Ux7H0cRxDto+qXvpNliWczhK+9lC/s4Y5+LYyRF1KRa4fXewKqObPkxVxe
aHwSgGZhFNwUyw27Ru7ORBzViQlFPKhiUH1PjsZj5bfjnQvOXKjW4ZKAbEwLtQsWX7r7G8AoP1Ug
oysygr/KDgtlxoMlW2FkhuqDTQaLmsnr3UFcCB6kXTmxSCTtszpD+In8KXrd5DsMzfHqulFOviGy
6nQZFn7PsTvmXp+VB4nUVf3bcHjmd7UynBvmGd9D/kzCTmpddCVAG5i1LENPXllQpJvvnv9WanSU
1rXGPpiRm+RvPY92K7wRhPBTFX+a0cFrWlJFqgX+0huOwOdCPUxyzENl9t7m7mtlqIFHwdoREYga
dju4jfUf74qLjFq4VtcaWS6Q0uEtX244SlTY6HDAxPan2rnfj/vBa0CNofR7Wkt+e0biWMnW8xJ4
fTjj9CrCNivLuNciHV5QpT/ZC8STGUtWmZ6W745OFgWceNT6sm5AAf45+DIt0kIfnJ89bUs/OQKL
LqnfYvXHtaJrzwSNh8Q12N7UllXPm8H9+bS/SF7RHZuVKHfL23r+LsNp7VxuF4wFEgsELZg4AI7i
2NbI5ejMJ0U72F2vEoP3mTuobI/TqTl83uOhG36gOgMzv9HvUIMD3PBKqv7omgYcS6hNpJtK8j3r
rDCLRAiskV5qRpPrFfo/rjs7sC1KdJQ2Zahi9KkpkCRq1Z6FnyVVDAxIqo7UB3EwmmaO7TVe5+8+
hTMcZT9xCE972tlk4+1BU5ye+3Rmw4/PGOh9qMv2DAcWjF/8lfp3xsnisZ3+YAo4nQHq/hW7nVL+
706QTBgAfrVyQ2vMfLrsYrcsr8pn6bQYdBGyZAfAvrnbnDlMA24QLCEAU17Zau/FXsxQIzmnOAjL
7Qi2msS4pLNhcuepY08TnNSmqYVl2mBk/pLv3nL9+uifLbrnmxxxGJC6gEtShn/qEIy6gbF/4b89
YI6Ary+gdUhYWTuNHqInqtFZBMMJA7lPCSRryukLMSh4kgGneHAIVgh9PGZwHHXAt7n6NP8+tP5f
R/9Eh31z0LhYqsEoveAcPUxwzuQd1QrwFIvZCekutOxcZ2wcH5QvzUFlBLTqg165ScLpMtfwYu+Y
IRZwABH6UG7mCqrxg/Zbd6TBwGoB8qZ6TjOnmSTmwSW9Fvg70Ho9ScKbaLHesCW9Wo9CnlAKyy9s
lDsYnEBW9hQ8eNH7NGZ/43lgkly7ZIfimSrzlIelAtlaAp5WVNrPfqZZTJE0M/bbbJXzwvByv2mg
FQFC6ThFkzC2eAigmi1g7FGEyDxh0diYUFyUHXqUWLygw+vJjjcSpskARmHxwj7x0oxzIvLtLGhd
uv8W7UuFn224MImrVRmQ6MHotzOWMIVxl2aa7ExomH12zvrW0dvv5zi4ZHGRSn0J/hqLcwAS5UGA
nLSAYvZq6LYEkl2Bz283AdKTFkEF6vv+gFDZWvnU9SRKp1XNu8I8QBdcKTphDkKRKFA29nHgxqS2
gROGamXuH8hqQAjiGtjSbr0kV5+7RlqIVwV10i2A8W0eJmai0YcBGw1ZpgR12C/KL9llrd+8qAy+
isYucQva7q2MKwqvqt+5+uIU5xkoMBQf88C837BF0HXMXnZ3Wz2vhX3xI80ZVUD+Jr1X1sZsjiuT
1qgd3dpCZFrBxtF6KK0OsAlgwcAIe6TCMCLGg/TuIkMEZ+Zp3tKmVFe1QJskGIdjmvdmDDAy6oQZ
clbQVsHM5qVPDczk/d89w2qIop7ZOxzlY2vzAovyOtoL8aSwpOhNRE04sSAjWgyf5I7AHXkDO7gZ
3Fi5Ckxg23rhsX4Hnws2qDNr0Ryok+1RqCbHEGFou3/YsngPGW8Vep3limi6uhDWQVBx2fqpvoBb
sdUpSnqTmxki6tKhMajjm5LG4toMsz5zP5N/5PdFIiFmv0Aqwt0f8n/dgtTO1hdTrhF98K606FRj
1Q/lnlEFItU9QtMycew+E+I6/uNLWP6sQOl9r7UJgHDu8jug9fu8VzKOxbcttA0aszR3aG7PyZ7m
ZItAJ62y0ulPawNkp/B+18ObSl9FHOfDCb72Rc1XK7wMKE3u+s+rwDBmkWpKyuoqVDgtyjd2AUu0
KzF9g2u/HtSFT1mVLV50YhUvAxlVL0kq6iwe9xRFsunteZL4SFxjlxhHCDMkzlo1cKPy6Z4ef65I
ZfUIW3Lve2FXeL3OhrtsObgEGM6MFKnPHymIFFH7CQpgKBj0q0vP6onJvg2lEMTRdy3YRXY3n8RM
bxnmUJXNCJJVEEydO7MuJUhI5ES+jfhbcy+98skygeFHPkQOSkV9uoPLEjpheAhtFiVORxEdhAfB
JfSzXEyJ9w9zYztwdOz0qCuo09rzzaUcnPghpCPdUybczsalS6mfAxkh8hjK85AdcXpB5IVj2pUu
O7sGM7DZFu/JKb0H+Hyu+tdBSqJx97CS3rV1XepUEvjtcomv3fZ7oq7GrvcQAIljMAjVPTXsL+xT
rMck/eBjLwzcpP7xlltBPBfIZ+Hrt5w3H3Lr2K5QhlsjNebFUiOm6bLAUQYcSyeoWxE5Bg+xEbQl
bZrIJNGG114FM+q/CnKzoodwTYwZRHnfzL3eV8Rbd7GSF8yXiZhhIxRy4iuHlgzKsqLFKGfVEpR2
wal9DHBGDmwjL5JGhYucieBXtEyAlloMZdg61SfMrSb3H/8s4cyT5SgSmxkT9VytdbaxCq+HHXO9
4g/D3c91IDoGfOho5aTvXstV+EX+7UWbjS1VtEPmwD++BrHAosC16kOo9ci/AfgUrxvZ6ixw0oiw
E/d2vVNuMlmVT9tbXzUJvODwouaBtOOXQ0+S4yztQKTr3yYTxBfUs3/sFKvMpOy6eVNxSIRIClNA
uA/Tzv5BrteVHMySWn5X8fGqWOi0RlnfK4R7sy4A9TwDh7LwQ2dF4KK5pwzIHX2q52W2ymKtJa6y
0fevHDbeSD9OAmWq7ZtgeN9s8SFDVVvkHqOLNOUQ/MTyjtUXx1PwYf1JPYFAzapKHIrC5WmgV4eE
yZx2aE408T8N69AL1Hfn1LVqXgu7v+ZTYjK9Kcs4Vu8+GNd/eZXuX3YQtAOPFxlt964sgOdPUriB
qBfBNdwiNL2LYhIzKVvI/BDeS83CXOYG8HBOr6pf27EcX1lAJyKj/5zzGo3pKbPQeqvlbI7lSJAs
MM7iyu1J0bTUIUrLgzDuuILrm1dCStBFYMnotRUrBG/+qrPKk/HidKuoK3668xAucnrgGuuzg6mH
ypFlEVltmPHK+C/Zb4N+mtRbqx/7oljg1yMO5GApTi4s2IWDK+Bdasm98fHMZL2n7gk/1TFGeanS
WUzJsog3wUsYYzGLT64KL0kbt1lxRVIJIVvp2cF+KUvuyCBIkXLN5xk1FYPMB/9ZPkiKEyCTCh9S
O6T5Al8JUil+/s4Gg+dvQCYyXEVghvgkACLQDvvyJE6SYbTfa7slSrVxqhpsY4+cw683uSknBkLa
nXBRcelimzyqvqX1kBB1JY8DXWweILcZoNwjL8AnjRjFHLTcN3eh9/87WuzcPjQ53nzOFVq1mwLY
qkoLXuJWoKnUb1t1RoZLl506HcjWqmt6UqKLlI+4qvCUMRoi7SrgQ/ykT7agESg83jx9ZM2seoOV
LcbNjpevaqQQawlFzTifmKgkMVSpsjDX4lqJm5SOW2mJoHFqXd+wSjhBltdvs+DH8DStGXLFjr3d
QDQafmzFhFDATJXa7Yz0CrySBVGkvnn6hJsClO2w/Yd4846kWg4qaxe3YtlQaocB/zAvba3D/Pep
kV9UeI7UrelYnDxRKOh8524u/G4bf7k0KvjdwjzJPVfDKjDwtRmQVxirYbl/Kf0uTXGr4KmOfNr6
ELJYRacZtLqqrYr4K6XdVUFUF36Xj2lTvCvx8dFBsSok6DwYaocLd4qvnndUbYP3pGaGIn++TtYu
BjfaRdp+wqDz2X0M0wvK3GLliWK0noQQhK701T2v/yC02J0QLWa2iXSKq1p4wRzWYyA9PtLfT6iv
9exV/ncLd76L72unk2b3qxFnOCYetHH77vVrF5JdhMjA40vH6m6/vfXBm64iFsMo4jEhzR2MP+4h
gE5p1ReyVgfJg6OwOZUn+DL4VaDvO71sy7YJo7ck0cXq7bwnv0EsbYrB4hRPVivzeiaBz6CGg6D0
F7W9nZS3DNDnoB8JXLIecGnMcBNoRQcnC2kkD1spFaAIEYDU+OO8hgvL1sthuPaNYHVjxfV+TUHr
Itsb05/NQeadDisuCj3iF75phiol88NJZI/zwIe3neqxq5ErZqjoAcJIBdRhrwdW48BeaSVvptD+
1Mj8dNd+O0Ko1OwzcbZcmEK7NNXSDRG9cl3optOaqCBmMAAJNn37KxO9TTUsVJLJp+Kq5laHp6t6
7GcJq1305aa2T9+Yfempfu5X+CXHKcZzedhZL95cY+YdyaOMq2PtTeSQ7aBREKNT0Vy1UhMUdkul
B8ZaKJumCcRTKbEER0dBrxPQOWUvT0td0vIV3qGEGlpIeVpLnwawYk6xbb3uPDzq+vMkxtPuVhCA
GLCqY+yqyEmxbVKd49zM2RFrhee3Ulg65ynPuAM4RaXt+6mDVVZQuVFLJg2H4VpqS3NEIDO/nkHd
DxYyiRzGHLmvP+FSzvHtzIiAcVc7qv/oclJWS4QbLYQve86avKwsb14c6OXlz8EuwaImGak3sG2D
3hN0j/dOvxwLe66SAl2hbIGF7NmLEsozQrKc3aWB7+e9sy5a+jHFZQtto4WvaAzy6Rf12cx+2uyE
1WXdtUYuVmNtR4JU8NatXEp7xFUlVBAVttiSHtT36xIG3sxYFc3mhy7VvxqTJvarc95ypQGoO1+S
aKpmsguUM2+9xiLkbP65eOd4nCjWJQyt/svMVHoFle1U4f4g2RkihDxsP24MTVvO6CR+wbH0a/iQ
/d45YoC0wAiD7KtLoWimwGRPPvr7OYiN/eSfLpKNu/1PP0tehuYrkKqmq5RiZR/rhpaL3rxpDdUP
i0AljPjdQyaE3dcOYprUh3VyGbISeAaAyO9s10gsd7uBK8RRtZ4S0MQmwQBIjAOAX7jicNn6Mtqa
VhGq1vH0Jn95eqg04W2wO0AkcypPUgCrYZtOEa6+QNMHr0rprM/jvo2msk1fmGTxfxA2l8PGvB/P
sHFJ+YqZOzgg3PQAWYz/NQIW8ma9Vk3DPp8PWFyhrvOiIhaOeCOA5LWOMBh233WLiFO1C6R8H0LB
nzi+QB0WE76olzlA9UrJBxVQkK9U9V2u0VbKRPeWoA+07sb8ih0U0Okvk+s9zY/0qg3t5PNuYbTH
wA6tCxZp5foZFDRfihrNr9WmAmmYx/9yh1ydYbL1hMLOWcdA1yrxov252GJsMosDHhD01ar40Zji
o3IXm18YlG8Dnhb4bCvc6SHJl/lxf1RQ3Qnb+AKqFgOPKKl9nsq7Zk42eHtNsZIa3QrItJQITYfB
lG0FTnWI12wO4l6WJOEwa+yzDms3bRwBNAixsGZgFhHnsN4aGxBOPHhHxIJSJwcf4Nv4UyPwy6Hr
fglcbQHhpqXhsDNOtXOoCOeeOGK0XvSBVBG75HhJcIHvFH4/WYuyw6FmHRzEsGxKvscBnJwYxUHO
MPuvPWykorH5z9QGjyMs/6ZU/Cv7RRMFiY16vN2wPvTrwGUJ2glO8XMxjTqGu+aono6UwOPdGylW
34JkTMj3Tmefik0AUfz1XWd9rIYAU/QAM6sgh2BbucXLagikv48lrAXT7OjvyxjFqQhrEUKT6D3B
4/ai5mJUtfbI53T+MdqfliAHEXOYYxuNqWiB6KYJ/ziPiYb8T8fCXB9gpIT2+ZcaoTHWP6zjzy0a
XUiu+Yz/wLEUbY9ZumT+PAFpIM27Sma93M3xEaot9tD74mLcyTj1gYVNHOAgI17L/unpGM6E1APh
Nog+q2wJfaUwMwjZ1HRq6DcVd4bCkG4cjinQtn/RtUPWEO7uR8audsXYNqFKr7Vvk9m+V3OMNS3h
75aHVak/lMILiGHj0Z9pgEF1GfhpumDDbAHKiWIbGW1JcjsXnNRUPCpeJ0UdGuoOxQmbd0TzQyTE
GBvxFlGpdc8XTIMoNB2BHPSr3elYKqt2l7OsKDaYvfz1nT2DZ1K9pRKqUYu8k07lKR2L0f3b11EF
3QMmzE1y1l3RnrgEZ42tPaXiTUIZczbEUIB08YVuLmdZyfP/8uGNtHRe4Ca6S+4HIHlv6flAuIsX
EL3ZvDENV5oWWDGKgMKFwxkQyqp0LEcmpgTJ1fVeSt3MwnBNP7t0b5sf5CkB0qSZIBFpWY6QOB89
DEdp9LRikMJJ3YdCyiIe1t7JacZH9nmLKt1kvKnFDPqs4TFoMibovKl9D/NGSAWJLKgoEJ2PoDc/
3YPLU17p8PpftU4fqLBqKkzpmu69wYdFnC2W9Iw+T+NmMtYNNMT4kzb/ADby7ucguezuusRiWV3p
6GFUHaCHsKRUayR/AUt4WespZCyRiEWynnlM5x4mfaunsVALP8OwOTWIWLx6mDfz/zv6/H4ZE5Vc
mLl+Jf1z1jLPONb7ZwzDZ2rqm7+zb9D7hnNmUtzHy9IP9sYMpk5qMJubNgRAsZDjE74FnXTlB7PG
Eq/HSLswX/zept1W9Az3H+XNmZKVHvGn7DPL8GSSh2fG+vdInySyeEjY48Vqlh1Y4bfUuQQB4llv
pRrA4EvhqCGaLr1Gwly2C9Ve1zBAgtAk4NVcQuh1Ao2eHrrE1ig+HTwdRGqGCkUC/6eJHoclltoM
LFUHkI/AAOtPOCOTRWUe63EqUXucKcKKFGK7M+zUxhlPNARYxHP0sc3ONRJQPjlB8Z2m4h5kYES/
Rgx6gTrZpFw7DBth4tu46jdFmDL78oKmdkJ0nfYBM7Wf+gF45juW5tkbS/7NaPgJqCNiyNq1VZsQ
2w6S4/mH03OmS2VbTIxJPF5TrsRdDXyEbxBcijjiOobseHWf35EOEfzMwQyYnm22Gc1uJzAR5qCl
ZPeSBBF09tk4IbHyfjInQDn0GX2dCkHMlXRqENtkDTziviMdRc9jHEQzzS8swVf12cM1aYxFQ281
yBAW6b4yH3TF1/oGNlEG+RGrFuWZBbyFCVDjxDO2kQlrfYz2KhMFkHxbD7lrZUSqJdb4DKF6AytG
qq9fpM6IxO3byBCF4sdr9Is/PtiZnQoCaho+dS+EbJrsHt2vSwPjAIvpTsSqOOtEkihOi+Xpssvm
15a7PJ9R1I066g79Bu2K7MpOKVJ+462nw7S0qMo80KvlKSellQTRmtEaDzDf7ACvrqN25O3kjLVM
hCngNUlpWvfJ098B5PzURaKqQ83k7eDgy02wd3GFh/Q1CTkaFTROpLJ5fY+2zqTcykjEXmi/E3cR
rQemDg3KhqGYxqBhDLMhI1PLcu0L+xeGjvhE5GW137mvlTzWAwS1PFAAaw7JPKx/BDLaOtFXArhA
7d/7Itp4V28FQfzKJjm/joxTD2SjtMDdqZKJy4OLjFMESlksq1PLthcBNq9XKD0kZ2lbfPcRGWSe
htQrM5BA5ftPJzyfd6i2eklizayG4K9fy7ODpJ5C81Bw3RC/FjWN996YPL51C93/MXF8oiiTPd4r
pUZsg6L1QzSpv8Lj8QpCewqgJFN5w55iYQhAPMKEeLnDXRxViivUyLe8FB7ssoX+Em6plb8KeJUb
NIwYMtlYXKx/Gs7enZZzRo3rD9ZAzhrDfG9BdX1sR6qrLojzvJMfOkQfkfdcGuPgjWF4xS0BzMrZ
wuY+glSO6iqnZlfURHlmVNQY1WwR3jI2r2WAtzKfzFDQLrEUlv/Q+rQkcIXRyAm4Gx5sCw53yGik
2erOPxqceY3KbKFp6hXZFQOAl64jz3jIOV7g+5BwFpK1ohA6xmJFfKZAZQJK8eOOo4wokRBKYl/G
/yvfR9SgtZ9EHxpZ5uZxqWGAORU8/rfdOSl3riMFmE8blFlf0l/agdWW9P58uPjYfadQQQ6qP8hf
1nQg+GJGr+YRsXXM/nZCnKtGSK42FSiLrcmbxfpJGPSkUKWeBWSflOCvuQOUVq9W9hmdleOloTE7
OTflmRzp+CpUmp3yMhdW35zuzsjUu0qWyabMry4q6Hwts/ZhWfQUhfUYlf5EKrp5pItWETppMSgZ
XHMHKRxy30noZxzOQ7/FQJzMugKb2wHRSHBvaHL/fzlZlM81c8IVhvw3toU6ymWzJggp8LaHVAIM
5B6LfrjYGdWQZTe3A+Q18K1hPKYJFDAcoNc5JZX8TEYrLbU99ZyPC6TA+6i6pHFYXBZ547HWDsMV
rbwBTDo96S2mv6gmXvqomsH2lfujxqPLZvshcrmv8Gf+mJU5Nq9mDrYFXRR3tz0SQ3CVXJaYfHKY
LllNlcNMHKvWWOBt734woXmkVHmDrlVcYMgqTNbVYaNlDpiIzUbJ4AtYDuOVMt1Lu9AmAN+35gi0
H1X0j0F2j29gjdyGa3BbVgf/+J02peP5OtrCvRjmkxzig7hE19GiZLlfeUD+rDsygF27biD6seww
xpcx8eZZv4viQQlc0a3pxzZmbS2Dl6AY4Yj620wNhvN5wCel+0pYrxrmXBflZax4Hf8kDrtig+4I
EMSrAqVoSx0xsmsEaqjdmrhMdiFGka2C/Al0WREAZWU+yeWz7NoUy51h290IRwEXSHpvFePAiw5Z
6oslNehXx9TE1jqY8syEsMvkb1Ma0OvqtwzU0NiH/HEG0xAbSeJj9/NvIvY9+oSCrw6og9RRqWlI
5XS+8GcW5ZTFfJP3S648SVSAywFMFvXHR79R/sXe/UBElrT3lKXM7npNXbRH0T1RanL6jI6mEziX
AflBiLcO9fBWQ2rH+sAJuwtknM9Ye9XnU1zofAljTsEAXuo2MhCq+I7fLdMVKLmVhm303MpbhXn1
rcJGA11lc0JwxckqNqFa4gCLGWZk2XyCZ2yTlNiXzfi6L+8laBw5N+EwLdxCkRhH0nmBzWq7YK/Z
9kgdZ8FoVAWG/R2gISR2ljPFgCJn1rHWs20buhBf4Hr+nKnH8tb5fSvSn0e5ZLOjbXH/LgBs9eio
0mQfStGxrRj5usROacWXmz+ZeomKGjaiNJuOrXrmzP+FZ6Th995YRdGk8Et+Y5VJnC2jNdsnZTTU
oJsacW3zitp9rcjNT7bCajkv0o/ClH6hHED0JB+uChetebaQoWvJcLYkeMPZSY204838z2CY8ItT
4TK41XVkDhWG3ITkazV25r//pV6aJ1OXM3Zy91J9Non1T7ESnfsmFVR1zHuh4Jwbs+jdd/acbuSO
rbLhEpHiqS2+s4NcDSinj4PFixcsnl2O/urwIfuH8huNXTNrY+58YXsDnuISWiG0xzcONea0opjk
x0+RiYxx/pMpu/bCAL2uyVL/8Ada2mniCWJoaaM9qoJtJsjHlz0Oi2Wm9S8cTK1YAizYxyood/qZ
5RVclpQY3R7OrVx1zUUStOy0ROnoACBmsyB1aIjv5/RhpPsvSSisOIMxz20Z1j2Mg6NcuqfULHoM
TjTjUn2dkCpe8S1MgQldQu67r0qmlbYR1sRHwqKImjKmUmkyHmLQ0EPNwZSLfXr6gMYMj2NjdAIl
knhe48NZ6fCpc1feWzWM95qubEWMmtMHLIVAIJcmJwVP4UJGexIZYsNhkCMhNJ5VASgsg8PPZOC+
Jf7SFq67mAWW//xnDW1H+idbBPAX6r6U+PeumALV5AR4e9jY3iOg77+zLCEVoKu5GoSQ+e8GkA7/
1FjaoE9KhUR63jtVPAdviMvlywdnWrTG+9nUvdWGix4z7w9mI+3hBwYwgfhXDoOarD3Kpch+ebpD
7snZXiPrKvR1HVXZWxyhvK68Iz5qLNjFoYnjyYTnpHCo5bajc6IF28gWPJMaxzE9HwfyMGC4CI/9
m53zUK+NDwpDUh7wBpAKJsiBKxf1rrDbREr3XOUVDBbbcByoUmke+5kaq8H6Wso5Ghc840spKLZE
nfM0q3DHN5RvS2nJcsynl+lGXCy/RWquGRsb5NJiS2o4ZfsrHIRkyPE2usDBYl2eaGmrSOHGNI6Z
MVKbOmVsU0XL5GQxsT+bmiVWYlifTXSbfBifnIfFf7BM9h97PWe62zMPXMzZDe2yOt1QCftyoWNb
ihQuYg4iqKad1eNzevmMmTI9ZSsiZGqhvgrVp6S8TzrSNYrk6NLZ7XvO3pm8OsQ92TJ36KqxXCXH
uxxAPlG28SvuJeig0yP1SwTQN7mSgj0u9FcVp1tlT1fmnZHHVR7ofhinQZHGAYzy6WyAK90YCq6/
fuIRdQ+SgyMI0ZXOvkDGTECC02qLnguyJxuPigWD3hx1shaRD9BpuDVroL3fXaptaR8lE2aQB97t
pBMddXkTXzl//bI/qgL9613h5RHjyMFT/oA56UuXqKfi0Yxr96NiWmRSxdn0BdwgXjawzs8Unjiz
LFKspLDoERREco4jbhgZcTAZ//yLHw0YDCUOU31Uc4hREL5Q1xJbO9KqlNmJ7rxyqlRss3okyYxY
0zwQ9/GxzbifXQzbTbhU/y8YYR0NZuRC3aDm+sssSrFYn0mQB+W7w699xL7f4yf6z62iBZw9lsYo
scO1LyUAPZn1w/QcpFnS/3Dgkqmw89KfplzfbYG7PBCwIMbuOeiW6hLVkEy14NqdGZOXdq+puRKi
8rESb4pYovZNeoAnhvNcYGwA+4WQpyKabGpGZ+e3kub174GTy5TIu/waFhaCocj7gKCcxU4GlfoA
TLyOaZC2aI1WB10QyypShq1tYgheCDn+6OkT30E4j2fTqNmsu3vb341L2ljTITJFOJiK0MUvbMj9
y7aLt+deSzWFoMJwInD+VK3H9Ua5ieeZUBWeOYgLSy+LRg/8krSlyOdbm4hXnnU5HWk0E/ssfTPF
eAy6WRpmz43QXcXyu2c8grtagSmxmgF6CgjeL9C6rUnRcDjgE7LeY3MTSI1fMUCK9ye5muejtenc
6nCKR/o5VQbzHRmMTQPytZh6v3P98rzFLESy6xJmmmkhrCArL2VNRg/hJDXdmccwNl65O28ije97
WWGXVm5GwPGTqxpoxNqwZtkaxHBq6tlAthZGkNgs1R2aUAC2dhT1wgQcoADnR8IqZVuu08lLQLfD
m3RDCMN4wLQYOyH1MltZrxsWGkoTbjLncA7hXKlxmaONz5lmw2+2tTdLsDZhexdioz0Z/tpzWWvb
YDn31aapERbW3HINYReG540LyRXEArnC369RyenT3eaJJZNYHDHrufqQjgisH9ZgZhXLcK2yP0Rt
bFO3OvvQ4UeDZRRDt3xB/lKXTsMMOxNZRxirN+ZPw8EwKphENF7ezi6O+JRukGAyzbzjJMZr9Hkp
ktog2Rp5i+OQHuViWaJtoqZKxKe0rAgp2uStHMxrlSf15iXVIuu0KmVW9luMBOFWk9i03/2GP+dX
HP2tmjGYJutjjLQB1nT4WjJXufWwB1QDTdXK+vtJUXQKKVX0ctgneYdV2beOApY52BN6F9gmGkE7
RKadeK6FgPn3pTzGVMmRHCNFIX8cYx2wNKzDqRW6Xs5h9Q0QPinNJ0bLWrLUL546oDsMsRtOrFJZ
A7kykRVMG7mCGqVXCq1TqDogHyt8Aijvl+zCVec4DRP6XO+lxi1lbAb31zplTqTW56tPEpu5L1PR
aB/YSO6X0P/f83yBLy+3fGCXENx0cPLjYt/w2q1Ar2ZGu3dHojPuDp+lziuuCK3QrW2GrHt77SQ2
M3Aw0vFlf5fMCoNf3pEiHx733r5yvFc8guCHY/8YRMDLSLN4k1WaKb6IX33p5uOSXWyMocguS2WE
RGTHYmBxa7d5e+fePwIAkAGUv8P9oh9N4Kv2A4DKiEZZ5pSev3ly4hFJBkqatijK+xtNW3lkv/Yk
XweFkEpZyQEUf3FKuxh9J4YtOEszmljbTSNSeIus1CnsqE4q4vWYTf+K5aRnUNIUaFQBHegQZzYV
0zWiyJM9oGCgfW07/6HCrxpKAInD6vLd1CP8PuQ/NYGLufaxH8MHIbxa+Q2zK6O3E60DECyX7lb6
c1wwz4iNlNZmFGqPfU5ORMPR0P5vy7B41eCSMrtDZzk9/IQ08Z0SgGw/xtv40XwVSknYB4EwDqE+
ZndrGIxhIJ/y5E7b885KTimLTRlovU5pcJ+OPmrvnUk4NB1EJlgUWAirSbK2SpNWkJBOJ5H+Wylg
rTZMuTePpaMEsKaoYk2ew4DIEIaQGC5dJ7kiBVtzcrBDTTb0WkjajxMUo+TppSV8PZYDwUKKb0lf
KyOR9avkD4doie9xlpXHbq6NbLmQBk+6GPWdgXIBfQcIHgfCRLaNelVD02/s0ugbeK5Jcwa/UM5F
Ii+9/hIi/SIEuKNE5ROGLnWE3fpPvF+XGjveTy/jYcvZ/XXtNY72QGmdIGdwIJgPAfqTQ9iPROhE
X4qfwm8hMK+tV/aidylSWHCoi//3zoE17ev633Hu9M5jcG6lXsogQl53MhOaj5Z79tfQ0i4E2zgJ
Y+yxll8/K3aeIFgg8TUhjcDcjx1z54kXO6I/VbCIj5Fvhd9IqfXFi4XKZWEVdILd9E2eblr9LMpb
GgUShwD7bPWAbUrPqd6n7AAl+Z8BUJddLS2qd6CrFdEnFr/8QNl3GzfS6eFho+s2Yx4mFRL036yC
3lu1edCOGfpKnB2AcsaSJD0BQmCvhE7q0iEFCx9sh81ys7OOzInIl8Q9zWHuXOxjAgru2L4ufyXu
m3Ab2VjsCjnLq3JIp9lDKTU3RKqBf8181XXzZdLhsW0Gj6ki52OJcgrmdNJ9H1fCTRuP4cqZDrOy
A0kTVytIBsyhWa0Da0ca+8ndQoO9bl+n+H7IT1+xf2j5ciAAeCArIgkbOHm9h50aPffhNK/rUhEC
oMJDbxobwPK88fsEj8LIAXpkxsMB9OfSQ0ZjHcF2k54nUbOUr8KtorgFaqBILY2XmrONPr4UG3ZQ
gi6pGQglybjGLMV/645jlpo8m+W4hPH6odoMc6Br9QRcKMEZjg0xxIZGLVZk1uqEzeJStMtcBM3f
+e7JO6mV3mYCvQPnV6nXhVtM047JdkURfZa8NPpz/pilWaYV+QLyAyswHsvbrcjwIZ4u68GwXr/1
wec6hB/ffmThc58dsa2bDhQsUma7zWVyr2awp+yKNY1RrVwZTiGHY8Lolv+OzMLyYgvzGv0IBpJf
Lvy3YWJcDvt3A7iqUYS3+n/zMyLapWm+lMT6Ua8AqsYpc4xoMoBe/U6vXA8Vbgg9J6myUQWEZivw
ZSPvLNfkWBH1V2IbmDx4gmoftvHeoppKX2uQZPnznBHH568tbhHotHmmX44OBMagbj6/48ifVmXJ
sq3tQ5Wf7h1hJ2zwuCXVMZs8GtJ6wWqanRkJQNE+J35JHk/WxJN50YL+rfvYC1Qdyfv4GL6IBzuU
gLVpHFP5aYX6dvGYdWkCkRyv/ABjL6sUkUux1ZWc5+qi/qf7gqSZRcpmg7sCbclqPvdYzLROuf6B
Le84vlfVMUcgo2T0lHbJadY96ieJ3B55gpZnWn8GRMu6xrOyBpCf/ePcQ4eHTcUALTfv70zRgeti
YRG66gejwhUgpvfEdzmiGtXUXkAd3LEeiMafBM17ivgXkoB7EiScjDxA3sYCaiCmuWNoovV0bjHW
5uObk2S7+Leic0z8qzu13sRGmjwFiHnKVhfOjk6WSe2CF2mr88aMxWhnU+4BajPgHLNv4CuR7gv1
TO3qDyzrOzgffWkFFjfCtlKlAqA0Cpo1icBuBrnj/p2SPmLkwWD1MO7b9ooNze9c/nUJVLTs6E78
rsmXT1qjRp66g4Su5SiBM+AIjlDV1KclMzs7jXOSg3GeC3QjjqgPobWiwImQolzKzU6m4BwqQJPg
ojMLMimVC+Vt2aK73qJqQFvRIcT6CxCZscpsRchTibG8IKkVjaD9b4UuZP8zPQLCZofJ8kkaejSR
b3jsi1J5MJRUNPmtPDXz+OLdlys6i33aspJubCoLj7s2iHn6p6FSPA1L5W9iArZvFZd1CZWnx1EP
X/2jD8Pdt5ubLo6WkmjTB6m0iwHDh4iOWOmJxEtKzHV1EkUIKAu/nvTK7CirdHLnpRN8kgy8rOGL
wCR5ccohFNNz5FUEFoCYD8tGgerpOsak8J545xrI2OkVns9y91dfWFqZsLkye9GrSkMuAgJtCL3y
KF6ybwAGnqY1lrNbyH7TYHoh/EPNSuX8u9ueWsOchiyVyU0WX3EHhY2YaDmzqzmgQ8aJErLFjkyp
7q/thUyvQajRT5dX8Ci/vi2lsjL1C779jOgL/Bme1HWRabTlZkUDQpqFVCBWcsNyUES+vU0zQXar
4mUkGwiZ9LA5a5tqVcCCp7Ev8UY2g4ZiYrRCOAYJRUE0oLlWGKLCnzqdtLTZjpFVSKD5jZVjAtmm
+IDBrVgo6VTZCpl3/rnXLlzNHa35vnPODJonTekJrjdAvSUXmBFRHyTKGGtxNCJ8AQ/5BWYpNQGe
5sWnDBoK1H1nglkw5OI1D61XJhB4+3CHmFp2ZadYNFUqQiKlcLrhKBG2n6oG0AydyZ7XpRvq3H+T
1LDd1/xcYf+u/gJQxzbbBujvfNQ73BQug9oixanWlWVhKP66wmvanNGSLWlPA/+41f7V7Cs9CSxj
ixRpSeZUK/Y7E+6g4J0jd3hdyT3xlNn6av50ZYecXWBafAy0CuH8QIOTgkMFg3l+F4TS9p2bGOFE
iJXQrNsoL7xiGUJhP2kz0Ukuw/iQSYjMGMjCp0fLrNZAceOdD9mhssJ6C0pOCbJzouJ8l2jmkyNr
88PyVmB+128C0Wf/x8HeJx1eWa1M+HfFacpAON9QYgUXneuV7PnfYLQBCd+Pnb6Krq6R1ggR3RaO
yYRpoBQVmbVoq3sZ602QlYGjTppO0PQEl/OMlz5Yby1ps1I+n7QqiIfaP/GCqnUCzrEPm/DG9UNT
iKxXXqJuVFTdEoAuY29iRfUbxUU+Q+uDLME4/8mkQX72q0JeZVdvS7LEj3bToU3xIPAZKq2DUWYt
rkohGsYgv0gd3s3u/PH5jfrNPcXcrJsTaMBcrTdaaEEqJJrV5oKahYVpHqgrtypDR7RJzNMnvD3u
BdA547eAJVMQKEzz77LkIHQb17Cwcecoa7k4keTjAlNO1UVMcGQU3DmjLBuhP6HcKnmcGbYA1DTq
/LVI1QEYlOpkJ9zwkNkJg6sXoYBGLeqMkhzIqaTLKWbPsQn/HeWWbPOyAgC2N5XPsx/ooIF7evvx
y8/4FcUg3rbjtkiKve6GHDOW3+0snFD/YJMLepJZhyGJ4f8/zCHhvgQlOWWvy67E6wAZc6rYmD6g
YHtJ1wOwFaZrijrge0mTaeuoCS/PQmqhpN+pO7wUXAXBVLn4LKECHQZ5S/LJNCilKrxJpclE36A0
rYF6F7WlGM0pPQ9rpsx2kImbOFMg2qJi+AJU1Y/H5wU3ttjyLFHF7rwWsDHsceiC3OQ+gOATrvyL
Y66HnVhIhs2UQ7fyed9HyecMaeUmYERQA0rmq0fjUKg/0ZbMhBlwRE4rgt0+6hL5lfutBuIAqSfZ
QFfGGzB8MdOvxza9gbawR7BiztG13sT9KuwaE1zOf51WyDN6jrQvsrH3BYWkzSahh25EqUkYRofp
7E0l3um/saPsg1ROKnUPlfysewPbwdpwZ7LcYXfMSxiIU7uaCaJffaiW8PHVxEm8wKpOhUWiqoMY
ZdXvpbmlltPDpvA51XYPRfUFyhS84FU9pEmi04k+9Jccwge2MVnHjtWI/dAihthPOW64A66ppBBn
41ecsXUuRaJxlHzJ6pyognGI92yNpRdZpmIKrSB1fCIra4qWlTaWJTxBhDGQi/9w+b2LfwdZGAaH
YNjk+naoEb1qTMQiLDPF1v4aTn8d1cIrdy8f1F8PG69va5BpQ1vXzlBucGhRhUv6BUD9sMGHXd1F
chrEQNd7vTSpNzWfM0Ba0ZUHerA9zbt1t+BtfTH3YYsPKNyHPCu362vuDW4oYHdFGGO0jzNxrPxT
6X+j9Qt4myjjCZu0JURHptPnlHYI3yRD1X2QZLXqj+yQ+hOt7Z8JJcKqMo4gzdlstV1Oj/L7+fAG
PxFQq9yfM7uZxaIq9HpCUoNQRbxIW1gzovvVAUs1WxyVtWN0gpGB3EZX2HXxkWH6siz17EaRPPRv
WGpgpnLqD4wh9rgOigryfd4reozF6jroc6gH4hpundR9kMy6uOtDTWftrmmWO5vm6pB49D5hwVwE
yMtGv5oGbVGD1IIZzUqTWYMl1HIYkiPCgDhfXgHb0BZKFyKdsl3q303shfajnntwkV+rOfQvMUvd
w6j6cACtle+Gw7NXmuiSXGdqTvnwD7wUIZoTT9TGjVd/N9GyF+x1nKKzpsOQZI3cgTx5PZn4XYPY
D7Twj6LZr+otveAzdV1M0pXor6owurZ3wOFIPWCwZrbPMq6VB6wwAU+SbOnNDdbq7P0DSYf4rWV2
bX+8tWt8GRRVHeRAdSABrSiiwVLU7P83liO6e05gzkQ8u1W2M0OZArF3RjvrYYAz9y1fRN6nS1EA
my9ucl+DUZtu7X1RYYsoEeT7O5d3cx1WOvTtxNEvlhsaC6CcMrnh4PNXnqZFDEyoH4mgBMh/lLSH
uCSkSDshbvI8RWZpQLOZDVhmrmzGWlN1EKFnKSDdO8A71fIKfQHJx0Ar/RKF2cYOIjLlb18veLre
85DLWVfDu4xpz+PQzZXiKan/zrJmbqGGOxABbNQzBLajy/ovNeEryQOp26mbtJsDH3ZywEgUTRJP
H3c8bBTruUvvM+i19MMANmh1yb/vYjWe3aQX7wvDMz1V8UiUrrbTD9I66ecFTrLYcxKmqsS+duFm
7ZNRWBISLAUN0bY8sO5mz5FhVGcFH3bbeivFboWP0F6VTupsNBs55RV1YP3er3+DLCae/l63zKtd
jPMcxkSfdsj4fELASZqjBJ4qajvOQDw42/oIRtyi5mnFVO0v53Ah0FOErYQ0Keznp+5qlME1+S/m
QxcQjkBs2rsnAEsdalmiMuzI4FmC7FcMzDka7rlLDHSonr5PnDAxTHw2DPg26Q5lmb/8w3LEP99R
ZY7VJeSWGTcS62x9Cxiy14o32UBcNrKV1+u5MUQ1otgal0YsAr4ABVDJTK50u94dkleGGNZmJhAI
fXmVdPyrqj2ZsbXDSbaigJva9JKesOJd8Y5pXkanHLlGU8FONuN9ihYTu8kZDU/WDCDFZd4ajinZ
2IYMQMxSlaJAFjOm2QxUi7i8d29ajcHUts8WdIQgViA2RynMTojLW0wUZvDGrsfEBAwLM1sdkc+P
jh5eM4+Kre3boIWWPQxwwG3KK/3Vrowi/hXiDg6a6wB/z+nc4DgB0dYpe5iPM/piF+HV0DKyQ8Zk
p/PgmFoLsH0F63MCctX6cZpFu2ZKDpk1NkNAApMLvuqYtZk9D9bzn0PLDGg3ylaLN59hCqCx+zSl
3GiTntXf1qFRLcenViowXHNwA4yEpkKi8ppdOizEhQIjwZPWnxVQnvikE5O8pDi/+2ac/w2kDOYT
lTU3OSsE1ZgxbHPjG7xMXSVwCWj31XOSleUsfGWIJZ1gRX7mnzhUYrcUHOth29TPxX8fD/okA9Xq
reEKAWZAGOaYR/rKc2kO+5J8T7ur7T8P85x0YZUF7r22Z4QtgQiH14hNGjdNcylACvhgWL8vk6Ze
8klRnbBNHtpQk4LjEKZG95FmKKplkSatdtRCMhR5EocrpOwywlbNaDCTT1WQGVWOQnFrtallwfhD
2ifHKSuzSSyJvmtZmiqsnITGmZiZ63z4e/z1uC1mJJiJuuwd9Nege1KPDR23ZRtg/scxMkU7Iel5
jr16w3QCOox+EVrhhmE1gjjoRmZ49SFjdybClM/Sv8l+iYmVDJs+cRwNdTKiuftoO0Vn7K41l3Z9
QzxGww13sIPVNmANSKCjE8BmpvpDClVh+0mKHmDZJ4qzcZf0/1IctV2c/A9ivRL0xUntxEfIgQOL
KxF4L5faEeDmRtVfh7WPYxdjYfTnqXcn6GiG/sBe7GzdWjQZUP03Po6m4XnaW5idwNeuqMluCgJY
7o5JBxyFSQs4cfquVEzkKdDScKtLkcX0qZ5m/7tT+yA3pbUSeZM5IHXrHHp55be5Vjj9OYNTR7Xf
d035U+Q2G226/7abjaVOrA2wAeKdmqJUZE3JTQN0ehe3KSLpL6nnFjN/Z9O5QtARDU04pWBtEfkH
NrYegeGrubfYxDTXS5jqEuAiy7dV0qDwRZLlrf6TwADbcrEG/ROh+YgUANFLmGScZXhIuQ1Bh5l0
qE0g30l1OO3tc4WnuShP5VY9OvQ4ggC2MS6NvNBPR1wax1GYMNxcfShAzZPL7V8TpmsSyuWLxQ8Q
p6BR0OY1vjbSrgqCxkGiU+L0sNJQ6AtbTK/ywfI3iFg7RLAlUXHoAn4IBDHCakIzX/sCa55WdKaG
zJ7/TJQXhI2yqf+bnWu99hGZC1a6H6sP7O1S6V6DpEm4YN+QejsalUVzlDDgv4XD3TggSpcRujOB
IgKAB4C9vXZE8X9Jdm0zGJCZgy1W/kh4SvDnviHf8h6eRZZCtH5ujY4YmASrSqVLSkQE7RT2I8vP
9hVWyuERWo8/37V9jOGU4dIEB/cF2ZvfX9pSI/GulBBlN4R+IRrigXqzLIF1uySnskUwB5/dMT8t
z3hixe1mLUWTcKKj38fQJm5P3J34kVQZBjDyHpwkdK/aDFTrCZDfNF926HEGHPdSxIjjUkp3cBNk
t7fsGrooF/5ZWIUJYNySDwq6hoLhmSUfBAjlXnNry9I9sr6FXkh/gBoMXBbd2YHc1dRM05o7U2MQ
NWB7SlT6WaxHDNEPBq8k3/5T4GL5+AhoCzjoJIAn6XTIchq3BpmMQ75AD9phxAm69h32e4pYSHYA
ZHXITj/kg+WR+nWVFUcuvf+D7UV2Ea7XZB/eXdENaLPWRov+dlfW0/VkSs0jPKBUAr5AjAFDcSZi
QqY5yC86pT+c0rPOSaYjmdngux8QlkOSbWmXOWKUnZZ7ZAK05YY/c1GNuBEH0lTA7ygRa19pin02
6h3fyo3HZzLj1dC6CaQEiA+68IqBHe3v0UBmjAQDYGLmsfqKUZQnEqXDfJPgU3DPpobvPW2lfTKb
dfk2/mxu7u454qGx/X8gLAGpSwy+s05dEvK/SFoGwrWG0dO8cTip+xkXIxuAovPCuYkdDHDVSYDq
d7YUfoPrvb8qGimXW+/XfB47nCHsHnl3kxrvipNT5pxerXb+HeVZmpGooodUA0k+1j3wlRLnaW9D
FjtX/gXiXgea0RUFlIAZiY+r+aF7+xk5dXMVOz3uXjtEmeD9nl4u/DTnvxoEAMVT1ARun8w4zmi+
Uop3/wMXrN768oPqJGNW/GOb8z9roP4DJezYsI00wQB75j6XMdXJT5cZEObiHRI08QmEG7A2PkDK
CHMX7qwWnwweICPCwfxtBaq7/amA0GebU8s/lOdYpWkQAx8Q/JWcYtVVAikcsta68JhVkkPg8qis
HyQuiSERDf7QNIkWiNa3rx8YsAXQH4ZDgHA9g6kOdLPAkYWbxmEpKNuW9cAe6p7Z+Qg6GI5W+7J8
x5y5vAYuNJ2CUW8vlno7De8wKbz5oiIALc5ivRAorRAkCzhZ1XADwFxo7edu7sZKXUV96Q12XMOI
rtAdJ4yaGVCsfKRrEyWRXvGTBROPJ4TaQ7swSbS8X4n5hmOG5DTqHDc2vyVotCBMlIRICxfJtOfZ
vplnJAYaliKIGCdapOhSxzxVHgN4Kn0dGYZGaen0WmxBVqTFCSQBYnfa6D6Ehcm4YGg0KcuCbWzP
ybRDZxFM7DsZseGWl+Hmq9m5sJlS5MiuIUZMOkntsIWvjEWYXrfBpIVzWHaweozKAHe2l1by31xd
4pr0dF0pnjNe9FUl7eIPQHznY1Qs7DqGZH5ogQKTp0BswNX52eZNj5E/SnqJnoZVVEjGrUfl8tnU
o/xswLNJVhmllC5H1CMVmdGq0S+bxW25QpWBLvcOm3WCu4cyHqLzPbdpI6NFRsZsuOC6XhIcZu7i
ee2HrmGwioLE1YQvrpxkGNiZ5Hqed3/LTtvJwlcZ4WGsdwy4zeaGIQMOLdMfJNvPTvNV/bufUdFO
c5Ya7M+JFYYWISubHhuyiuyOBdR51jCudsQ3i1EbYGgDrE+1zBq8dhI1nd9FQOoaSMyp5cLH1aPj
hK3xrTUnRuP7R9w9xhjALwaSO602SpQgNGPejPmAhSOhZSkPEMiRSwT4K9mLevl8WI0YKrFvAGpz
TFeA8QHp7Fy8qcqHn3Zw13uZiMJz8EhYo3lWt/8xGF40H76iEbvvn6f69kgtdy2mVJ06nsE2ra75
mKIHNieRuyijOXnhsFoSHjJMbzzRbHGUF0ILxgwx6TnjFJHiBeiR/6naJDTY/c3VfN/MGdKJUa+8
yZxJnV9LQcDh7IF4YpllvFDOZBWucrFcH2g4T13Noj72khizjNNdQCJYeYdaERs7CYRI2AnVarQ5
VvTsTwsWgFyOYnPPieqod5BZpTGaIlk4ctvi8NZ00dN85glj4J9PasX0w1UjG9Yq/OBy2zLTEjP0
D/19ukNegyQat9iWZx/R4Q4K6p/pCX3VVKdEz/+dCOO7yzZV2gHtVol785FPPF7QPB3Mm8gHbWJc
iHvb3hF7hAvUFaM+sjk/8lhhE18P3uSUfJMxoTg1jXKmb7qOXyFTu/Mpu/IQVUv3SS2tRdPyEz3i
k0e32UzW8r70kApYYpRTIDbC+hV62+NZnu1FRHsF/ykbbO7N4d21N95y2PMTGzBB0TludOYcfDFg
8ZccBTVahnlLLacI25JDqKeSNzckJqCMtWmxaaHZXCnkkUYzoGQVOG3cvF+WiaitM5fqYEJQunvH
YAHb8HYsVAMeOm2YL2FU12kyYiQ+/sUmdtWaXIl03fh6xwiIbutMQiJM/gkYlzD1n2yIoTtbK446
yYyy5m9mwejQvcBmhEMSjp5cTnSS9R3owzVqH/mZLlwJ6XvzN8zNeq9ENGSCr6S1jr6Caa81lWHK
Ft2WLpFAuvSjIPLes4ODVw5XPSURPQ4fGdbPJoS54IKz/D8yoUA0WMsztknCohcg94DjM1r5fWm2
+aiJ/o4ASfk0qLvuLi8oWBwruBb8YlbUmY2ACbBe95DelalCSXII2eHt6pLwQspo1WS4cIDCnMsa
ZiC16dcqFz+fDyGMdn1Bni4BzxUBU0dFbEiPEIWbf/Kmw8Dvw7Ha05dfFIns5HZNjKQF3dScRzwL
yEZL2M6aD1NY0LB+xKDnHPrte2TCUl5GT5iqaeeBDNgEobROKSAes72fULsFV4F0YRLwvYKEN/z8
JzNwLQ5+e01kPJZE3/e1Rte0rYCXwxPhIZpe/MEiSPWkRq5mj5KgfQH9zIEQOfkx6WoWSZZNopRB
DRBmj63xDAol34rkPVB75zdV1iE/rO49pp6tH09TfxYy1nX6f6tAvoCrnQpcHPQ9tGFgVqA7W++r
1Wffwhonq5vHK+5NmgySEZ68w3CAIA0bdNfQnHFLaamm/7S9ntv1ywe/q1INEqWJLATdMcLaw8EO
nsjmsWSEl51Jb4vwJY9EJli+fnHqQCh0LKmIfEVxyaLV9EghAAM8dn1I3VpU9UqtjIkEMRdWnhKx
Px8VocaelbdtS2xAdcOUj9ug0QaOEFtILhq5b+NuViwP/qHR+M+ga9Raaz1pUN6YGSiwf3/v91Uw
vsdONqsz0eHIcBgrNOFp7Rlq3QTW1icsVmr3d6l7YcFLEd1AA3U9UYEM9ObwV6W4Ay8wstsVcnxW
pzx6P/694tZJrUW5sK/kQ6smRg+t8UsHVfdqbLTkAALM7g0tRNK7A/9OpTWLVy9yAX7FgFrglMlh
naf+5VKXKc62dblX/rpq9icrHrBJdFLABbh7wXDJbvrRUt4IY5ofN59AbGtmX/vUEM/P1hbzskOT
uuS3/Sr/jivYfJelcfxnhuTZi0NcmK0O1tFAUSqO4V8tG7uz1E7SlCogSywpmf+Wq/QRMausCMMy
yHjqbns5BR8y325Nk9cxAflxC4j2SGH/3sdbV6Tzfh0CMsq9qIwDxG7haH0dAEG2lPrbhsZDwAmm
trk8gzGJ/aGjKKYiBdmGfKRlG3MoMVfA3UIai9MDbHawgDh4cbzdRDe7KPS8MNfGZwF5GxVDMRtc
YtDInp1pPJV0K0LkD/qk27jsN8gsYfvRrBVL3Ar31ng55Ek0fA4LeTUnhxzD3167+yAU5nQbyVBQ
MuDLPTKp36d3RWNu4vem4sqeEmJnttByE0HfQHNzEBdUfSEw53xqFTpFg670XgVvOaZWvK21txSM
iCjVdBotOddmyHv2Kdvbj8wKnPlbQozEA2RobZWE/PjZh+GTVlJPeXNDfThI6ho2+I6SeAUKuAOg
rYOyZIpWdHE/yESTNzpqTRhhFWPEog0JRWyarlfFiJ+NRFCIqGnGQtWSqn1z599fmT7SSC9TJz3v
K2N7TVu1Rk7/Z/sGdRqS1hgfnUCzXDphJEdzOrfgt3j6NRAJEntO/dRkisxKPQzM71SAtjhkfkb8
7CwZyg1WFNdbrzLBO8EGxbcJnzoqwdQ01qbMEvw6webOhhDuOQ8r+M96+B2FMuak+xLUwH+1ovFx
8XlZVeRcirm9Zg3uDt32nmAcdau+lJWlKb6t2VmLxIgnEfWVmJoS07jj0Ao4XHysrU/BZ02Qnh+g
BclG2L2wVecocvTTLJkC0/MP/YkA0hJUfrH9B90KCdhabb6zKrpJ5H1vfiP5M2eh0YJQ0AOWeAJP
rm+Mdp/0F0nVGh/R5PL2oIBSfJOkAcFfb5LExvETF2F3719umJiC8atITSYsh5get0BSTBDYqFZ4
3Ntulm8g0FbtfYSlxIflhxs072gRW0nrTaYQwRJPi+rfFXCcuQtEJJuSFT7wFy3PAdxxIFJSZn92
xNL3VuXOVVCoNUYB/+rhLy4HiEDkCYqrRui253E5zc2kjwXk7YQvnWeEo5jJ4+cUkW82kXpus0qc
ot96ndFwb9bpD3hVhWoGCvO43oNmwzEM46fVb1aab7VPD5soAqCWjwk6l6oux0NOdkHCGcUZULxW
ujAg5sbbpldzSYkXQCmI+MQyRPjOxyMT/qUZVgKt5Nzn5xvsrEIInKFD/GV0aHwCLP9SWWIjPhkC
j54dQP+g6iD4eigy0LONj088KHxeyS3MEnG31or8FG1K/kD/j1HybHev+A2JqJoWV3mKbkaqEcZI
+gSKG56AXrBEr9FKeJnHyYAia9BoLdw2sYmKlQzDWbxmSc7E0ZBqSdN7cOXCPxsM0bwHbG+3X82k
vpCDFAAehJop5iOdzoDBnmTM9nP+ShUfKbHsV8Z5meovLSlA8CwHtvHf1+TETjebV7yXcIwOwr+T
h/jm5eACIkzBq7m9Dc3uKLjkmyEH09xnxiI2gqfugdmGVvsOtXrjf6Mb2i/W8+YJcbh93yD2sOse
EStFjHPoVz8ie0woC0UbvPZcDMEn8tc3ff0pg2OBKT4LuV/2xwTnBpYUbmr8mx5ZW991Ijus7D8B
3PU1+oLqnq80mjAIr6rnXHUWp6kp5vzrYDI8OdDysukKKgmERDFulGDfM9XKu2zzSGZt+M6XESCK
rVQxhsCJlYCoHo4gthHT/1pHvwMf6LFbR5FpMm4/wIELbhjMD5rJ1Tqs7VuhSqr94vBTgJVnROf5
cGNlFhzhhpboCbi89Q4orO2EHk8L3FLotTXUWWX6bwA1A9otA9b0OKa3fUMaEksUB1tiRVrOOVtS
7VcyMfD5pmHwOmkqgBnBVsR6/mWo7X03Uqs+H1vZvqc1DBCChloCn0AU+l2oE0xqxOqInJ3gGHDO
hAtZrXjDdIeW1yQvR645YK0vtEDpWYk7wYmZULtdl0AmTj45dS5Wd/g0zuxEC6u3vja1rAD3u48R
dphYySzb4OXlEn3FpmjeehMxdfQML7IZ++a5CzjS5qFHBotTrxkaj3iXerflBw5KBi75HUispTwK
55B21p2lj0MvP4pMKV8LpTv8DnFNxx+j5UpjsI9s8qnxB/LHhDxrpBzpJdhg0MA3j3I8l86HtzDV
z0M8Gsk9hOD43nMoU86bkp/RSlUivP3BHgJG5W0xf773MoVX5ch/BIWPnziAfby3Y+Enybu5Cswa
K8rutbReQ5a4G+igK2rnWOarkV3FZ6hBwusqRjHC70mECEnepcosGAneToP7OM5jZqCp4kxn9HOw
kWP+DMzQvtLm1SfPLPsrO+eg29bHDaXvLz2EYCNQefrIxtEfDBWtNyBp4+uNah1UQ8udd89b54NL
+u1gzLBqX8IiZvRLFiAq93TZ97LsBpUU53GD0JAX4/5LQddju7JtqDsOTb5exxVfPQFt7xoJ2ivL
QEHJBl7qmZnEiepRcZvZYz63Ns+fpiMnJUKzvfZ/z/OlXD3Wpb/txciEx9Q4RPKcOrEstHYRsMGT
UnYsOnYUxFfixRS5ogjJpyQmfb+3hA7TLjwnaaJVgg1Zof95uKbzdbsTpfxwl90AanCvDBXl1EvE
vrb9OB3Bv78DCqWcgs8ABBtaggjs7STKNoRoAHlIPpJRa5TX9lkt/WtpXPJ+iX80qgCQ2bLI/np5
RtcU1wmWSdGiSkYFpgjnMA14tfXgNvMEKR1Vrf86uwm4bnwkznfjwkpVk58giRDPX5AkPrVrP58i
HnaxtZfguH5O8y3Fn1ZKU5aXiGpdplWoC5UNzPBeTQCKkGnKoOVJu0bf9pABCGy6OE1xBdok/TxU
AnTm1scxCYtAS5YM2nBf84aH1oUYDW8ldhV7bu/ITMHIyFEU4iI9UkY1E0TStdeQcM3mccfdCDE/
0C6PVrNgmKZxlJWJmgizndvIx5gNq+llrIBu70JgwwR7xWgZj6wxiVfqJpOe4mGarpWF5B/AkgN8
IwiSD8lwjCrhZ+hw4RiPlBC/xBSZ5UnDlUIFd004XSmDjQC49WknMzxbWfG1a83Q3f4xTLmjs1lh
ciA1Rd9dSRT9Xj7dUqyGCm2053rYUJqg/NsQnhZlDvN22qCScMHwA2DJdPcZ1ZY21FtWXw0ovXoM
z8+kKkQX7JCt6MJgGR0WSNfkKm4yzsKIQiCICRf6MM4TIAYV+dfw3LmjR+wRfiLbvX/TKKSYsV3n
6dF+9a+/QFzYxu5aBbYLfAOwkl8Ge1aq55KJgHtUkTpKl8jnTwoeVIIlIxuW7yjFQAqOKCLIOd9L
+Lq7pqv+pDwkk3R7nnRfzy0LxAQDpdmPDraJaYHzOyorZfx83fdfOza0doIlnMa6+6w/HzdbCcJ4
Udj5phfhFE8buPRW8fWuvzwI++aF5Q7Bf/eToLKmxwlWOtsDYH2/6xK1OCYgaCW53K3m6aM9yeYd
JqIrXvhyxEtnf9PekuAf7H8TZqlaFIcpV30uB66//UwYfpZ3lG6IjzeedRq2dUt/ZnAcpHbZdH/D
/IBVIUUoMyLAN+uqO5d6ljby8fpTvDyKNjlQrjjc2OVWc4xBHc4TAAbv0nZJzpeqX650gMvaZ4F4
ESITrg7TgCxPdnXMGrX/kjM6cxeTz5On2jmroLLXKIgvCvSiQE9rjbVGSyilvpTH+TQ5b3Pc6Hq4
jExsfHX5AeoHdAQQZaumoLP/eKsgGAtLgN9xw8ewE2bY1mIXKiuWrgPSEJnn1yd/S+PbVccISOQB
IsA4+8fkotTmiWkHNvYavo7lPj7tA5ONtiL0cSEupVOIKjE4C4VQyxbj8EH/YF+WJNaG4mIJeXzk
FImUTyEXndNgQIQxeg9smWRqAUq0+QGYtp7RFPmbizwk3OjY4zPti8xMlYHJY75Ux9V0W+hpiKwE
zuy8whX3l9sP0cLsw9BY4UGypTFFqKdLhmoLt0UT9YQLA5vrnXcwi2tSy8nJ8LSJz53OK7eU68gZ
8AR05GyESFGE7ASxXi4L6wc6dAgOhO8HiHmI9kw40ElXQpbEgMdklf6TNfqIXb7j7UL12119BjXg
sVbjZ26Gw+3nBZGDIlXiLnYbeLbgBGDHmGpdwfUIK64VbPW2WXj1qheYsXy5LKTJfRxmUwPnRqx3
YG//+jG09C0wLyxFtxa4mzx5byPJvKmmcb4NTlGlgj/3/yXPOiYDXDWq6muvyem6jZ+UZAag4Cyc
NAyHt/p2EmWwgsCzmjkOgOr3xSMRyUlcQTjvy7pIXbNl2oX15EXKjyKDy2UTm9sedxzBxAOTvzgj
lW+hCiYzNGNT9iqWSYeug3SWWcaExgTQBxQuXLcCKCS7fuXB4nqLtHut/qZ/06uWvrakJ+46uQ26
TYwP41u3IofMG7ILKdtjBwxx8OWCTbDy/cmkDPVVyzXv93zCQejHi5/85mH3PQC1PgiCCQdk/4iP
Tz0MqrU8AL3vVsALbs5UJpHpFBVhTtsTETV5RN6RlxOiHEV5E57AKTg8luSVkWp/sxYzlM9ZLxbR
P6JIEpSzlMeY8YczQOsa/DF+On8AYwCCQ0bnEQkkkSOHXfH3T/mJ5fk4NRTJlEhM950+IGa2kAho
8FOZ69tsNKfBxrCtkU/fp8cidTzCCZYTtVI4f4NdHiYl6nb4UoMNZU9yotCLXAvHqKy9YlYBtZu8
mXXjDrRYlH/i+8r0go01bp5BB2oX+gAtl0UUJtUP7y2nuUYPGmK0+28M31MpCfdUDXTXrWIAXcEw
SM8zkezKyf813U4SeFT4Sq8W1WIsA04ONCKvu7mCyWUZAgu7zNRoWMKF6fvongrSz6aifiwaFrzG
BGkQmYufTjgtrZm0Wm93Zriamw3Sskyhs6ZcR97vuapugUhq/zeB+Hu4VrKZ6YkBoki8gNI/4KDs
wcbiM8jNu+LsnllFKylwI662KgPpjPIaPoP2NCReSMHmBAzc2W90YWpu0MBxma0pPF9K1//D1jMN
Bpfmrqa2N7YrKFevdGaRgzAQ7MbtgYX6l3LzUax/aOZmoisZ8G+Ek5xg6rIdc/4z8cLOabashdzz
HFNjFMTGcE82QKVzqSC2RqcVCMS2FKO4kmM6BskQcTRCBlVlgvEyK07jioq77AdrPEa4LQHSs/Ml
7cgv9MpP3pzyXrJvLObyPm42lQsD49KYo4pudvui3taw26mphd2TF1LR7v2L562akLVDc1b4YnKB
3N9EUh/8lGrjHX5hfiKANv7iZWW6JpAXt8puQXqHV8YfAaud3CwxhOGEADhatDnn/LUD1sISMP7F
+DhkbrXYNpmQ22X3LQhxqopGY3qG6TlagwwsC9qKOlODWYYtWqyG8SmyDmnrQ1bNDmEEU/V2JJ3q
jCNnEwHPTJquHYl2EyrpXe6aXIYS1EGn71kQNsWS6ovLGGWdAsRd9+da4J4GJ93Fji67+Ta9SgkV
4maYQAk/pzwoy8f7nQ2KW+duIzpG62EhkBKQZzxWbliBk0ahGl51++Hcwy3QRbPZKmuiLKM7n55O
HeXpMMoyHqpRJ1XP7ZXKp8GIFUR1+W3Ac7gMg39sm6wum5MunvM8a/qcFfD15M8R4cyPyIZjKbqU
JYLDa2f+5KHtGBull1YemxOgnUieCymzmvPWDuT1G60TAh3zg9em9Cag6eF11NP9MnNZQIaJk4JA
TAAKD/1Z6f02longIkG4cWzDN7I1k/Q89+Qy4pofGxkEhEembgQQSSXD61gPhgestldpeL6uxvSd
Foje8uhXk0CBOFof/S4iwDFU/3Nz4hz7H7PYGEiAcTG0SYQKsM/StzR8qN9TH7sTok54Pn+j+Ax9
pLEW8yaFu3Pwb3l71futNfy0Hfq6lT1o1Ae6Y/IejUeiPNmxX2NIu0wj83uJfdNkShL4cLoYqd3R
RyR1WTkbI5Nwmh8YeImyxbxAwVgqpLF78rfbosSI3/Iuln7Jytw4Y3IwV9rK0zB8Y63OFuz1yGqV
AmCDYNfICfAhks7+rnflh592cBCGVIHiqLs6l/SK0SIrN8gyvAqgL2Rrr+gAEkTesMJ5z/catTBa
G1jMWJohHBXmmctcQNrtF+fE3PdgDUZiGBmp8ZS7Vj/SR77lFwm5o5JCN/C3LxIflC8iwXA3borx
D7riJ54KEA9GG/NCj+0x3OH7qDE3rUEcSc+nbFZvve3vul0QENJ4IRtcb7mMcSmKo/dUhZ6i+US1
seJqnghqmDK2u1cCQk/LfOyW+GDrtm4CyDuKBYtTelxJcG56gd+fUijFKwfNqeEehy6Yl6aoRCx6
eyh/Vn07wYZ01FmN6goRz9tIfX6UOQpoFoLyHEMJ2vqpX4DVWe3owJe7TrT1m/lSvoh9QqOeKOHd
bFm0pSFeFPAbnWwErZiGUIFJUJvPcyJnHjB86YucS6XPHqk8/Nb4AKvPsugY8NCZOEc7fiR4LcIl
UFfWCcOC2vGEaKCyCW+jKROpm7JWYwl7sQ0AUWjYGuyiwFTPWI6qgzFD5yEpOnCP0+8BduSdsFB7
LLVnLhrwlUFDOlp0IbgTc3JmDEj9vND9RsweLwCo88j7oJ/PoLzu8w7gGojkSxcsbqeCJKcrIPoP
CdMHOylRRTwvX17Y/AR53bGYHD8GEULO/DfdzPlSWG8+tRb3iaGNk9xUTlrvR0rBcj5KRH9/Cgf0
lDSmfs6qTtvGLQgxqSq8bVSyfYVWJvSmOydxyJVfljRSduuo4HjbFhPOpvbj5BYD+vR0yw/WD5sR
0w9GdOxAyMyHBttJsDMzSInpiHh4kgUmJmwClN5pm5/Vrt7V7q3BkvpPnJk50ws4TInbCYX/D54R
2LTTm/vuhgG4CjrjUAtJXpSkvYx0enCqAh48NZXv87Ytfv0NgAExyYKKJWb6zsai1EwA4OG5sTFl
oWReoem7eigBCQ+J2u0+oU5K9isPd3iVYmZQwLjILFwQgSAEZLXgsbZzcLAnt6ncB5qTmvUMcyqz
SOaiENNfgoTSInRh45+ndH5LOZFQHLZLTLkn+DClRd2DUF2R2Ll3JTlya4KOpbyUXPXWaBWoinV+
aTWLc0RG9I8Bjgy/LspPr+dolYA58CJDHng4/HLgJ4AkOo0up/AVR76qshZi2VRqDi3COSDGudpW
Hl3kncAepJjUFxe9Ix1a/Qd8GNf//YZoCyhkUe8Cmi1a21UA5/rs3QTYhAGl3KdPZcGRF28bYiqa
DGvD1r6w1lAreTBFHrAc+U/GpOryzt6p8IU5PdtK2oo5lZQ8ozaN0cv3IdIlpc2jeEdB7lq+RbYU
ExYeGQ5LoAxKpljMc/vPgn83mBfyXw08V7WBzvBUj/XFjyVrmOeyidESYj2L3QXJBGk61fMsKA3N
f34Zj0t8Dl3c+eCa63pVDtlcKbaVh96yTXrpAsVtyicEkoGZsI+jUZZUCGV9KlkhMakGJUeyZAoq
Y0z+D98PlLn4/3hBQ0z3s8uy42JII/ZitZwa6KMARzs/u6qmpy5pCRp/ogx1pRiNi/HNFD9iqFRA
mve19kcHvHu4hMNSM/wgyzxqgmt1ZkafhYhRyzeKgPA70J8LnK/xlaSLTDQRsFDorV4/S1G+TM0N
OupLPE+INzF+/8gc5Zx/YO4uZUTSNZ0G91Kohw/mzvy6OGLeh5T+KCnuFPLFQ6dJDsyMrl5pRhwi
qyCTbIp20qMfkigpgIiHciCFRMGwV2x221Cmwheo8Uz0j1tTj3Q2mRumJ+JjIxSrFtkUpejjOJJ3
3G1y8d8daXQz3rPtZrEJda4x4RMjyR71Scp0LfMaGsYscyCGM0RRE+ilrNw10t3vQB5RWZqiUDGB
Nj0GTKdvwkR0ygj9YYarPPDUSTvAnLsHb2d0bi53ZLt4PO+PkYrm7m8SjZHq/hhzgipMoXH/nOpH
fmx7/Kme95uV0jYOeVzXhYGr0TWx3MLNTPoiGFJunuzHOzVYcHB6B8IeU4HlpZWi8mQx/WlZlDeW
iCtg3J8isbwqLzp6YgHZ4jDIGKsZrgkSUWnP0c8lLRq7mlKV5mEO4lYuHeVg3gpcbDgMprPCgCtQ
nHXHnPb5JLPEX/2bq5plMBJigyFvJ3AnTaX2z9pTt9VRA71yI/yKo3NJR49eEXuVp1L5HQ31qHYU
y9btFk1EE+gtYkvg1BWmdriN0YCImAQbrbqvCffdLlK6MWHgGr8hVGFx/YBU7ovMS55K/INnCsxL
bxh+CY4kETAN5Fdw35h3SDdqdWklqM1O8/f7e8keoWB9WBHyGHVRdcwR7PykEPR2YgnADW29kUbE
KcHJo4acMG/fkcK3TgiwjhSJFolj3KBTmUOzaVsWMvNaQqBlK1TDbjnJAGlYo/ej+cHbAqoKSEbz
stshqvjmq4sB1P/Az4LEp8py1pmm7X+QBea0RmDoRrqH7oW7VYQRThrlHElpk3jYxi4MSFHivUO+
25esEFE2j9q3QbwCVDaaT3x+Xk02JVHQLHmptF3AmHf8l0Ori+M4MX53C7an+ruU+mXrpOaNXNc2
4Bv0GmwhiYDWYg/EqDuOIU43MdgAIx1mIhCQOCQ5JxgNryC6YBim8qhG0Tfzso9YimvtLNCLsuVW
r2qmzr5lDtGH17JyDNQzn8P0A7mHzN66DFCNnC6FG4kdcifTejbS8AeBUbSeNQr4x7pOdfm02fd+
f28tAAyDN0NmMmgmbon8IFXXIw86yXkiu4LGgAnuMNeVRUBTzXgUFmMncl5+/NrUF2mQGegUDFfi
CM/REgsZy2NCCjuF29IpDKXKTsIpikT5h8CVMcG8gFe87nJWvQ95SlnyG5sgd+9fHJWrOWyZu3EL
A4lC4XPchz1wOIVSgUVTOlTkeJ2I1L/dkH4MZA4gtSRzy3bWfIKemQCYgsTdiEKFNwOJmAXqF8RO
BPEHwBQWAv2C90Cj7Dk9orjNEylHm+7XZeS4hy1uyYwZAy6YnD9XHcExjPF5zBmf3Gs/sULHGoxA
jie3NC67RyGwuIjz6Xu+8wMsK1G5gz33U75L/HDAoRgXo5kLdQCV/v5sd9ZDhsFrB/VHbLlb2DIT
9djMiZXyKZLXN8mX74iJQGVXS8I6hkd0Szw6XEoJm759pjU8iv8VDtFSQgjSiI2f4guj+E2aiQjP
4e6mThXty8Lv4GOy5O3K+wXu3tlhvVi6vExvrFpzrLbQTAPl/p3ealDvXlx084XAwBEDaX8VpefQ
VQF6VwIIJ1NPKzkI6mbi8ElxkdI50Oy1B/VYBft7PG2vREx8nI/n82H0novTRcJnlXenEYjta9Si
0s4YwPiV6LTLElmA4S8ZfUDEf86O5SNLtHaRAbQq+hONhN4p5g3btUAxtG8vnlubGedXtKyQnDnT
4fd3sbke/r9KNKMqmTs/MGZMX9zdC4OHIzfY3uLH212SDdle0/m/no+UQVvpEsTVZYl43P5XWQTx
25SniO0xptmGhrODBNcxUGjEWpainhtULKMBLQ0a3QLdx/pS0k5xcdXhTxn2NAtNn0vCqumqUcW4
YfsI6OOj0XzWj0qt2ljirlKvu6lp7iPhHheZ7iloAfs4CKTL4bb4hI0PMmR1JMrFdtLrG7JHIIqs
6nbbUvfPWgBg4aX5XHJgfqP/PyWK++AsDp5DQhvHQ29uEo9L+82REh9bFxGbix3iG1ODp8UTrxVH
XIhp6VxpC3dahX0o8bctO1dKjl+7oBsb/JRgfvuSsmoKpe2Fref8OV2JKhsv0ag/oCwlMyU0CC29
cB6bJHfXdFuYoPwPDkRNLeN6CanBcvwot4hactVMaS2Z1texeREA5rPAjRqgmzNepwVgmwiow/h8
ysVU/AQQphxJlUqKOrHgnzVQJmNJ2wIdqzM/JhhpA5vp2XpOAEDqhTKQdWSsowYHap9KFpW3xMXs
WDzzF1g1HXpz5/X25QwZ67KxKR0EEZQ0hK3G/GqFqzxANKSJuDdH7gO1lhoDV2a4/sQj3XJIg1/+
tI3uEUbXFtVHd4rVXdF5935+pVei4DaXhtJWo6WpRRZRMZ0h7axfpyUAMPJupWDbTuoTi+VnZOtr
2xMUqz7/OrMsJXfZHO4ECz/kIJXXsjnwalN4G1/RVNSqzMwcUyIUp3p2DNXNuxNt+Hcj6uL/M8dq
CINaUrEC2hvuMse7pvnDrKqOsit7Dwlmp7hDRGsgx548T3mHJKAIfPMNSleTx5AZIDHTABD1vVwD
sy2hNvAAUF3c8JgIzwdhovNTQDMDh0M3bdjZsIJ7a5e0Q7JLkIcjThNsiVcRB3/hHqpEgS/Jhqfj
uSO95xHAq4zsI/RqDkA+2Y89A/RTDyspxiJ0WjGX4UMJXNCnDnghbf5GN6c0zWtS0cQN9G38Xfg2
wk2v2tZOgQYnR8qQ7dRBIiD2+CpvbIfgCCVJi2KiQKlsGh8hzBiR6EZiwGy0ipMPNXf+GuczWe6S
DANlNipZuMr7oeA1uDNFpVlMYf2oHPJgFtXv4lbZ9iBN7edUFe5wTptqEb4fyl5wh+qipAzBjWMm
mr194Z8K1/+MQV5+RggZ3aYtZueR2smmgaVr89693GpIUC5+AVabvhyL/XUKW701jY2hmC6Ua/qU
xV0yWuUYe+PueHT8AsKDyg6c2qhLZ8cljiXK9hKIXTxChF2kb0AGJ5SDe84SkhSDyQmKo8KBOIO+
dYqB5VTE9yNJYIoU4XRoWsf4FDmWO2hKTL8CK+vKVgSVJerFDGmqQvLDooWDbGHtbOb5hobqMcl2
lhAdAhdvnFqSgwTRsAi21Rw9XtWp+Y6s7SfhGppFX2z49UjRf9MdxgqjN6yoa8tNePpika9FmrnW
W5GBSyD+HN7S/yokdDeewRgz10IDDj3pqhtL49coimoB/4BIdvnrLSzQTAZuiD0zngRmrwoo3DSx
EHC2JyJwwKym9tGti2hT9OtgaCrVngJtj0kfF9qLPXJcysR5MeWgxi+6VYlZPvDlsCAsL4CT4a3/
2nwgkYdnw51nvjQr+kJ1YoZKyB294iktoZ3fBJWVfBEZkRay3Zlc8d9adXkQ/wrLliE8m2CqWghk
5nj3/Lo6hn7G+BqsVHqzyJSoyadEXIwSCSXOht3+HnsjNoyy65w2Qc5QQ2RdTVF+Qg+iYLFK1q7F
w0pkErCFWnT9TeIGiJBR7qC0ho2aPNWbzeB51zHA/jv+P0iYcghHs+j/dizMmFWWl8SZIIqoaxDW
mswwF1YL2AwCKkpPPkIpRutQcbmkhmNYxFWHiqjM0qnqiuoV2Ln9xS+K42+3fKqVWoFdcC9xV2bT
zHmODOvxOng2iuMC/WOoXSVDeF1qAGvB7Ya8co5J9/nl1Ob+JjxgqUxiVIdpWWYQTrrzZy890Arf
DzrwyC9SfRozPm/PLD10ia+1rmuj6u/iASV1T+K4R2W47/q1VbreJgfkOjodYJvLZyfQQ7bIW8BV
glzg34XOldC1fxHx/9V27j3BWG9o2y20IoEpNVSyuMbnOqxgR6bf9PQIcD1lJPHCChhqYzAm6XjL
VnnervHlByL67kvVO9NlfzquB23CEfNQ4FFjZV6vvNSffSgiwrw1/GmQ33PHtF9MxCG6eEPIp2pK
uJYE063Xo1+sJ1zHHfaJvQr0RX+fVTDhpn2bdkPtJu9QOvZV10+G7I8mGfsw+Vbs9CYX6aThN+u4
51sk5o0gUT3b5vLNxZI7pIPgMOSGEN0il6MaMxcRV/ZoaiylrVwdzllUsDfZU4PcFQ+/t7gVhsxd
VjpVPLZMbEho/iP2mdaM3qnFgGV2gbUtgzAdIFj58uHqqA/FKdbCGVypcNgmAdGZVk0zdjTOvZOT
O0mkMrHGCegiCFcebnUmzCgBPFExhJ5uwzdmqsYhj4yznsb2/bN5tDaVNVpWtCKe4SbCwsrg08xM
JiejluA9r14ZgGP6fqD7wnhOg1PX6EVtYLpBLY1odp28HLWIRNgac1Gc0hZp3O10Lqm73g30oG1u
kvxkBIjdLAKGElRy32XUdveFIQ/Hd+4wiI5VCij2N3y/WeZkEHRU4pAobhzi0cIoTMsFew9+abTC
rY9pxwN8bEXjS/qZKj5Z+BN/KrHflEkpZj0z5o06XW+FCBFrRFoNgxRU8zjqQ8GRcqLHuvJ4I5bo
AtjJxzXqgclZeY6cNBFDqmdWQP/ogy9CltTkRVArlmshxaYjRoZ3essAaQSn3fpI+5JmK3IbzF9A
hCcBNMlAljqBsBVCHH9itWmL++0A5Ysvs67tVDMhPis/6Csdd0V3ABPaizMPD7++FHwCDJozWpWL
PJAuC0rMj68Y2GE/uEmg3XTNzjaxEYk098W1o/dqQxvWpWxcWmWDQ1E3EBdx1tkAtKeKapw6CjKi
NWxFv6L3b88mA+qODA7LVyT6ZoqHub4OGVBzL/QHna8KNxlyYiax/UBtpzisMfjQ53BEoMPy/R4D
IAenFwceBRhTkDrkGUvekhXnwL82LMpJi0N5RbJyjdFGawgzFjgV/R/9Mff2Bpwdprlnl7AEijIT
hItQNgAwry5nrpIkoJL8uY98gCqu+eIEzEJ7yGRoOlKMb42YortjzqCYVLrGT/RJly9xHIWiusYq
QARGOi5ky+L/AoMLvppmY8eCfnJ9NT/oFvN7R4bsHfMq9qc959WijCtcxznMAZEUeTkEhtcFLvAN
UUD06gOOysHJlGKr3jDF/LZ+dNh7pcX29ajXwcHqIdJNSkNvndW7IvEXAVsiHpJM3jkGWuWtmLd3
UBCx59YRi3v1jiWrlgAT+6HX4bdbeGyPdBzUUKjP04ujvC7PXhPlJzia2X99kqAJ+zKpc58MmD2u
ej3zkao0mr2jgjnTZe+9V1n6QAm42WS4dQUIC7LGrY00V/RQfRR+4tFSPBoFo0IzIvuIty+8M8Cw
iPxllS17Dr4pcfkABJVBRkqZlr7Ft/mNI/y4ICgqDQtd/CfDJinACLhkiGqsOHJhXJhsh/A2S7nn
bBm6wOdZW++fZjCWNDbn9Xl+p8kvAfpnqjiInpogoWtfvMbfJUyeuQUx3HskFgIvdSxLtNC2DSqH
9uD7IDYxFXISaUYgMFflM43Y0qcJpzt4P7mWgzKT3LpANFemjHq9+vKM2WI2OY1eRJfLfrB+wmMv
dbDDejIZP4XvukLNhRBOflzaiG92k28fvVuqNBsHWQD9dkqPpnWjKqPReOcbL3qw3kmRBV+ydtFC
z58dmZEl3XPB2HbJjEBN1+Gp4jfOrKqksa+P49f223+yhONrUSbVG4EQpjI8pwu+vyKyuWBIDTLN
8V/YUFTm5D12jY4ZeAkH+iKjGqP7GiwZsDBZChzXNqU3mwD3TF6MWVOBbTiPU+m5mvv74VD8wVpw
VsrBxPIkHy8wxWhzHQwH4oxAOLqTaJychHALI0gcL/XKjZPuFjMinWw+mB8uzXUyOB8Xd9jMyda5
1gGEHVWV+XTm+SQsxX1wBbGfnC9cCPZrdLrital9PHqF3M7EoQU1qiqNLg9yPAvAYyPKX51fk8Ii
IUeUk5fCg6YbaUMUjQWLIocwpIzU7I4BoIRJAXuSeRjDhT2dYGZPtdspVZbvMNsDfn3U/nxtAmip
djpLBcNRZdjhfTzMkq2XaUNI0VMN8ajKn3Actk1dSs1LDqelK6KuPv9SvZszihjtMQkho8ZYUuef
lpKRz/RPz1W4eTaMsqWlbU56jS7Vqs8dgar+Y/3L4vwC5CKZk47lnaNFzvSwLbC2jSDV1YXboSiw
/01FoZv9z087xN2R5NV73xJB+F2FV1gsbpd0jPjWcTPglKB9Qaq62DBlPeBO8fqgUslsd70lTmKM
l5LGtNvOqx/JwWLBiOoG/Seh5pc+x41n0UeDEMNrylVW39zxVVKrse0sopv/w6lW7kolm39ougJu
RELCvIYc90lIoKDwnc713RGCc70zPnQR2Bo4RlomsesNJ8cEs8HFchFk7ZcNDawFEk5Vhz8v7pJ3
9NDhRZ9BDzkD2uuqA7GXADdSw2ZbEilNe5f6rnClsWvMQ3Tc6xeBXBfTw9O7tpmH5fDczTeJJ6HS
Nd8FAJjSx35UUqxxiGXCDqf2wwmKzxhYyLhj0Ea1OUHSAhrWFJ8KFhQHmcHGadmHONbojRJv4TsR
QVKQEuW7mWzfsRSpeyuS882zD/5Az3+DOrGQlBYWI3oMIbo7opeXcn7eQd28b8onAUOlnWGSwwKa
4o98SL9O/sV6GOdmO+BSQFcMn4ghHQAtbMb0xKkbWTWSjk1q3fiAgNmV0BHwrDSnraObzkO0y0yw
NEKNu98OX0tYxy80WjkOKwLXRJvxo+jvmICFKhgHTo7n5B1b3SFVc+ecGdA9KA1U+3wiTWDnx7Bw
raJlJueq+9B0oKZ4VPI0Eoms+Ug6lRmBicqFfQZJGjN6GqLk3xQLSKjDE7V0FjDHn7hVmrpiBjns
mbCAbuzH75BNIL+XT2RfcGZ9eqhwQyfoBblnb2tzbT6ntQJVc1nY7DRFpo6hLSl/jzPn8TkQqfHm
33IXJQJ1sLRk3NkuUQhjCXTGmomOP6NBPPcFQkvXTHHzhpIQnti95VOmyJX3PwGn59IlX7GhnXPc
kQKfrgtB/Cgurxcixf5aoWJY/DnW3SeDbcg12T3mzLin2PfA7AS8FsLCEHaPHKUKtMImKI1ZO4Dw
qvt1DVOfqRk5yXnEG2JaqRqF6ivLvwg7YuDxWhFbK8Tt8an7pDcDFgLTwIaEbQBB44ZAoqCUd4Or
wOczflbEAioLbXzmSX54bUw2OM4mCyPrYiApumNHGLOiWHewrXkd6netdhJEY7w0Y8wZTyH/DaqR
TcMzfK0ttouha0U3cnqHVVL5H1qaauOYgjohIH0ac6inxPZOk9w0Y5GIhlt1lsCWpWTZ9sw5AQjm
h5Q9QWFZt/z5aCkv3AaV2ozFWc2N0Zqi06xX3x/y9fcfzdKcg2fU8QWxZC8touHHaBMzbKzmfB0x
njKn3RfQ4UF7M6B/RDeHyGxRavHNPa+kd9FLREa3Nb/5+NUeo0yH8+2PDAz8cFL82+1hQakbPzMv
H9lj1zUH6VEJa8rLH2xFHrd2x5JmefMXElY+URMgjfhhlXy6yVIJdD7S5bITHEeKC0kj+/4Io041
SX/PCPbOGGwtas9IBle92JcYUmzpXSTrvV0w0PrMiUXu+Gx+liaqMiIqqwiUJcXKkK0yXuKcOSL0
wdGZntHBCEFMn8tsubOjuzH6m0kxavb3H3MMNx3esav8DjllTPL8e2mzuxmpQDsEvbRMQm5ZL6TE
LSZ5jK1CxEQXACAYV9dHnihihmr9TkV8lywC8R/4F2MvmT3T2t1XAeB/TPwhvsCb8OIJ6WaUD1he
3RF5mdth60PCdDwbsOyVDCf3FaQPpEZiMPA3MwN1bqUwWmgsUi3ySsOpPWblR15DVWweHFrzY+AJ
2E1/BUvS06VRyh5bvgB+BtcApz+xUcmjkr+2HqHEp/uDTyhXPT/z5eyiEA8mkoFZU85YmwGgUZIb
NgfDRrcQXgx5u0yZIlYVL2i0YCCYC5LN7tYc3x2NkJUQd/tFrMtB3MW1ZIEd6+VGCbeTHCrhZy24
dx+gkTaxo18cYebilhDAdUe9Gd3+wgUcNp3E8gbZclyDR/IPVSzEqQX2LOrfByTdoOgoeKsTQsCh
IGM9oKvhoOVeIObXfTaPu90F9cPh06wgJa4FJiabQlTRkotSN5BlnRz5MF0PtmMhhDAIzjMY7SC3
5jx8Z8YxG3OUvUN/aHERVcN80tKIgqThAtcFmHK2JAvzbLriKgza3jSiWrji8CN6kGr7e26Km8JW
cw3o0rUwhnkGs5PoubHyJTDzTsF1z44SnDG7KqjMjyud7glw+LU7FxzAbGXWBvcEkp6EBG6XaXVY
DvJv99z5jBG2h+ZO/dXmlUEpqyAG5ugIt2chxGFNSqkRIxT6udVA+ZPFXlj7x7uds25qFrM/2G+c
fvVnviDKQFyjuTLAzpNY1gwLYt6y2YTugwSFdWXLodR9s6w4i17l7I9YjBnHCkTluyALCXTuW4x7
RGbKKKpwNGzdq++ZPqaa77DoNPpvQccNqvZ26bpZOXEBvrJkk5h3BIvCMo3RsM2g8WflXBH30dXI
ttHAKJprZLInzReiWe1ewE3Zrv1TtVGrC+AL1zqmys3IpowLxAJfOjjgIXgap+Tfwx3ZVAD8WsE3
U+FsLoesQx3fQIbsWz48vIUuHuS+9hLjZZpUt32uOhOo7m7EtoMuCAI61a7Zrg1XycDtkLe3E8zP
/Iv7QjAIBtyNTi22cb80THE3k4REk1y3OP9HjwLYdLcXiwpDZfTDPLk/PJXsxTiVuCcjdW6wQJE5
JhNRtkPWLrDzm8HvFQLK1lrXFSRmA8l6S1XG72KAPWudGBeIrEogGPH9uQ+UE5l5vLz5qP7dTkpG
vQ+G4kd+oc/9ve3GVmONrJR+0s6StFaKJRChOYVZmY9HR1zh6vUbh8/FwQ2o89jc6E8F67ogUGK7
m62Qp/qnImlUrsRR9bD55AHbRfJuWtYtcJFcSEcMm5Sf3zU3l+hL9vQXUoIz+VvCTZEBu3kNudE0
V1J/202e0iuzBiPTJaEXu/ssx6a46iIMdcJqd7t7Guos3TWJH8M7eIXV02xF173IHXcyGYcRMOfU
BUmL9KqhBDR2F2u9VN3u22NmV6Xq6o+4KG7CVeLmIxNx9fIyYcQjNt0li5dRa2dSc6+zeGi6HNJq
VWxNtSy1zO41Dat8roccihJ3hJJIyl4dQ9Lr5sJSdLORcm3bbNnVE/au9nSfquIzQx5XMBzVP3N5
FrmlCgvPyi3/xVKVXb2w28nMskwRGGIodI9FGScDXNm8uQwao6sJVw+pvtPGJzsuPp+3Q54vRsMZ
AuAELx8DwLrk6fqpHcAzigfJ90eYgnGyennPB7FFiGKzQoOiyd2O4hYHhOwbZsMCrUuOmMaQkkc3
GkJ7i7ZTd7uAVq7FNHafVWOaqPCChSUvJqKAGyWARbhAOfY8hl4eHZ9Bka/Ezm6xIL91IfjCN8Av
U0YC34SCZUEPNbJ2JP/uVOyenGExy8JanoewRqaH/7zIH4T+3Du+gMWwVz10DJNh7dRSh8n1Dtpp
uFgqvXHxH6bVdnUrbbpldgzKohpLNE87woFCvlSHGqiwW+B5ukdAyp6GcEluYqUDqI3cgbBtoc6u
Zd0vpnvIFyOdzkbJPGnB26g4lbprXdhqNsYAUHldkBZ0QUri4kYo2au0+Dd/9S7dtxmzYyN3fdWr
RVyZKwzLulNEeCnj25l8RZLXw7USHydHDPChfbKPN0XZVnPFFhHNcRKVJugKWLWxdp4bMDEa5J1a
RQXzEl5PTeNwejkZe47tRljYcWEiXci7aqB5jq42P//LyhuSKa18Znhu8VJIHmcthmA5ypmnj6I+
HO3/LQ1xySRUJGmjyz7i3MaG6usBA2Zz/ljEUdZfdNme/H9n0gXC0U3ba0xPejTxdh5OsaEonaBF
vF1h4VD2wQ0scxz19SVSjr2XgJbXrlZdaNakp5HMr9ZK/B5AGHYkFgSCUx6+OiYjL6H60Q6G9KPc
4fsf1RmjHrP9iIdR6cxC3L6BL2crNfJz5P/vtYAG07HwkiJRuxeJ2+X0VdQDnWIGJu0m8lvAzLXq
HcQJ2DueTD41iXao74pcKDvUURXXX2YS0AJ3VVo9KNhQo5pzwIrDJi6xtfBz6a+mJs6Xfj5m89XO
OHqHR05d5CzPRn4cnHD5zQE21N8V03KMjE7vGxhKbVmKKIMLT7bOoMS14N1r5g5M3oDwPbYWu3ej
NIePrjxSkdCYWz3DwXONMG13O05jApGs3KsKiiZzhW2FfHClkYBUrhHH0EvkJec1lUGlNn0OfeEk
04uD1Hm+SZAeQvoQVMAsvMv2dq2RVqqgTGGTeaVVik7KnBCI7rNVGwKVamAWhrWi9rY4P55180Eg
ikIq4xikkAppxUxBk2eeq34flSocng8lMSBtdkBc47NU4fr7JlViZgInRd4Q600qz9nqqqQ/54V3
wDS4VHcDG9DtvUbms3xSk44HoOVG0vvhYmMOK9g9WSnGP5r0q8+u6WI5wutBAJTqTsU91WUBeTqQ
FDyhD7EatXyd5KWFJ6HXQMR20xIOR+0hC/RcPL8Y0HBJyt/a0a1WBwAHWzgzBebOkKlCQcBXph+8
rFIUTo3K/v0PKDsbnRYb2ajcfOzWHGYSVmBL+JB9+ilNOKvx6i5ii14mWTtugwYnOyS5BDA1rMbu
xm6NKYyBM793U1OB1GBDqyPeELpnNVwVNAtOa9ZLl5Jkkec2JTMTj0riMvfx0mESJG8xylKJDC/Z
4j9f1xjzaZECiNpKKW395paHx989R04gDQNEEQe1v3B6kLgcKvNh+iZOMkUYlsqApgh3Uyoi5Syr
rI97lzQULaGws4n65jFU/3dg3fmt3RNdslfhOI6eSce8uxcrfWZSwgzVBaKtG/3GYYJJKQei5vi5
vWQR1bO9xA6bm5k+NO8IB0jlRKwiAQNVTGeoAicwPK6wCv6qPz4AO8CZYOdpqRryoioFZIdwSCAv
1WG089ZMVuEf6e6+/y4r6G86IFDUzilM7auiy4xnivoUBENAoOmx/+F7A8GzSk93qzn5qs5ELPcf
0OzLQsv0tX6h6YgjynVVV9kX3G4HBj7qUWI4Vse3VokfBPVdXkTOYchTTWmGAmv3eMJf4RH0Ys1K
DccgVFXWNo0xMHA3LXCmcGFYrose7r8apuJcasV1ozz/swBC6YIqgV5eGxSEc6fuYwyho0IoRRxw
anu7AFNdD0NPo7AynB/66QDAQ9S7jYzOqwgeHr28XgZdxdBETBV6lDR7gVr84nUm7o1ge3VRKzUJ
hFkZptSF6lXuGmvJFzpEvYELHEOXjaA1QjvlISuqPGJCXueWuuvHHCJQZoXDosWDItpcoF8jyRQr
+UO9UytGMog9KerDJaxN4oMJgh5nEPxDNgDA6R6S98xt7ZUM6DpV0XLjClhQvUJ+WaAPczPNVZDd
sgxYlXyHpYIKdP66zqjgwOo0wCHLzbdtlUX2Yr/CxsmcrZIbWchRQISHzBMZ3ACtSKu9z7agTOQY
Ag9Yo/Tfwp/zK1tR9E0CtfsGMYIocEF3SvnV9KW+ymkP/3bCOgpcG7nTkbJ+/8e4Zy0Lfxnjo/Dc
sZqp3ERkdBnFLG4DWPoJYoDXqC9M0z5ZIOoSVuCjtEo//JMOBYhKaFCtGX/ccnmeW+SHXU3Lpggp
jVsLiiiwLTVBSA9PwdHiCrCfwQajZ3be4nq9masVaGbzkI74j41uCGeqLRTGov86NuofF3V9RzSk
qdmquNXkV1HnhDz2UIk1G1VxYqP9PDovCO4w5SycrvlQMtPxphiKe+crcSmKNNmxD1Jr2Qj068ma
S9SEGq8HAVE5Zm54pagGF391c81xQEfXWmeiVQExWgaKRt6m1epEANQP+RSrzP//Sg0rFz9VjOeF
u5tuWV5kWLy02cAX1AUYw7WqT7fHSTxdzgRzANbxcp2C8tVBuUjXvqgump3acZfvEiSIefsjxcTz
Ah1Xbf7cnAlAeZv+SA5OqY+PqUn7ePItbeFvJ46VaJADWab+dCUJsK5m3D51Onka0NdYn+jFoErH
9odPtqSbX7N8wB2aG6lTe6m7YcaoJe10TFHo94fiKGpIdpf22F9TeK2mkyaCfI2whmNLjkUWG4nS
IIpv1Tgw2J54iNekeSFgkJ1Gc9lsGciXFb9phN24uB3HX0Po3I/8uDRbyQYM8S32B1JjwRYQXgXp
M0hlUJ8tX9XQFhi2NKv80JSBvsLEt+3p3d16Q3yKOgQTgwovV8f2Co4Dh/aOw8TpG2mj4QaN6FeA
X6712WUF/9l2zSOiJU/bsnI/oTui1wifyLdtepTgAHbbywqFLUoj01EjuU1/hbh6ZV7PfMVjbQJk
oU4icWP/DR7tGRarrHyDHBlKSaavlCjYiBtZBjsVD95Sf9iM2aASF25Np8MRGHCTKNaWSu4USZ+G
4HttRTBmsnMGECWtcSyc85HxeMj82FwVHkkNme+WuIxQe/8DEwpnYSxnL2omcLtBV0JCIv9NxiBW
ZXaJRSLjbA8i51CeG3zXpjriu1OFgQ9aKJbQPHoImKpR5y6blqRwxAyHwQnEiKIR66FA0iJZOQti
8ua5q1Lcg7h4GdApnl3y8l/d2XXlEl2rJQKEWsHFGdFU5TH/CkC6Paqec6YP5q2dlfSjYLIkA4kz
Ski2HU4jV9ZPQeHMJiCZ26BTWYUD5M9u6+CIVifhM7InhVM3YFvtxLlp8u+BjBBFBF9ZoWQqwQx0
pMeoq5bp2RAhfqTOM8OPSvsx6H3cz4m+Qa0A3z/JaR8PGy00VyzrAhTDyRHprPD58zyljssnx8Jq
crxQ/F+C1l4R/Sby9Zc5SYznDdalieHRCCgNsx9xTgb6EShLscbm8O1FUqC18dvTJAdlF7S2tMBp
v/j05rt2ICW4qFU001bPXMhTmDNVkau4h1BRz+dRA1OdPpeT6LSCkQNyMBqI3gd4d5blntARTfpd
QBeRUcMV6FBnDUSG52d+QYnGZAxO4EdYWRMi2XI8DQBmv0VUphCh3s+Gt8yIdrUa/bbx5v0oaqQW
XGLYN4tZaAX/y6zG+17YO6oSfECX4YUE1mJQyruTGAoNcJ224qUkKb3BscyyZ2PPSRiiz1W9ltIi
3yFxfqruINads/cStxi9pb3HDR+zJG99rw3crvnQUjYFcUg9DKVVgoOJSczrob3QtpzL0w9nZLc4
JF7ZcGndTIqEWfhLfznWlfonMvHhZphMyeLsGY83T7r6HjfY+zZUGQ2lF1N2VSam6f3MynkCTms9
XTmISraBYd64P+ja00YCDQw2yQBPBvXSm5/kTZEruMfVMhkEki3dGczqAgCuHOeRxXMjUuHExIP1
ysP+vjAAVU9jIdWWS4YoHl/g0ABEQJs74jmoSNnMiMdIkluPECEHdI3aYCT1xkBl8K+Hbj/dm6si
LjTwYfq4GhBg+czV4txmOG8teolDxRB7pSZBXoc5gnILbhnJoAXf4cjn+EL7VzBfMR5QLDiS3ye5
Sj8z3TcteaxSU4ros/3dPe3mk2H3CV8jLYPpxYiW8gqaqlFm9wckSlaT3WP8VR2YPU9y2SOf5JCY
Di6hPCyRh6RB2/C2RKQkMbvpmi3sRNbNNxVdwRRrzOWxK44OwGi6Ks+bT7mxnbXHMujqqwOCtWPS
GolY3tmrfH8zCk001+hpWWCxElPOH5+x5ZnUmxhRTsF0uM6aXFhybmMnDN0HvwBTs6/TQLLgtguN
+xlymf+OULVUKhdAYopb4/DgiaLqXFUamqLYSt/Nm6a364yTEjRyCDDdwxsgyd3fGXteK1SnHAD1
fnUknQR9K3Ri9AZRXbljzOBwbscLdPE/5Z2b6llF45zmj3qco3cixGHfS6JtOdoszHRJPGhwMf0a
hkDgh+Rj2qTgVHTmGkikBaj91yQn6OFmjb1+71uFM2gj4pHRhI9b+iJ4q+Tx5qA4tgDPq3TVUgAu
B88IOj850Tdtq629P6N/CkBxgtE64970qm/f1eRBoZrERjSnwkTcCwVOAyjYZOU5Jtr/kXY3Eqwe
lDqcZvmZQfCbjMGi5wcoFU1BULd2SG3hYmOtQT5utPGziE1vzVk3P/6gR1iLQnHbzPF/fCYM00kF
xX3MjR4sTKw31BXDfKOjMicbUu/mrBRY80j03XEUqeB2fEIqtiiFkB/1jpO7bZJfpZG3MQhcgbqb
CsAI5GU/QbcxS2OgYZv55r1ZS4fVYM2SaG6SJtr7YhiISh7ElignBtJ4HL9fjfu3w/NbIuAbdTlr
xtZ2quJhQfHZmWuoeuPhF9+SmUObNTx1mdlL5rn0JWNNgToeGxANBAfhiy8hPfo8ypMBc2owyyjn
fMaLH/7IIaA07qbzmBlc4ahyUxefluvrJtxNovZAmCnGtvgjdQSZbogeA+4HHurVuwkWyrtUu8nD
ED4vFoOfFVVVZ+q1sJu0/Ij9A/KRwD9JgUQbwxHG7lgkT7FlUtVr1NxbgT4c7p+NPUmd+o91eo9R
/Bndpoyd72dGPbQmZ6d1IVp9Hybv7+g4Hh6eEaATNOEEVpswEhLxFnpiz9yfAcuVw+Pfm1FYx0zq
dC4/hCBPQ/6lmH6EfLm/R7OvWACfJnNnNrM0VlD9bOQEat/ubE2dAxIcbxr01oZH5ntauJ7kLkIe
AnyFmZ4R4H+ifgA/vkdmP8VKqzrb6c84sopb5ksKUL/4sgzqG2RWZxOqok5JVj+q5lvRNi3RI+Sj
PO8rLmmX5/hZ2g80AgunVMUE3gpLm2KZhO+0fyAcvuqb+6CMDq7IvhNSCB1mDsCMC0b7Dxap37pW
gafhffSuMnp5HrZHD/i94sJJjtXZmgUeoQIh4+ikiWla+BE4qQi3D+4EANgwJBXdjbUDsQEdvYBH
gE8oGlds4qEubEn3JhZ90RKn1zCN3zuNvkbPMzlR4xbKzWaTSQXRd15JI3bBHLo3u2/EK/JkRAKw
Ad+TRh6C5NjXxiV3ce0ictqBhgl+H09wpTn/VItgqnJ8b7J6mFsbZOIMeEr5IWOdjb1FCtc2O6k2
P/OcuS0CkF1tjfDPW5BFH9fdqKFqBDpLoF7q4IS/P1crYSMmcnOG8ytASJt+pppjynHyMPX0MNXe
BZG0zz3hwplLxrOT84tuMeuJQQQvblgJRh2x0dKBRIQMQMjNUJLOLTLoAO3X7B1Rce+qLO5RX3bn
8JUrlgM51WKRh+h+Ef1g472Pbr7T9x8hqX7GcCOOclruRnVr7t9xeOZZO8k8FS9R9dTogtlZ7U7/
Kw+woKj99FeW87iUm4OE+lxK1/dBfJD0QWDewSVJD2uxeVApOxxgqui18iJLuFHCuPskzx6DR+kV
/eIejzKY6xhsBk+Dtj0dAuTOTZibGJUa74beIztwmmgP6jOvbkxqS/oITgmCnY+tbYYXyN/YlZsZ
uNVi9NJYtHRvn7Wc8Yf1/0lYiBf/Ji/VvOPchBKXTlvcyq0y7CZBIEM3K2GOGi9q5ZOC53/uwNI5
vYnepLZHdsN/fJStJPFK8EDk+G/m3GP6ZR0DZyng5/kaULaQJJ5ifyJRSfFU4D+cOu9xPAYk5yHe
DIWfwKBrmOqq7MGaINKQhwiJzfsCCxFuCUdlrM7RyKoKYBJb++nO5XAA7uVv5RcprIFBwO04ZZvp
nIKExxX8A9CzOk76u9I8raco2m/BSwnpiJRTx31hl6jHD1nMUye+SvdWLpiI3fkc1AK2mBSEMjvx
NU7R/96P5yDJzP3AZRekD5/sGTc7GiQX5J9gK3oalNrW/ys43mch3efCUfjG3x6fvOQseA7gWozN
fkZ++eNqb4xrBAuMpiv05wTVgzG7GTDBVBUCnbqqwU4FuF3hsoizIXzMyV7KCImCfnxJs6VanLcc
TSty4kRHKDJAxKArKCNe6qW3ctHUvUtb0uU0kR/Q70URqRFPQc6e86kmFYuEbBw424+LOi60v7aD
z/yYjOpjUSjUEWIzjbw3kO7XG7Zcti1e8AIAkGs/iDg6As7CTtmZHeVN9deYL4GzuHZLB2HP6p/z
L8cBmPR1/wvhRdUOxcRKIpld6JvbnPtV0yG90buHsxxMpQa0sxryUpJfFYBhiPNR4H2cCi7NqRtB
0B5HoWLhxgT8D/Md+GUWb0+tBYDpAPImowPE1yeg34hBPMK9+q4uX2KRu2zNF0iPZtJLdSuohU50
NoCYIrZFlcAS3nxKum4HYpsf9FLAwZ0zZsLdYkpqUHnILev++ENsTNnKVjqLROCq65/XUF+zdWo6
GmmzYk74/ByAJZfvtUBIo8mTRbUh6GUG5Op27vv09cxC2Jml3ATab0XiYQzFyayQ4cQu/+AJ7BUx
0HhScYGF0zS26fR5U4oasUnbcJxONxMuBloGMTsmyZ95eloVpVtZx8en3dYAeeU1wgLZncwJo/e5
bMoRQSHnrr0slFCjMHbR3T07I8216Tfdic13NBRIwzQGjVyXjPPtJyvMf12s19ZYewfrvH7tESVq
mSvgHmOqFD32/HJVTSLjE/vFQ6lfMbuNVBXffVWPFRqxOVYcVDx4XshDEHZudrVRxL40mBqDq3Ng
rLIEj+bw05m/43qT9FEFPW4IXltzeG8Rm9m0bwSmZC2IURGqTNJZZbiW7mWs7HXZajaiPqqFH+Ae
7zbCIWfuK6HoU7i5Z4QVb3WqSV6guHT+gjkpR7gmepKhEdb6/bZdIrpoYQWD0Y2WgfO3Ni5DnjtM
KrXfEQP7U3b13B7HjO5xM0PmqT7tM4b4s96r8pAJUAvXwzzuXanjdGngp2lsw0TR3Sj/TygMbMAs
BZjEdHhH8AlQG7Kof/e+bxgnwMHix8cD+FCW5Rq/4eKdiXnYjcQfBtU2Qn7RvX32FzVqprmfjO1T
yXbgFQwMZBCb+I7tLRUSxfJBNx86UiZJb/BUpoYc02K+c9s2WcvXeE3lW5NFaZ7N4qdTe9JqCOpH
O6ZBb3YFD0rEBUHVABODG+DE9qB6b1iBnE2ew95RmMYy3Pq8Zhfm9JVDj8hsESAoWSuS4E9c3Xtf
Mqm0zSRz00VIKZWcub8OkgEQPiW2H8F5jsFbW5ewXJvZFwmeEMQJwkcMA9if8BsM0xIMPMJgH/rF
B1ohCzpk4ucFnha41OC+i9+bBan1LmABurTaa8D5db+znU7b/KQ4cPgCnMH4e/TSjoZ9sGqJPivT
us+L+Qd4fytnB7UOfqCStx3Nj7xJtfyR0UnHYP3yg6du++Fr7jGZt+wQfJwytuQM6kMkoVCB1Jze
ON05XDiALsMvsuqOYIBg8FLdPs23G067ta6sI4bl1uoihbzoAHI+GbA6SfUq86agg+68JXnLLKeg
RyNl8s/kTMnNHTkS997xQ9TY0h46ogCZZgEMZ8+1knKzfMb71L8evRAUpF0gvbzX8cVstCGz+p36
xc6nVJc4UPE21W4atPsfMaE6qBWpexKw5FFo9/wxqghom32L4iteQV9baVr53HRPLK6nnXbeWUzx
QbcPzgTdVB35HDgAmnfF6b+psxASQQ/A52G0vlFLU79Kii7jM5Bq6oIZU2+mWG50Xy2LC3poA1/q
ezR3TWzuVIZArW0Fcdi8TEkl26X/1DeKxAnVR8Qm7jKINUmjOhuS0hkjMufusS5SFTciK7cyCENO
Y/WTi2dhU0Ma6Qp1HSjZBRrsfQdxeKUhJj4ZUuVcvJlljZT4m+/CbmvOQMQo4ER7HlkDWBUOPUgT
g8Zwr5zu8/2wKmRId+xJMWbshQ6OZYQB8IZoRV1p3ODYOXTjix0QdK7YcgA2DPTAgFqH6qUsg9FL
Io6Id/qIABSwqypK3B9qWq/qD3VJ94SmI2+75MNHb+jQGZgXk6RBfFst58bcDpp6lvO9nf4OW9qr
XTtGh0TsYcTqRjm3gmWkvWSCHdT38Z16uGwlw/FKrwbvRc6109lAEMO/ZdEpnQaf79ckuAoX27Pm
5X9g5sV8N+CgkF7L52LZQTJJG/7grgIiLXfTcFJhKiU5Lvwb7liaoybXljjlZC7TLDKPzpimIuwY
p+h/jE+9cGBPGoXmxooXp9m4vVgxq4c1+MKLMtNUn6kmAf3hbFWfI6sf04Ih+/Shl1ocmos+KopO
PrXwD/Wj9w31PLa1NuwboJrfiLSrTQSPq5zzenFk+YVK/YzXBF0WX/vs6O+U5GZJoqsm62u/Jtu2
bIY2CrHShxVqfFIi4/fb0n6RNxYpEhYiOGus7V0LdBeIYBrOnGtMQLib5A/94X3BOhib6hhW3YA+
CPW97xnKUF53Qw/I0Syj8bEO7TlgDuRtofo8wNY38lZq7OaeSK7xwA5MWd8MDOV2qiB0+t7d770j
ak2+Z13GTVSD7Od+066Dedui2ktIe+zIBza7S48/UB4uOYv+YaZDsLTwvqrXWpzLh/+fHaei9bZ+
2DC5I6QdlpWbB98rfkQNuk/Glezmg0W8N4wkBoETXLZiVImMtX2ht2loNOr0Z+cNWrDsZW9Bj1FD
yxtPPfcuibRwQA3oqpdZdI4dIqHri5DAcob19pU6RBTIDo57/uGJXTNt0YztNpGkYn92Dod9OETN
bk/FYASoumpfoHo0JCXYed0n3HN/raoHzk1alKhturXkFFHsV9Xhn+Zv0VghHedKEKSUYmIVcb7x
UCDPLWj6qLvmGiIgzNSF6yzPqnIxivfFxjecVyqfH2W3CX2/OuQ/gtR3yQCR3nU/XbWkvCYIxrxh
F2TiDuPRF4FgUtedSURzoEGnkWCxMgzrMjXTvNnhF0oUEzP5COBtwPh7RXuDW1ZqFEsaGSP0UIUj
rqru5BXrCZwugXLXF0SeRHE2QkWt6pP57EBEW+XoJ3fREcicTwiG0V3dbX0Xg0B/4A3DFELxQAn+
M0ZcKYfUaWW3+lALCIyoqAUH22QIbYbGNHqrZuPttgg+HRpkl0GtK9edAg/00cGoRun/rf+2MjGv
MgDoe140I3Pr1koZqt/UXub4iW1K4M53sORqiHXlWaN9miv4iDOKq8wZDPVh+ojQ93qbzlvjjs3a
b3te/SPZZZRFMesLVljacTCIW804F8yU31Ip3gKZg/FM9NQieCjChTiEmftixYjMffdilnLX9FcA
Lm0P/ElzYQ5y1WVFKBW8eJiT/ri0kZ4w6U6ShQ5PQoL2nY5/32bnhlqrDbcVWH06ustlVIK9wz9F
RJ8YcrjY3z9sZrbew6clroHDChvecab8GibY7sOU+uW2TW3oL/w5ZTcF+iufSccvweLQhOg9lf7v
mdLkyyb5mHJOpI+b2lN7pzIki8eS5G498eeEAkYYmKRWPfedgDbUGnSnASLzZice1wmIZ/FbUGXt
aCb+85QjuGaKAY5Ljd1RsOAObStGpGSEw1kY/VRh0oW750BfHXM0ZkMBD24KJpeXaUCejExpSJUm
2YsLUWzpLw3EODweTtZSUZqGOgYETpGm5v85T5xguZZUSnugDilOa5Wlh0aZTsZ37fioV9/wyLMG
oULay6Z7Mjatuqloj6nlBmcKm+FGlQJFsqS6c2/wNZFfK8K3oO3B65rgCdu7sRXc0sWHndl0CA/6
CAjI7ktavl1XpGYGUW2Rgflr9KXWYNmsgCBMdymljewSDhWG4tDfLeY7U3wBV5PUqPXPLBvRduZk
E5EFoiuTdLyW+pSm77lPPg6gclGQ21rEB4qT0MeXT3Y96XuRguEYsVMcD+iH1PUGZK2Ma8iyNZK1
I5kjRuyRCrxfvhfdL9+Hojwj21FRc2/OZes7OcMFaepw1d9xfZSUr+07JJb9y2UOYFFX3xANw16h
2gk2ll+3CsROYPiSHrdPjvdgDlrnF0NfrOG95M3U2n/XTWUlNhtMYa8qlMevxbvoOiRdm5J/1qWz
nrtADo6V8XYNSasgWyHpb7LWVoP75iVsMG6+Cq8wWy+CzOiItl9UfwrSQFHQQIeG3DhAay/CaIkY
2oJSetx5XeNA8g93E9Vi+SgY6TCQ73gk00R+ShXlW0Cf43QYiQkeuFKMcjSoDCuAfuTvLHh3mdFZ
LgDnGNnq8wHdC1IsNo7yFD958+f1pfwCa0e9aLkllvfkkjxM6iZHiCRGG7GyGvY36AQjiSItdeCl
6a1X4iCzuKV9BkG4i/yfXvr9TfTJWdykuudCY3aDP5AHuoafmr+fHAtzSukSFTL/HpR0j1YDr4dM
rPWlnDdCyc1SPdBob2qqtk04ZnFgmubHmV8FHU2P5GfjaRN788RdrWOYmX1E+W856alrP90C1wBr
JPb0CslVoub1W7Gd9pTwmAgrJs32Bs+zd3Vun7KDAT/sBx15HodgxmiL2oEw+ctTrpQo0MVE+g6E
kE6Su243M7+DXtmdSTwuR9/HI0jkRhiMUSvS+dVW/AZesj95vlYrSRjWmZjGy3Q2mYn4KCu8lp3p
BiKwGawOTaKHE5usCA3F5BKX1+Z03AoyV/KwWWIrhhj/kRykQwNMOvaomvMdvseIETazwksAHHh5
Pwc3iTBQIlwDHp+Wslpo+A7wozykEvKPgHh84tAfZhTOrZBxdTx8dr2m9GKZ17udAU6N2SH7qGKP
RH3Av4/pnc+hbZudqph8PYpHMDseQcndwvsmopYAROsacXI2qn4Vr4MHzlkkZ7Hu09xqxGtVZogC
86ir2y+hAepBfF+JGJvg/6zRlrsVJX0WDJApy1nMRKzmgDoIU3vURDS8M6apPzsY9D4/NXzMDF/w
bp6xiTj6jOQgkCHnaadHsUfkXNF32c2y0ZtJc0MI4aINp5JPZEBG24noou7HndF/9r4URcCXThUi
3BGsip9v5lN6YOAK3/enuazHSCAmqVyvsOjnCsHtOMRTlksz1XVoOTOMgRFnnabrgC0UOoDEMrrd
dyE05wvV5zyC8CSg6htSXpA6Pbtexskd9xaT34pYO8xHI7wKFCClX48MohPnK/kW6rrIj8bmeZk8
G71TLygZMMEnHyr1bRoM9E0RBMlGGrqD3zVWALSrt8wBgyz1c36r0+r95uulzuQTaED0MujHT/o+
OomaorMIfRyhlttXNrSosI462dNpLEf6mWzFHnia+mcPVZqj4uxJyoyQDEfYwka7mPjUuI99EOzn
GH1X5b0WVU5nJyaTtEZUkqfbHQuvf7mI26yBkUJXxz3twayfg3ePoReakkKWuyc4oobKMPDRQeVL
S0DYJ/yEqYb6XTF/k12UxE/l+RGjFftjwcXpty7xbVud2SiUtVfgQXE0oUYjl4nzvdZTfv34csy2
MoltbvLD+s6yStDiN2zgAqoomUHyrw5ZyPaeiPgG1zce15n2r+81HvLBa6mSQAxKYDBG4qhFasw+
uMKKefxbe2LzCOf8Sa8yW6r7ogVkMhF4Yo0CdpM9Ptw1LPjcuhVBIXfum2WdDPOxIxSfpKm+gLsf
fNMvQ9ph/w2O1zBjzAxARYSjF4gR0JXBkuLWaxwoMRUKENdzCPBzVTs6kVVL2uqyfrj3MDArql3e
ZFAGgPdMkycCGuwJ0ESbD5NHdRtPD7Zv8xzmbvqhOxYAZw7cvIq5CnfKZNcuE2FDnVujYhfQwDCo
X9FFd04HaWoJkWsJAuRhkNGJcjntchDmu0ZF1j0vBafYxXoC4Gx4dt17wnIH1ueVuSLs8ay0ZVKL
VN/zY4CB3PV4RGwHbo3T9hmD43lVpX6wwUEYr1djEzx23au3azT3tB7gCRanr1/8hNrU05ArV5cT
n3LPrFP+8QRYi03gxZzT1qPNWakrbDmPYBB+l0+5U2ZoVx8WghoXq/RdE/MUej7sGsgeek8Kjg76
TELnJpJE8ITeG9rMnWpbmszhheT212xuV4mXE+zV9/yvLv7InQYk9PiSRDRxpMuVU9qRxXOvOFXh
F9meBuv0UbgpvfCmPFMEv+BJrYOnW06tgFXUgt+FWxBDkR8YaeaLwtb6oMEuNHpwaPHdhfROXbKt
SKjvPzjyaGLhbHSpusXPnWWBlQRjgCLUg9RVCWKDd3Xrll70FPz3PUbcr1doYzApSIIXG5VngbnX
UULxUuhkaWFxD0iByGWpLSRe3512RtcivzuaepH0qidIz39Hhzourh7KE51QfTBR0murMK20WrPB
GvKIEhLP7FyJ99/qpCEQ9QPc7P9Y/kUiHg2SIVRuHT50TpswlBLV6Lx7L4mXpOnvo2rTs/d4KjMx
NhyvFcJ41h9M49zk8/6c3w04MicH/M548XYGVKnTAL492BDLrhtAP004ttNs6GOfb0KOkyrSEVWO
/cY6x7/fGT76B9nbqTQZlfFAFjwSrv9IVPjElL9cdZBwjefgivnlEJhzSXgUgjWrTXma4aIrpQIT
JsrNoJIauzs+WVcmGKOEBNoJDIenWc0lEpWbUPGB4nekencQd4U20QKr5H+e4whY5CpzlyvOuxyj
fm32/Mg97aR0WjgZ6N79PKLobULxygGkPdsF/i4Ye8omuyqhXJS8Re5Wq728020+VjIZDbb5zBsi
+x+q3xr0bbRKtnlOowjHZ8LgX3xdd/CKfdyZMAsVZsGyAwC5kGX2kUrWi4iFHbE4WSui2VfB8wyJ
TMWOK08PgVUbMo7yLVE7ikGehM61jqR7/Yo4JMS4Uwq81TOM8pmaTp1vwzJ5V+s+CvqiZBUTfGhi
FUGGi5dJfZxz8Hd0wVBfq+qxNz0mfry4ouNiucoqc3yyUH10zcB0eM4q42mj93Ogw8ax8Ur+9Vv7
S+r1b9d3rXsSxZUdnTrgYsZe8ViRnEbtVGIhcCK5smUVG1ODgb9ev94InmJkEsByt4NHPbYt5buZ
0/wq1G4jZwyi+5yE3gkWuzvx36a5xmH3NuyUCQ+bXCKyGnurCuvx/+HosDTAIVhXsoxv520a6vVk
e69whXhU2avPjyLCShVKk8oiqaCCjmoBzMRHDAQ+upr/uIn7pB3CGfmEHKNTpTfNQnnquI7/dghs
3LQilP5aw9kTDwjtCKVeu4POquVwuX6jkQJ3j4sL4RUXFsr3UfqDwccPEMU+DaMqGpylV+6X+v46
EjkLK6PxspiY+rfDg+CGffdLwUPM6XEUJ5eYcR7hphaJffgissiX9KbO7pP4/b1K9MbZ1TfG3GuG
WYOrVEl04xcX5Yo6LiXfDh/g1cMV9sxNw/cAjne9li0m2hjNDuWSp5YzQGqGf5p/vhJDSwTzTc7C
8uALL9Fn2/wEUi7Cepjt+xaXCGy+c+PSgauNFXPXuzgTimip9xqLRlI2YZXMplWv3b3UKjLLB4zL
g0fzNuFpz4MBvYwpFw6TwVkczGUEWNjFJ/9/1wX9tzkTsHDffKrFFCTNvwNvTkgkejMdy6AKJi6m
M0Q8rW3NCdma+9CcVamsGJCiKbT7DnBSbg5GfbUeGmOp6ycsBv8z8TxVaCZIskASaNTX/INPlExE
tFST/6OfWZmpLyWHxgEQkx3AN3pAhGfzEN36iYAODFgw/8d4EaSk0RrpK6BERBGydhSYGLgQV2LK
t1RZKY4gfb79mzse9JOE52Lpnaw6rDYgrWwJurYbr0fqV1l6BSNpvS1Pb/4OIwjUsKkNMLMXEnjY
2kCZ/msGtNLLsGp2hCyplTnn3rP+9u0tNQQK8lOsp8bpZcRVIfr9Q7fVfdkjPDvoymZWIUmXFVRp
ifAkfEdyCjT4lu0YCQp1EaaUhjECV77/2zKKFGYT8vIz6/0jtY6ykQgHxgKrSKwn2jBDxQIxSrLU
+l9S2xjsYzegb86T1ZiYVxAXEjoyr5NPyRcyUtxedxH2WAm+omSB66ex1+cSkL0EhDPmWvqPX7oA
wJ0HxbDOTkX4gLmx3h8N9/Skd1ELhcDVc8eJUDF8c8Gtsfg+9vzS3fwPqdq9D5I6IVPHXBfTHaPM
pyPQb0jSFeEZfi63yXbZ9tj9IFbs6XDsR66lIvnocM3diXUyiGnSxEw3khQynvk3F/fWM+FibMnI
boCvDFYIoSDDO0v32BQglyxsMpviDG0d2PsstYqykSpMw4IdaAJoc760Lq18jw+577eylbmtjTBN
a7i9XrgPB7ifIoUWH+nfgORwSE+LQ62GBmBf26iycTK9nkE/C7nRSlbeJrAJt/MnWjYK+dkLEFv2
xxTj9zlIlcyNUv/WDin7mgNyEeR6bnMRhwgxcz/TwjofLQSMvRPpGu3s7wRsISw+ySfzZnLxpIGn
+k2OgWrmTmklNiSKqM4wXuRqcHfA2xgikcgn0Kl8sO7stJq0ekoFFiXi+vopBWJq/yZt0kqZFJEg
Ml66OJfaR9YpsuQu9gNyPSx771quurr+Ydz3rTeExBvj65BN4sXfCpnIDico5lFE0BDWYMsB2jlD
Z/LaQPoDKJh0251V+KNlMCVscaR6+8rAeL9TzuRFLBhPL1O68zpfdhdICKJQ4Ja1EYkRCEjlcVnr
+VBxFKUMP53QxEgjHba9Yp5MdNKHRAJXQrVCSEglfePMNm2Un3QdsiN8og+X7YSqF9WgebatlFee
CPR9CvzlBtmV1vkAcWKUfmoQKokSJmKKzE7WiCgHfs2pnWtJmt8ztH34wePZZ7CUBG/wRtVR5PmS
rfqf/5gbl34JRlXcqiG8mn6+c9JDTDIuevAre3uAaHAP0Uk8XWdJSZOyk/Uy6rgIalWQUukb6l95
j2lBpL0ODLMIJYESSVOROXqpHUxwKh896tcTAavx2KfF4rXunAsBMsO2TtzLAYNH1oknlHbEPLOW
shUUb5Ds4zJaQb9231HudSkJZ4wobuUmWUXr/FBZi6nlOjRa8VppqzJV3Kjhoefpz2ucCRX0Oy7k
TkNJda4Us/MHkKJlTdGEMkYRaRnJJefajCUb/cGCmVt4hK4+Xc+i0HQ65GflydoOTi6whH+2iclR
kfNMQT3YhjvedaPtU/tRN4AO6o/iMWFoCG2t6VrGtHgyJWXGCkzJN9uVmeUv6RXOrMcybjBTWtxX
6YqOvCWfQzSl9tWGHJ0d+1GElZafI14uswIFKnwWBhdIcg9p6ssSpF+wX4qAvVSicJvx7p8at8SG
eQwM9MLaYMyUzLyCFM5cKjhETTdK0JulhnttFHWREMtHSWajCSMsFXLBP916XqLjmSwMz9v0XPV8
x1s3oMKd7ugifbA1TMTZb74R0v8iwlmUVqigUC58d3FpXXyeddIfuhYhpeMFDnOsmlyC6m7JWp6z
LWsBUF0IZB2mOus8ZS6ltgV/bHo+nMrreD7xfyWeUx1mClmvfczNdaJEP2f3ilbPq+fB/EJIKjgk
yMqJyM/fv/oFztpgY7Mc6z7LZraZBwIlC7rd5oexniN+G+8Eggek+hhBDDaAnOaaXSzkFFmbVmPi
hld5hHtQjbnBolEhZ9VrGJJrAeOTRvl5TAgUraf3tJ/vXcdLTn0lA59/27bobPr+u2LjlCl3o7TL
HMAl4awiBbZ9WL92dOaJKuWM43+lbGJLcj+odfmKdxLmSqYCE+F7lA825/FkjA5AZ/0F69enjfNv
IwMXqODowOMR6PZKvXWKQr6SLkEOPYAZw3iODpjH3sM/zuhV4yNdRVIbVMIeNDBtj5RLXAPUDSDr
QFIizUlxAxQY2JikZyfMpeo9QPIKLCF1j/xgrxs4heHq+NCkrOIMR8o2yWM+TzqnLvEUGXSe+JLa
Zw6vH34Pn+T4adBv7QTHPh237DNzXuobYMaJNeSGtS+hANKs5+cbcegu69yZSJHnc5GCGkDuUHYb
egmO4WUl0NR1j7uDVLaofYaryZtVubOvAuhhYMXFsANw/g5IOXSUW63veGvFJ877mf9bHcApBHVd
UAhuNunPpueDuRmy/XpMm8GbKgCIIiKRXc0RLNTm6kk77/pr8l/Ju2cyZsCoJybi90nq4CLw8wgj
ZhNM8moIUrP8bvUdCinB7KXsoagw07P63UT7zB7hzsmnuztj6rZQIKq5+BIcoR1qX4+u9lCKVWTp
TIjuuPEdEIjIhHJLRvrHAoAxrLjCjzEsBSObCT09TuU8Fh9b6/+0hzrcBliWFIl/K7+gnhZB+PxA
ZUX6nky+pkZlH9r+2aC8DgplQ/+Qc7Xz2KZFtHYif6zqUYntjyzqnQFMMc6lwX5HLq2AhP5sANLS
B3wjyvzQuC721DthxyV+d69BsxC1nxP/5u/IERr0hl6qbJSOwMIh0S7G4fS9MguPkUxv9eNPcQAf
rJV32r6DorzMncYMqCUuX31jmf8NoksCuGYVM7V4eP0zr6ytD7wzi7WfFrxhIorRfMBB9EIN6ENP
ycehPfVY5Gj1mSN/1wokRfqdRdLhOcLRxhohA9DyzQYos6pU9FIqi2m+MnRUS9020tXJWGhdFRj+
z5fD1Uzag7kYjmzhbPX7amb6weH3q/Hzi2DWKsAWV6QN8MpIB/VaS1CDKORzuiVoAFX9E5ot4igC
eb/Zs8XsN96D64YptmYyyIRmhUeYszwzYPkYv8qfy0wkTq17RbLMBPQ0MvkKb7B6QVGBBjiIQ8jc
eabMqI15/87KuF2ZdNQfGm5a7vA9CoKUGUzcH7ombO+aWOEUYd++J3KlLyi/4xrfgioF2pMjiZwt
II4FyTgSmHHosPQcnBYc/pCMi11U3/nJGiOYIp+vawsubeW6CFCvxjRO24Ue62AsPPO64z7GAKes
JKrgk1ee2UgMn8zjcSYQ+q+qHrczaJaJA4TaOoAE9U5bwvBB4m0w9goMAb299sPmjZb2h1y1bv9p
yC+qA3PPZR6vXeiY9mPZmkJOuaLs/qJiThUKOnqfYhIxJxYX6axUuiEt6dim9x3dFLTSp8lDoqNG
sOULAN25D2yekcV00rbm/6weIVg6st7DIoLnySK8XmksEwixkfedM1KOeSJtbnxT49WoylqbGNx9
LLgd+ly/cQ9J/riolRRyM23hyxe2jXnxC8wicA5+Ls5PPtOstflpFli031Ifj0OWUD/6uqgEpinc
IpxENf4JQRvEftdBuzUwV5Kl3QMSpRd7/tNxt+C+zp1DldY3kAxW9VpU3V6KyyKzeWErXc1COW+q
IYjfzBBMfqJBayjD7gZ9xX3mnK7nFqRv/8IReZIsER+Oxiv/g+spsWOQV76cggkaBbVblUoVbeFo
AdInp9057UzORuOtTuPpMSk9U2rNAimaVoxaLtkK2ksf2FfsXU7qn7uFuWOwc9+j6M4SOeqk9obc
dMDHk2uVWzquFuJt1tQlZidtj4chDlaRPHynlaXqn8Jg9wlHwuKH7fMfy+E5Kc6MDSg5ql4YjjsS
rPGS/4/pWNeRkwH2bIhIShASvqij6GHhCjL6R8byRDt97vEpSvApN3388HczI3mjGrEBX+1TgFrq
FE3Z0+hqA/0n4YDEYQ/qaLzd8On3pPlXv7HBEuKC2N0JV/wxgw/nr/ZvEL3w8x4ZLMS5XxqgfYvY
qe6QkX7DRqr8Xg0KvDmJ0NP+feUzMtyNAgl44WNdYC//9FoSvNdPy1kGJ5JN4ex8+MMTANeMX4nU
alPjLsJ/AWTaeJlfjyjdEoZCu4XY46dW3JKe/GSmy2HzZ5lfxXx12IqihDX3zoqSqT1Ygtjj2rTb
IOXN13PYBvG5Xi41XGMcbNHSffhwcYtL4tvUEVKvglt5kZLdaT/sADmmMtpzi0puPV7sW5OXT5yN
Gmwo3ez5nDEsg7UFQ37CYnjA2i4zQwQ2e0FeWrY3qWaEaGvoOXU+uZQ45JoDe4CrfiVtcjpNeHIQ
B2vI60WcAagFY9hdWlX3hzXXUh5wpAFr23w6hf5jZ/IfReOd8pgtjharCcItIIEmk7RW3RsgFV95
I4zRUTVjlFhTx7ayt49BB8AYtu9qYIK6IvBKboNN3VVG/a/bY2gl7Mj5C1NF92v0n58TEbcVXQJg
mZufmslWHGCU7BY9zeZuC7m4hCtkuNlpnfeyWdvDb0GrYvO2c/a74KKF2B/LjHoTYT23N+ZtySZ9
VUidnvieGpN7S35BLrUnBJIE7YyRqBnKTx9j5eIDCEQI+Js56ydAZlFOAwx/bRRho0mMfoVU3S+j
+nEmZcruYTVZNklfLLdORIudpzBQL2Zxi6BRK7oYSqt4tTDX6tHomMS6h6ouM9mUGhzMN7kwMGf3
Gy+8qiTnR50/CTeDndJCW6oW3rRxj9Fp7PSq38AEoS2AaMLHqEvuEiTIFn0EtwBU5fChwkcpCUWs
iWfolvLnG5bMMJDBiUaPjxyexDB2jBhhCcd87BJASK0kFe5FG6gfdMMOHEOhkoLCkItcdeKuHbNk
4gtimFkYU0KBD6dYQfCuqeU95jVv8iqeyxWrGfucjG5bvAeCpeSVRGdJA6WwhsHjrPIbVaxKe7/G
Od1AcFzWWx/ofBzfod43NYwu89JihiNboSKEuQjGucgg0FhgNgoeHljm9vqB/GSMCQ0rSkfSd8cf
Nt2tOSVK1JdVVUHOupDs4R5xHgqNudjw7f+GwqakuZmXOpD2co0INmxZjyYQFJALUJJi/ytrueh3
rcZca9gc+ArhHbTDsD+SYjQDQfmzyjYJsb1ZVJpurKzGZRVactmzwitL/wdGtiRAk0IWfj1HM6h5
0K62o6gFANZu3P3WKwqGSbkjAtuIBZuXa90MHTylcFdlB+vfqqSy3rKImjm1tNYn6yGLF/YqIabj
knsctJDdauE/++DOblJt8pf35f+skJ98lZx/bcrJGdHBlDfFmannPSqQpccJp0td4GBb20uPMweG
7twW94yAMrWpSsfuArrJxQX3KQgiudiVwJrlwJCzIlUqLKRoIGhNdSrHr0TBxoQtw4J3uUuVc/o4
b1geExjehSFzFcHqDbwyqRAnub57x+SwoEZ7XU1H+2hYUmgFr34fkfthT7kZ8xEayTplPnqBwecU
RoABRnKekdeIwULJ5z9R1JDAUO+CUG2McugvanJTANtt0XSY80WQK3m7tHwL3pm4xiFg3GXxLY0b
p/Hm7ihY3t8W/4ZjftEVJ4DZy8SJqjN1LDYTNFYPaubyyJZ39kk+abKuXJBO2Txbdk7QLHslsLn9
FfH2R81Pk7dSj7q2k22s7CulDMDnyCgEpt/GXSSdPt7US10Pz+swgh71xcu6FbUjFpVGRAWWgbti
JyVzE/DsaysyREGlUk63F3oWNosTH5a8nnp6LAQE/S5aU9HU8LucphcX10h6bPEvYsxAkXB+BOyu
8K+ZopBsMKHRnvTPF2i3Xjb4b2t2+Qx/DS3EVrQ6SRjSQx6qVUug5rxx8XwjMlHQHgbFQkJQKmpf
hMVI4jZu2yzFA6WOPe+EJfOu86gaTTlvsSi00Y6cHUp6Wh2muiMLtf37QxKjLsk1BzkZH3hamm1C
hMZO8CpCKcpmG+yfuQjiW02wq1e0F8UjxcLBhVPBXh85Sj3lgmHtCCurVixQ4i6Xcv7DBV4ZPD9/
If3QOKTJu7OJNneEO7YcCWxDADf62cH+7vfSuvnGA3faUX1D7pK04aT6IFE/JoEZ5oUDwhUlmgwJ
0I5qdwzVB0dtIRyqx3UHhe/jl6MtcmMX25/nArXq2Tuojvqxb3HQW2pmXwGyHrL1RqLs7ilHeU++
lj6tU+yzdmnle+vSZROaem/heLXmFCy9nMd3meHmb1X6J0wLGMpWOAZ4uCbKFuGj5SKDUKQkcRte
IEQ+N9E1qlTwOohirUZuw7ET8qtE/hKmEUx3/cpstS0cKFRFmLA6ueOS4Tg/tqj1P+Nt/AfAsJS0
ZdRh1S0sWE3jMCQKYfRnZct7w52Wm97n+nsaCan505ndPTYHK6jPMSLGp8cEtXQ17xk5qdwa1F4I
s0kLwxI7jsZvfRCKfAmQjPifDcvS9EoRB//ONEqoWTngSm0FDjZegnomvSNmNZyCLcDuNKlizmEF
aZ2q+21Yg/OG8mAo+iyj4HOtfkHBH1dpwTlJHWM9gub9GXHqD/299xfg1fxamEl6W4DSKG023bDo
p46MN2QnZTc1gStApRGRQju6YDtkC4YDBxovJhj0mE2N3VlnQB3jxWhPOhPXCMcoICPpTLU/qCSS
4lf3IRHBglf1pzLxABtgZvtocf2w7uhwDC8oJF9VJUpXhHDhiudsrVi1Gw2zx05Qv8/QWqePbCeG
8kISg8avheoz9RT8b+4Qr4wWGN/7ZPBr3J1PF5heXTmMcbr/aklAalt8NqRMcPNqcLApeQ40nB/s
h9DuRg9tnVjcRQn+q560OhVgmVYVmDkGypIlQWF9cSQHI5GT16hjo6x8lV3PdxEYbAdH4UzUOmY4
JRhJ6n0fxFINQ+L0AD/gJyigaqELW5scD5D6iu8LwUVuL58THWQj0lFVOIolmf7ZDg73KmRJ6KDI
mvkoeF4oyYXsBCGqiUAdXJiWpHbIi2VgeloXPXDU4jmG/fZIDjw4/RJVf82A5cm++s5CWfzjz29j
nXonaZ/cYONKj0xxHKZ4zIXy4ynxnRREa3RTGvIZrNimrQ7UGPeRp5A6mnhQT2sKaxvX7rvuN7vv
j7XDKEhH48efL9E0LFv5eNY9E5D1lc/FnAaGkNL0iyEqFLHj2K8X9gPFhLJ9C38KoShiA54XXzAZ
YCFGRz6QvBOFV6wXB6LvcNvtndhBzRsLVSJYpm4KqM+VQzmDUrBmebNJwdBd5Mvd5PfMCCcmsaCW
73WZTQ5m49gpJCejf1HvO20f1I+wEgAHuAAuA60oBFHMX8t5aHt69IWXUIGbzweSu6BA71XzUpoz
3cHYuQjbv1EDsqgqy+NAR7yclf0zMaCTtHb44JBBIw06Y4XolLWiSlou9WT6ejzjx+WiF48T8u4T
6Y6wBUz2bDVI1s3yxguDLNj5lPYHCYI3yYevVCwRqfB5vXjsqKekkYQAfUVABJCqHRL+UJkavHfc
NmJqIRXRn2sR1PmRKjD+Q43GnzL2Kp1g2ZIUGcBKVE2r7RQbprNGgHBvKMyMaf89UKGUjcscuJJ7
9yA8H7Atve7viA4pgkMjnMNvLiXqNvNNm/wxNJToGSiVb+f3VnDJxuJpgmfOZtFJodB4mMw4Ylwl
aTe2OR+QOXxXOQwN7rrgo3CU0lNq/Nbh3WdYUaj9yGgjsdaJV0qYD8XnG9sjP/ZtUu7dYF58wg+I
r5SGXM6HG8UPD9Jc3aaum5UXaq8Aq34QzK0/oZu+baBlr9RY343+zLGSrBUWs5dOPwCwpQrVlbVg
YLLQHhhRPrGUFx5YTS487eUA/2D8+6jqRcF9wXiDgXiayC84T3xStAlKqPnwVaaOaaNqyuegnt05
VFoMsbZYp4yB/huWBH9xKupgPPE14sO6hXxBRrXupJbVOqqEq6pODvJ74TRTymfuUv509wxJWx4e
EaKMQs9+j/Hnx2EMkZfxxjzTHpZHL4CFMnHIaa1S2SC9Hfec3CH4ANfnOgOjJ7A/TUAiaTruckYK
tV85FKBj+8JJy4IYtTzTZ5/umgwWjxsf20aApPVGQ1ishe12j1Ifq1r6UkAGUrXQNTFC1WgIyHmG
ehWx0MNMain5qbpEuNApdMb3VIR3usP0QcZoaQ374DYGYu00I1LpxTosqS/zMThlEN0lt5BnnwNp
eE4CwuRMtZB0V4lHR6LbTGmOYJ7MVs2GDaKEXvS4Fvi5h7nOre9mDJ2mF3RB55k4bmgj/xLB+oDz
pyABnCO07IR3iSN9BAnSsNZrqltyoVjcteusrc8AIWDKHseDyTdabmHmjl/ZBObFE91gWqIHDLAx
oofbzo7QLyOGpm+jxjezUkTkCn+kErpcZcz9LC8h7aaW6DBCeCXVJWULb4NHpC33eX7Gx0lph/im
rSUUlPNMaADcAKFCcjCZxz7lv07nm/HVDYzg7QWjbz4aVGNrPjk7yDZVYzKJ6m8SbrYOCbTGN/Hh
OyQUDvUXj9xN4p7gM0dld7RfYG/0kTO9uvjLf9sI5Z5hoP3u/J6Yhw+MwZxuVpcN4j1NHdBNdofe
rjVSPMzMRPEEPZ1pZOFyL/N870XpMfooO0jiGzNrJteb4/7SqdgZDRZOFdi/FxCjaeakpQenolUO
DiLp2Whe4FQN9va8p81nibPSEkW/CE68gEVmTHawj6SGuG8m+aLdjhejWlehN+XoP0+1bk/BW5W8
Djnxecvy+4dI2Cf8CJu6yaiUe9OVKP4ov/tLPMp4DOgrhEWIBhW7EZGoGuzwngg5uQnEEanfGFM9
07hVcDKfBPXG/Itivc+oEW0hu7BMK2giqGL5gZcKipcBPND95hWmHcxRqRC0eOglYZaPbYoe9VYs
a9gjOxkQn6lPWdoe88Rbnc7I1KN1vvj7KVyyHMMVZyvtQr6uYL/FkRucOqvsihY05ocDcGGbNCHZ
UV1HGTRfH7etp9OninEM8JSw5SGtxUruHeS91TVf6dBXQU5OS5aY6rhqtgOVoZHXhBm7uu77VDCe
Xyabpo+V0QiV2rPcYuSCTfWNjIxsN+bemAWPLZjL2e2qLQZuYQjhOTqnGWxfwxkPDgExE2vdHdks
OOmebFL4SbsBPVXpe/whpm14jEO0Yisga6i5hZrsVxPN6z2/ZLIEyvM7l4GsJ4OWtGOdLZccMQ1s
y4NsOHnbj78FyW4M8hTMCbnp/byG+vQRx+PWcagxX2sDVV1xKpd3cwF47ZNvqrF3oGOJ9UahhiGq
5hnicSIDRzD6RI+IADLCJ3x7J0laxSE8KWO7reD90/r8yLbXJU87fkT7zJtFl3KrUC2RUT9L/jxY
nSJzsn8Z3vrSdP6PQXF1hOeOMjWSLz91eN1Hd7sPesLO1Rjy+DGotziyZptYQJXfMaht1on3VWvq
IZB4kXujojzbzRIOTQRi58j8FJrsiKRc50w74nXjNxT5WlKpzmAALyheUhMhQN+/7AaQ4PF5uuWZ
5ohl1FlKH8NuRGCvNd2CzXcUgiWl9J40CiUbvBM30O7ZITxs2myXhp6tdT1hZ7dKv1GXM8bAC/FV
PKtDFIlU7G2+Qynci7CX7IX9T9jC2AM2zIwe2vOPn9Hj60Vw/6GR90FbcoauAtUHKXMQV/TsNTW6
TUKILfVBb+9SHb3Fkv1QDNbSNwapznAbUiguCvXEuj+2kys9Cq5H6M/OPme0+luuORDfF03yTmwG
vCcZ/dLChzQi6DY1+PFGmXHpwTrG5knmVGk7FPW2H9+fPpV0SvmH+t9V5MaQngbWyZQQ0i+6y1mC
YXAAqgUBYelzWw8qHvoFECRI692UATn3p2j83/hmQUZ8d/mfZFZqXbq1MmkUNtxXG5WdbR3Hd9DJ
uPTy4OQ47LgXwp8F5gP5zgPo7vLE7pk/ijjq6j2+XQqJPqVciIM8aGDngmfhXNNbwPqDUxIrX2Pm
rI4BA5bU1xoIQ6usk99DoXqD6imZuImgo15TsphVBW/AOGNQsGV+sqoWWMqmrI9+o+SVSa+oLC7s
bn+353nAM0nY0m/zli+XGbIpm8QFMd9dr0h6spRKh6PFwMEgTfKl/ScrPRG6Edc1WDJX73NHiSCW
1RTcnvdKFXV3RJr7Gi/njUK032Lk2Plum96qmISlJ5k17POzAPPu9YgI6Edt6VBrRb9EINbZFt38
CyyCD8k1xVCLcH4rCvi32KhEu1CiICnj6pcYHx3nU6ON6PMyWnNSG98X1Z5X0hVcoThHarWTAIFp
zf3tzJYbXKNoSE0kRXtzi00xFZUdegRhnQe2ziXN14VCtZ3lpn0yIVlH4hNCo4SWjviK21P61ZoV
cI6t+dvdDAHw8YFKkkuiPjixzX0zj5m4d3Qrzz9ZwEIGnuMWSmNKz37A2dqO12LnPF8RC+Jx7WNP
1WDGygcJVqefOsk72PmZUbbtAZejZUznmPVP+EqiGiDAc64oKx5e0v/HC3gYDcQcRw2Ivg9LEgzx
6H3R1hXm3EY/oq5jPjtXg1yydMPVNCQhUg5yyTj2V34YrLH7E0hGTArZNqiubpRiTOGxJkB7OmSD
AFzpBGe8aO92CFsdhwhWANEO8Qi5kAqJCylvNkB1EYdO4X3RrUUyMOUT+MBg9bYFm+s1jEQrPKk6
DrxQ8oCl1wrJ+p3ZIfnCZbLj5A2WaQSJbdwA/9TKqtaRsPI3iOeH7CYyixFB1ds62rtPyFRY5rEQ
JBzhutiHPOWBsjwqSdQWD87cj5WO07Ju/nfzD2i3pa9CfVQKmmhlSY6qmaUuhDZ40kpj1nu6YmzJ
k7AlNN+vhW22REmLiGO8ICF8trjd3EnAjHUv0SM0crTSVvajMBXwOMFraqjSJQbbjhjcIsfrOlLI
5iiF3jpOfxFyoUpyhLj0Ym3Uhqq2furgkdqvU3Q6Zi6yndBilp9CKx5oBVZW0VRfaPOLD3nP2Qhi
sZnRoAqHXF6UwybSJ4MtZZauZxEs9GriJNSIvuKuz+T+6DFKdr2Qgjp/cYNqZDAdbrOVScng+DW9
kZgjsLn0/5wSgAQ8O99sGrvO/8LEjbTEqrYjQ3AQYzoDdWs3P60YcGVv+ewQeuWmow/+xedVwaJh
UXjfwZMqEh2NWA/7r6wjiWZP/+Ie22dJf+SJjXzmFCAinCuC0qu8INIiaOlIbVW++pIC/7wOHgJh
BQ73a6wLxTSKSjmGFxxye0u0xUYlVsBx70kVwdOZPXYup6QcSgTqxBNQIS6eSDUXt027WjZp2ZeR
sMxQny5sRoC2FptHpGbxzVaZshgqLeeXyzwBtEIzTr+iRaicSLCgfeKgVb8zSbpJ8YjucSvDpR1p
s8+u9ywt3jjGFJH/jOdfomcJoMR7QWzYmWPd+ICZNDp9VjR2t9jphAIxwPaf4nqJzEKEYqHRyPhc
lAwiW2UwWA1jdLnE+Ox6izYusEF21B/iwRenVlV4a/tZMPWB4D5tMN16eAQ48CEzThkBuEatQ4bz
ocwzNHvGtwIaDVgYx0X2o8n/218cQNHo4pScTOHUT/FDO4s1GMqe9otX4W46XksBNz2DKRH63i/x
uk7ixN+fCelmn83r8S4OJDEMefYDLoks49AF60DtZRtHaMLaoA8wVdGKP9XqpT8OE6MRv0hHPU9N
VMwtCqlC6p+IqMtRsiYVvl/QDweI+0BcSffg8EFVe5CN7zp9Ib9fSidzc/DWOdUqoJ78DzLPs5pI
l167ljrlmgRXYwWaPtmXtThND3SmdXYwpGn3hm7KkXOWu4//MLSXDtr8z5fTfvTASSxYB2fs4v5U
Ws7Y0omPnjmU+/QfL14nym7gTTvJABhbzNGM9Ti8mrzMwBcTCf7loiqSYrZObfPv67jFqCA8tm66
1WaEb03Gxu9x4ZezlF2J3rXJgQzS9iA8ncdu/uZNQAuEPVuhhdotc3jZCnG429tFZlOFzB1/6hms
KYG/0V+yaK69fiugaep22ZGh8kJDBdJO62dy6DTFRZm8rwfVXIrCdFjGYUxwjWkwPRRuGbttNm07
A2yGl99Nx65MNfippBdzaIIcDOLmSTC1zJUpOYuUtHJQp7aXCJBw3OCLN6Zr4wWDopYPzifPhe1e
tyxv+XxEgwFSG257LlWrKWG6ErW69/CIqIpQ5CAh1vHkTxFemks6n7fqxr48W+rJg+z+0hD72iYO
0WSjxqy2MVMNGiQYa7nnxUo8nn9835fTLextG2kjgP4e/0ycSAP8lCm5o4X35aRErZkZW3QauYGS
+qAmWj7Z7CXzCJpHSiIG1QdH4oVI+TQeSsvNdS7m+Nt7ARTHKSAxCLgEe526Gx2vpm1MhvcwlJXV
fYu4iIErjguskJrLQb+BMp75Oj8ZI5T9l7HDRM7aV/fwfxFXRGmjENfWqXEL+ni1vPk3bl6iaRl+
+l8VJiF8mSDSOBK9ML+CavPXeQR/gOsuVWwNPe9vbbRw29CWIlDlIidv2+i9/klsGoFqK26PgyDq
vTZKCxiyTfBUkzcGqGjRBwCJs+FBbtk19nI352D0N+UGsSyJBoQl12TD8CdjNCmZjKpeAR/s86x+
SIkbKUCL2fO/P5ZJIywD5GywZGu0PISvh+wqiErpGvzJhTgkwTL1zz0MkBzx7DjU2UcKw/4R5MIa
YZXu6mHCsUN1QYlHuPWWBHwXHaw3jqynE8+xrZGvzChoIBfliRzHENtPK+czj/OShxveEH1OWlfQ
Qe1hkRkX9vyjwTje+MNrLidw2JjSNzSCU6o5fYns8bVXClqIHC0Djn6DxazuEkYDUMqHHtyLEpNj
oRW3PPZ5O8de8EM54gXun7qX0UgTG9LQOQVJk4ueAftP/cIVly9rS3dRPFy8NDMHP4r8VM42C7F2
EWK+0nYeE0fP9p0eZ4vTJtRvTR3xkKSLgbLMbslMBu3j5huDj+pc+3XB/ff5u8BN+YgTf2QlXj/D
3plpocuHZh4X4PaMWtjI8xBp5tTOlFGa/RKJO54mzzULgfX6/plWIzZXw0guzTG8kGTTliPbejgZ
OwEXlltmWQGlcHl6ngHM6cKXRnzmeX4uNa6DYWMzuhwtdWaDvBKGKOe1ivx5aeGsd/n+sfGbAfq5
cb8aiNyeeOOqgVDmwhCOB+pg5ZiqTFne5i3WXBW+JFgb9VDYzJEQrV/I1qPHm9AwPNX14+pPkrLw
WeHUYyKh36CGr/e/yrfg+wzh07Mshao+NgJcmtbjBjAlAT//JPZV9lnce6SpqeRrnp+fqmcJERhg
su6sPufk9o/jKw6e2Te3XIqsXMtVvOZBS2FNp8ONlYttT1RgtSg2NlUWaF04hq0Jfdifb6qWGjTT
NMWYdCyVMTtPhPEdhJtoiGycgPJPq426XHDe8CHKSPA7X2R9INKjFvSEXoTLV6vU3caSXNJVBYKb
yHqDgxal1mt4DycVy+nEEm3WImzQu3rUDaySMEW+8XdwUzY4SpgkGTBO60RHbH1Bvi/oWvK4zrZG
K+VW5pv6VENqpLNSSFCilWsmBqYvnKfIj3BArsNTtXUO3jMrpop7ElK1u24YVQ+COpqVGKbyqFRi
qNGF0tC60RXhmZhUiVsEhNuifbbyiSGPOY34B38uJcn96j72WMlqEx7Zo7tUdg4puMX7ljd09v1a
EFuempQK4tU+GfrbnGWUOgXHhaprtvplrcUOjrfEk12S5zUDAgYm/rWdJvayc2BlUGpLj9AAzD4A
Z6OCHBBizANcgny6cFX8oJHVlSEi9XT4CTfxdy3B1YldFKt6JaPi5k+lbUfmXOp/6JTrBjBdYrmN
gMlAtd/It30y/0XXt0l1pvR83CCs7tFkp6/wdjoACMRmjk5GGTzwUIESYrEj5mS3rqeu6wVP21CV
btFUUflAMvvdhs3IEqeuf9qtzgV5T0P7U8MYOeeW2g8nppTarAvp
`pragma protect end_protected

