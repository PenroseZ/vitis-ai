/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
aB5EHAkrB6NT/NTMoBINikqg8EwKYDaK54FjPax2CptnClXJaFSk1P6Y/9u3FWJjIsff+dSOe3bi
iAx0iPp0pZj8xWoo7D2kuRg+plJgYo3eEH77LyOgJ8X7XStkvgjstpA8MmqOdtjObA2+nWfOXV+w
qbssx3RmnSBBdhARD6rqOFwTf7/3cDuK7QTo3GD8GmkOY+DCob0TXNl7kc1BlYaNbdaJok+U9OEg
YjjGCk5uikHjY6JmbT5Bd71P+OPQhQWHoUBkHUIrhbxZIfDop7LhnylOAsOUmH6p7xY7O9pS50TQ
NpvG9Wsvg8pUSyb0Hyecew+1A6TcJyANzCU7xg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="MxahWTeDMTwz2fyFkxR0OEw6OdcfpBcLNutRaEfsJI4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 301152)
`pragma protect data_block
hbfFuBI0Xp74waLCAt9YsBXmHB2xoohavhi7cP3UKSIDh0stRX8YqDx9Bo4FlPJxsfRdN9vKqyUW
CGHhcfQIKgbF2ejABT0lZIGNs6xP3p+q+AoB//n8DhqD5XIncI5fUgbVYKdqZgG2K7nt852TJkQe
2uweZ05qU1aepvD6ogwcuyLTybgVyE7iQqe8vfiMpdygTgvdhVU96b7rkrIHlXwiPBfYcAmnwD/B
PIB/1jCmkHk3E/y7IUnX6dfekC8UqunmDE7P671usmRe625QEB1cVpuq4owZ3XNJi2ZdT73Zhinn
DdKNMLg1ZzALC+qnSnOpmc2f1A+PsZDLmQN5WVCI3ULZmwMVwkGO8X3hOX17WUIa4mT8ctq54HjO
yJKorn1iR0H9jsx/xkyY7G4hZyXkiUxVw5Y4lG+50hu8njx2TCujUImU84PixFfZfllsTLQfKYW0
DBiRire9et2ko7IV+mC57hz51QI8bbIhHrBBRsv/DZEOMe5h/b8+vv9nl/4IryHneFdmUnjOfFoh
2LTnZ4Zssw3wjRzRS4hGOHWuTFO9i6yU+26dlqAFHrTLLmmPOkBeplg3Cbsi2lqhoBndT1kIKrNc
MGGN1+ZXOrMwFnQIwakmT/1M6zZhV4pytfevz0YjFQJifqCbJIsIGClw6Cpq9gVOVg1/+4LAnxXz
SBkgDe5wQGADYFH+c6tAZVjXkZfgn08WkrlWSxEODcHvHeWfec98n3ACA+fwUs7uzmQlhJXQt4M1
AXJPVrkwmmVw6A+EBXoIUVihKBdVELIBLNjndAv0Fc3Kj5CIM9VvcDaT4kwaPihm/yOn8zdk+yfu
4GicLEROVlu7P0MrLqmeV1X3HHG2gd7/kgIDAqjxloP5Nf7YXL3yK7/tfpJluB3o2MQPmQSPSKPS
RPOnRuEw5EWDNcY796UYBpafbZDFq+GJhmZ1UsfFYjG5PSbYjdvoxW4Ys9SmLTm88N/wn2AFBBi0
nvUYcFNG9ArmLx0/2u26dZk/NzOuwiLu5DavCdMLGGdrSUZeKFlKpYUT8YLzx2CgfEbbOEy4wtis
QMZ9RJLlq6+ZwjLZYubHyGIQj/03aj/ijF1sR/qGw5uI0eUk/2VITxlvd1/pMLY7j7Ku/Tuc1pLQ
cv1anppCi1nGnsCFOfRW9Mkm/Kp4VKNNNw+R6IQr01T2nFTs/SE9Hy3nlyHNj8j4Arg969nIfnGK
Nxpkbiyn0mdAUAAwCDRHT1P24p7byFQRZe009LQe5OPG/Kw5BCLKtzskVkOdwzyMvxjqy4M8ZkkB
R4o5eNs3e+LWgxWKx6liWHfoyFX05uQRtfiMBdmzhA9Aqv87Ave3y0yvDwBxKS/ii/Qosz3f17RM
LD6vwA8hSrNVQc63on7QmEikpgxXV5ab2qQC5Npn4A2QPlmZf3vwIoMp0Nz8toWlTPqhHks4ITYp
x+/6OntdbDuIJ93+yqAexpdt2v61lXAPLDlWVGh8QK/i3MIXD3ibkbdx1fqL689NSly7Rli10V9z
krGQVWMyx7Mpe8gedPzdaKylWsNCAVPOah9290I4MdtJslJg+Znni/ilf68nanTZeYZVDZWp/9YT
G06PBYd0Q9HcOEc3Bu3T4X9oEfBZdIj2mUocDIrigGE4elDPK5guuvrFE/Aua5P9KV8eP6d/oS1s
WIqRqMBBsgClCmnw/4iXX5pMAjzTIIBbTQASsND7/aRxxguwkFWrjKUZ2+AnGEy5czVltackVsy4
f8w5eQJS81MkqeKlEhrV9OCeIwOtSNx5JPTl+MaWezcaqCooMVsQBLyzgxYUWJKz1j34+1fCcklk
a6/aU4n8UyoU0nmg0tIePi31rremjE7/9X96EaGDyRJ/MaGRqnROjhgdGrlTGFGjAT6StpRlEdk9
Bcf4LT2H5T7L4vt54zxR/4OjJlFh08fiIwXv27fhg0a9y4ccMRiHl9tc1Z6AsieNqLdHZ2ECK7po
T14APzhg4cytMJ7gKxy0NAIlCqPaX2jFMcWGeVmiFkBqjH/yBAuAA85FCDiGsRxUfi271f6mSLjE
EkyELGiKw4Bg3KadIgkrzJQejw9a2/ID9b4Ogh2uM4LmJpkbeIQ/90nQfhJ+1TvDND2+0HJPAe7F
tR3AIYBj5ccaDzQ9FVaaI73LEKxeC9Rceijr7gLlBOfIbFQoQl5WDFPEul8Yejz5snPwFbo+KJkz
xmBCoDMcg1cq6eYeJ6JTZDfsbrVEbnBQLhPkr7vZPM2ji0AxwZAvMbVhm/KRuqejc6pMmaS4nGA2
8yQ3LYOv4l08HZH2wpnYqXmNkVbhJKbTpLQoLulFvTBHGTYsym1MacFqjkzZGgLbBZYTX4TKbcj6
QM++HuNPHPacHFUS/S4GemeQZ4I96tK3eMtn142Z9qY9NI1u4yL7rjobz2QDivOPqn9zF3Cu9CDm
lCDjUZgevQADvjmP6yetPvwIxVKmZCPwE5ALeKsfSI2lQtigd1r9tZVxM9yLcoPOscpunGZbbIrH
f1OgeU+cY1lP1shbBet1QiquRmDdfgZLxxhZVHZ3357ZAdZjwJ63sNkYlmfNcs9Ze4iXNkl9u9yV
fNfwJLIlHpL34yxmRxjYkSq6GwbJmK31+MXvIkzMVBwzJDTyL1pVydvsaEcvRiEXJ9u7pgvnOuXf
LgH8qw7x4Rsnlr++nhVOYOwsPb4Q4yesEK/ObDfua5TzQTmsNZF08+yXL9M/vHOjuMf4BBPXdQj9
On5UHoppg4sikxWz8qZ+BXQ39MlB1ImkM4Cwto5vmhzUKmpsH7y3zZfOfWbh3tBCcwJsBzCnQIyU
Bj3vdUlTEMG7defPSKolDFamWtmKGTnNfY4HDWedJHT27J94Uo08xaX5gueoOllF4FZp6hrF9KV+
isVmt6dYVQa2p2+vwAG80lfJVnctZf2U2fjqvKPiQL2Zhy+oLtuLK3Oo7vRaVvMc2calWfrxDYBl
w4I5AnLVTE80FkAglp++wH72LTw0W/zg2/JPILRIuydzFfam6vRKcMgk9dJNUEgusdbF12ABYnSs
BYib69Igns/YqfPptCU6m1hh5Cg23emsfUjwtaPbai67UJ8RFHZN7bNKZA+PTbGJ19XqD13+DmqK
/Y+yvMiDz6XLgPJ7979MERzGZbygs44RtkY//0S7vb6lPfyKSs7zSFIEuuqpqFT/KOZFYF0dUCYH
l5gt5wMzjqZxqjwnrma0OfeHaz8pCbtz6O4NVqphb9pDzsTBgeVmMlob51SWj7vFPCoyHhQ9aM6Y
+JkoSqaTJdUZU6JMlgDm7vN2QPuetiMQnnu3KQ8enw32KF527Jnq14VTuCpq2KKm9uB1o7QO2LKy
lShddZj3vQMlHavY1sR6KmzTJhEHfptL78Y2X5n55oy6FTBPKGfdqwa+yHBFLZ0Vr0SJYtUxnB/G
v8KbYUaLm9IXhi1JILpxFy+9i7cpfy0UrqiZGvrm48PfOA5hId2eCQo/XBna60zO/dtmFBEhY0la
o2BykYlZiFHJ8KHWRkutrV9ctlWwcBx8hz3KarxSVHrDSkz/yJvcUJAZMDVjW5hFaGAfW4QnFVPB
/ULsq2ji/Ab8VklOy1nxfwZjhmB4Phks2nNTv+T2cLjEwv0xqbvUFPKxVZ00wPU4VkG6iSQJPAiF
LveoX8twF0zhum43FO0XeDU87m7p4BU3Lyc+kakpm2Rpy5gDiWhhNPr87+4vZUNJb6rRtSGng+rq
kVYp0rivcK8fDeToU9hc7id+UCyB3lHKQG3DJpfEW5+3dpLZm/VioouMBBGZMm+Pwj9g68lYq7oL
nRmq8LtZvR5Is2f5z1rmdN9wuIX+RLguuYe1H8gritSK5u0fdv43btTtD9kGlj5lMP7+okUKvxw6
Abb10fPqFlrJ5rmCZHR3Q30jINDW2h/TCWv9lcN7rMCmcRjnn3e2TLJBG5a5wjP/O3CK+eDJUTwF
glEvdq88oKfozo0G1fVdxBHWGwKIBaVFGQChH0SXwK/4o0E4S+8ppwad2c8vGjrP0Ww0EaMBh8js
fYk+sYu3GA/ndpnoNruv7NGy8fkbtQMUCm7lkXNA1DNyIkx1VMs9ysijilISesmrsM0lM2b151Jd
aKnTcK8N/XvGRGWCIVYwKoSDMFrJQBiONQARBqtiUu+plbmLnIj9D+Id6ZOXpCwHaPG3leLlX5Sr
HcdGHIiItaiNKQxGBfZPhxWX+sVoBCedtzYkIJDivIUP6BO1k3pAa1yAXptCpPLYxJC5H5V63OKy
tUb+l3T8QDTmAO7y05j/rePqDvQMYlqxJ7RZX4d6a2ehHpNmn41XO/F+UNC+Fw4HB4CubdfPV/aD
t8jdJnlt9w06ciKPgn08h3zHCDC6NLiYBHKbs43mGeNCoC2q0yd8M2nbtexdFOjMGex8/CkUIlsI
2OTlmIsrMdXgxq7qzN1ZjT6e2+aunkUZ8mD6KXN3DCc+6i77aYqR7SmRyGNw6o2wI8ZW3obpp//J
3SV4+QpYLlvgdKd1w2GVscAyJsx1KIR+Zpx+0tlNwLT9lVO19g6n62ZPUK9GDnwuJPnTa62AOmKc
h4AHI22RvdhSiErLZOzPtmZvJue89zI1LlsJ9EPDG6u9zEgMwEbO6z1fxpvh8gHfCdCGsnKARvFH
kVaMwjDIWBL8AK7f0H5hf1nDikyvL4xHiGcyZKVWih2yu8JglZItQe4TgyFb+pcngcdhMD3igPlt
v/LLqvpEwLtrzWqIKKyviIt6DoxXMQhk6XRfIbDlSoRnbkSUz6vnYa+BwiAoemCa5iYJsfJ8jx3r
bgdmQXawXBSIydylWTVzIovnu6qB6srXR8jNYsGgXcahdy4woJK54RCfYv9wscHQjDazYl8pwGXc
rO/bO8mUcjr4jS6+OXJDfRcB5P5TpbV3bU00DLzDhSjdo+HrZMDV0xxBAu/4zAwFbuwe+Ai5Dme2
Kam+HZ+CC1DBacNiEOCLPC6rritxXxCofgJ2TimoitrG7/6RMkuv/VkW3B2rP3CY8ZQ8yqXZHMf4
dhwRKJyIWHcYKzwqMw+g1sgVGSZTNyDn0UScScVN3HbwYd8oQ4alki/Gknqhm7CCuJu2I5pVpTin
eeYI9jJax8h4M/0Vg1StO7+D4nEr5ckc10CSmPhosketaEoJ1eQllQf3YdNnLnoK0B2hqEzVEAXS
KtMsqT+PIjnw7FaHD+4/3rY5M9vaw4lmy/yHL3rU+wcwxdMwf9qpWSnghvccRayFEenepLW38z1L
blGi0KA3OxVdL5qJfOR61kw26Qivn4D8f2pHg+rLl8NE09yU/pVECdqLmWGsiGXk9xbJNaWNd7DC
YW2JFDzZXk1WCRUWnvrCtPLgcgfuPLzf5CrtrPtbQ/5gNKvD8WRck3bcKUnCfozA8X4iad7/oQMi
1vybp6OSM3zsRiwIJU/pUjHhuv678Tk9d09mdk7usiFSLdwQ9gXnJIPSWS4lXlTxLDBwWJ/n8PGP
ziw5kfKRN55xiGAono9JMoKPt7v34QflHyAm6nJWzmLCi9tp1+O1/+N4OBfpbiMLhC9ZNTFOcwtA
iM1yCb4xyjCU/5Km0KOVe2fX7El3wfduYYufreSrLMa4joUKIMryGj1X1pe9b8WSZtZk7MfLbx/P
6fbFoBpjfrMQOJ6Oyvqxl2wlEP9pOhCDLfcmZI1ZGNO0RAK4FNxdqpQZJAI71xuhmiRy7NDhNfAk
uE5u9MQ4hfdU6nN4fVxj3aBLWoD85TGWfxIbDcNcHllBtFP4ZfBDs+m+2gUGI2nBErvY3Hc43a0y
SB78m7E2ZS4/Uc3ycwBo+sjkFRBwQpLWJQ0nrFGDSYaV1ec83jXa0DM84oZu2xv1obto7EKkxiIT
ipME9mMm4rGYMTHRNClBR32X1x1jViKKwf+83VSEmz5dkjOgtEa8VNf4BmPUmXM0ypMlz+F8oRCv
Nc4o2/MHdSXbYhHJ425+M3isuusYBnPiFaXKPFNiMks61PXopdpj0porzOIaOecCSsxtRWEDlQqW
uIc0496uVzaALAIsSaTNeLEi7mBpqEW4TuVjSYZP1+AL3PFN3Qc+mqEO8Ug4w/Q9JjrkViRYKMbR
PZYeVx8emcZ2PJCd8smtIt82HI3YIsLlf1XP7eM+EZSdZw0cxiCd48kqRNmfuibjIsDiwuCGq8IE
FN5JRd84BDBqlWmj9Ix0e5MvXJiKPigXNsH9oC8tQgL7hlwVuDqwT9zMmUx7pPuaM9EybXSFRIUq
9z2QjMB28d42GZwKVn8QjuuSisg3vYMEhtQEMv/J7lgMogNemw/bF+lD8ZQIzvHiUCNXl6E2+LNu
EEn8rSQM08Dumsq9/+AwgwCEkd3KYiBh1xDzFunxm78FtLnheG+hXfndsB2xJJYyRy6SaOBXpmm1
y7llZFAMxqqPNfz7Fb8Z0jIwYkf8+Tuumfv/NEiBWeLVn+LXZKRD7QqtJuf1e3NkhYmSZVI7VTkR
7xkHG2XyiKj81cL/54cGxUguu/qf0ti1hqIayGuXMoKNMdPxIVbKzJVsaRYG06+p4Oa6W/w5oNP2
9lYTvjh51o+eyYuP18bkuTX2/pFrBbt+kfmWH7mJnVRwdTohB4r7yKzzHwg4+ld+pfo/5tLrgjiF
uaeZ+H+lk9gfj+jfP92xGlHfuUHZ6zTrWfAaDOCb6zC3ohFvYJW77qvy4piEwj6yUPvgM33J8NK0
pB0dBPleBBOwAbsal5Kkyo0Tr2vb3ArC5EXWf/2YK6jdaBwTD1yuHlQ0Brw/4ninDsyFHyuW1nHg
VkXiw0tvREerPrtxeA01Kh93h2CHh7+FpYAzITj92ssFFfqq5Bjw8iqs6VcMiGPn4xo2XX+HBKYz
Jci6fN90VN+LtRpyrOYAObfhoONPlNxgAzQbBPaWHWOn+rx66D+2SfExnr67TcYA+CDfFxkaaOrJ
45svmv+Bx+zzgGaYoAF1THKpsc+BRgOwcJ9uc0hs6U6Hihyw5JT69F46WnOHR1pzUIjXXMNkNyE0
gLeXC7I36JYS24KZPzT3wPQ0Vj+AD9hzL0Vvg8xKguKAVJxBgXcHjN44nhvb+fYh3XOdG1tWG2jU
fTHP8yp71F4ygtGEmw+G91j+0fONL+G6lKJdWtwkBnvDav5sz0EwbRgiTQg1s4COFEHvy59mv6y9
9kwWIBhPP6arpQxVl/rrlvzliU7ESX8mDXGuCP3zFEXVUSMkzlw9+vYajhh6ljHWklnFReNU50mN
zKXxApJHEjScU1OCGx8rSAG8oGgMhovCCtMH3A5J1MtYAGDjckzxNOsNQlC9ZxFikOO1tD3MOBXf
sFEWoaXx6APg8z6a9MexF3fxliNsZu0YEslXmx6cI8Qxhd9nbRSxLBwvYjd7MOieiFxwe/TakgwS
yfZnMnfvKrQr5XRcqLOD55ycD3CA1Rzt3EOTdurdQDJaibrmTa3UePay02m/+VzzZMXQZY6zPari
NomkqsXIO8AjmgFhoE5GXiYqpcWHplN64SbOtodidwNNAXuIexV9qV629wCGYLcDlCZptC9/VO1a
VndaocC9tyfXyazfFRVPD3j2EuEL2uUY9fa2iBgRWWURDSfRgQMLINdpJO5ShntENnKbeSi6yf/Y
TnVpS812pYYCIaOVn19KG68YXMxeUS3C/PCsYqmjAwXWMvQc+8eHPGMHE7uSOixGBzDEZjXQEnYU
uTYGgCZtbZTSdOrhQEXEfv5obznajdraO7FGApJI3iirS0ZNrQL0y8Z0ZEdvXXHHo8KzPuagVEuc
syuYhIxuDLpZq9PcORXoAQyX/aB2yxnc2MnM4O+YdotIB6w9Q9vXs2/EXOHLwa0DkkN7cEljH6EL
t18Nm9FWQ7OVtGDS+maswGN10M+uI8dh3NKPyHPdgNzR/1T0Bdqcinak3QTm4/7JCUaSnaVajUMq
7j7EBtgAAk+pQm3vKgOFlitb0SCdwvRhhzavwfuUxKRnHuGgME4T1UooD3ISpD9vFyQdOgRqD4Wm
5uaCr0RMQzGV4dPcBkCmll07ryIP82onadOQCUHcH/K/wj8GoYF0eTl487BjuDU/v6hzpHLVLwRR
B2zFLwAoxfp/qY25CXLYYKEjkz0kmDgc2tgmT0vRwxidCYWZqWWjTSfxWZgVqP9QKCJbmqXWGdyg
JbrIMsQPyOU7RFCcYD+yeOWuNlfim13RyhLcgYmFYXyV3Eb1ezb9YXBXmUrPGNxeMYGYKlyrCyiT
VD9GhuFyW4YBQ7jnoqBg6TspMeESOqtUN0jOCliMvBQ2dpr6FLtdNqOvbUBbZ2+27z63MthIBrrj
Hge193dAbn3RvoKge4/lUFWYdfbVpvCDafKWkASTXbe5wzkIB0HPHGGfS9VLWBRj0AkkOkN7QGbi
teCkLc8eexDwBJi04E0km7s+LBxDhoxri9kjv4aF+nDjh5KbZ9EvsfXueDc1JCj5myImKMBlH1Ce
qQNdtVPViptYCbmE10U+5qftcfPmGOHp4nzbFIAyfRvU+butGSvK3fD0YB5PKeeraNw2rIKgZc0w
SX4tKwvozvPfsECH8ukhhKdZzkR6gsNiQkoP4mb0FN20a1cKCW57bcAkkZnH2ExHYpsUDtFEIY/n
FVeeLoghqfB0dPPTUXgZV0KkM2V0wWPjhwIRBRMdu3o33NW4ROKlglukvmKqF9sPEsYm8tZr1hfl
07vQkt+AZUt19/8SldT4fPLKN6JV+KBJHICRG4Vbf/TOdrDvXJqtL7pIbXQ3Rv9uZSaD36KduKn5
1/dqWLX2ycx9dy2xnAFsXOVcrdyOvNdGmseyqORS7S51pU/N+NhPfwHKck0/cPVX7X9JjqkHVCJY
rT4CFhsjYHmJ4eHMSZs9RWPZXhX5ulMZXlAXkek/Zojntpku9x8K2owxI7yHURM/erR3LoIj0KaY
t0gv2kFPugepszaqvzDiD3Ph3fEY+uDnNj8OnW+Lq65mRrCd8+jY7Ru5FyX9EcmyVNmJuGFMtzax
t+B0DfRqRsn6IK1DqwGRly8qYS5cQIfJmXGLPOU3OmIRpJqOThBu7hvXNexqVn/Ri7ZsHJJ0ZXSW
U2aAftE4aSMPI8yUM9EVgZC+uOyyseZ4pGZqPNS+Vapma/MepZYunA2VyTH+XqCg663nrkz7j7CK
twomY9k4Exi9hXwrERogW/AdJ+bRExsA3INO8KqnwhfHTv+OY3GcXN6ynDJ2mI7zmFj+pfz9IfJj
uwpBVvx0gPexKj9yQ5eoaUMz86mvdGbr9VbvIj7cwixTc72d5qO8hEZnXOYcs7JVMkzSE7diHnBG
+4jqO67N+ZSVTvSC0+pVjTPeEm0k/x1CVS8Puqo4XR2L/Tukeamnvwx+cTct2+LuJ6qT6VMM1ldZ
5Wenstp4nWUSNQFM0mM2mngkVmbGfFvFMEOSepNHWq6iRQW1ZR31/a9CYlhI+K8UU2MsohqC2pOH
TmjmNG8SgyW+sTZQQRnOPUJqqExOywP71iqTcrM4XrUIhHPRVUl//cS2e2qI/yIgj8HKg6HAcVkd
Xmr+WKC2Uj1ClXg2WILN1UYnLbgOMpwnh68FyUlKUtBeSjNjOlVnnRWWQLu24kOELgMBX6EQkV3r
gnYzoc3g1B9P9lK4YS+xH2PdcPr6neH/403HTs1BpgKt/NZxJZFLP51J+ZDUKWPNChafNU8bzIcT
K1+Yx0rIdUj43vsoTEaQWc03gLBqwMkwXE5qw+ccK/5u3C6MrkSM6xIMVmp4+MkIlfo+eS6IG78l
Qgg1BBXCG8yKe724tqunb+giMG8plDSuWrju+hoqkymhfns3WUmebrM5raFeZdCTfQtEFnUSNHAO
vfU5Tv2EPr2ZUNGV9I91vjz3KAs+iQ6stdud0IQs4pP66fiqDNWoeXwL6XICw3T8O4cES6M9pC3V
gwVIneVx3K3nEgH67warNa3doUAbS4hPzgtqTIyPQWNr+FPnNIeAzdBhevYpg0BMmHporBU1IJYS
uoc9WnpNKw2hTAYIC9CMgqdcIj2cAH8Je2YrRZKCr9VomvrlCXvJ+HQf1SXt2YftebAvdWo/JmVa
U93YP/aeD1m2SltbcHDQ1p2f19/84M9okDRPkFuP64QZobN6/ek4WUqMEHA55Vz5CIM7EvOchiua
RuXkUssE0NeluLU1Mh+uj2jHvtVpXl8GEhQSUTjeC8bIDh0SPOEGlvgyLQ6sqna5rS3zhZHl7Jgg
tTrbmcluzfGs8LAGyBnCqkTET53Uvxnrxr7/mJKUtUXdesmsEuvpb8kTjRwJHSNJ1agZwrgQBgMm
DZ0ZVuHaYhULWMvIjw2sha29PODUOzQ+8IFkfnPd9q39Cu7D7+sz06cxeiN8mY761i8CePHBfcQL
CTN6t/4Q70N1zMeNbdtoNHGie1yt75rF9jr1n6XEpBa449bvagUJ09aXDWmC9yp40/kCt6pjp62Z
y1A5al8Q10W4Fw7lw/i6q8POMJrfBEeXn9d2TW74r9cHGOWxvdJuYuNda0TtKD91nIIHIDBzI6Y5
+QZ6HIvBtCH6FNkzRr5c5ZUeAgvo5Soj/O30Wunusivph2CpWCC/kX4q8OXq9QkqVFnMDTBnr/+z
XOETKwmZ3AnNKILufjdW5vghvDP+ZMUok4xWhkROTr9sLB60o8JuuEgQwa8umb/AKJZNonk+loGb
xqCpBEMFg/Ig0oGK+0NVYyFHNwQoKRwX3t6i7PLylsI9lnhkDPf6jFnGQThYUoHRx9V69vY++Pwr
iACw8N4pk+ddfvgmRYYPy1NWT2PHfqG/VbMBdL50XPSg7ImcJROPQBfBSTMO5Szuu7w8IXe6cb9A
ITMNH6nbdZ8hedG6kbBAGhNndXGgtnqqa8zVN412WrdzkxTdt4wlruvJi/VHY33g3oU+TbTN2+0B
FvvXqSbIL2yuGH8DgkBSs2AueNubrnZ5l/5ylgsR1CIUdJfB6E20wnBNCMjODIBwTw7oOf7CdYku
NeJ/JvLietX8uwZjTdj2VcFAfIbHmVOMOWLFbNRItFk/rDEpwcrnfOEVrE2pnC3jwUbv/myrqsW8
1dz2tDhxxItNWIiWHxsfzrn4DSkAtBJo8/8FekoiNXOSviOLdPRdWXlaOIkPIQdCQOpKhc9fVFb6
FpmEGEKC4NbwUBvFv4oHQQ2yiSK9aGHBFHwWkwr899qkwjKM2n27G3NGx/Ye0OaGjnKAEEHH8s2x
hNU4KIzfbfSrkyxIwNcQQAYgWbEkBroHC4/1Btv+Jp30LJvq+dB3tRtXBOVFWQ9masmGP8JixCmF
KYKPX8qempMbgbk5PQDhrGGjQFwgOVBQFYhlUEO0crEUTgqM0YE3m16dCQs2MWyzjdFbrmH+7086
fZcTPYLzArk94HsDEuaK5xWJsQ/G/E1iB/8Cg70mjvEn5XR0roBxOD7IO2g7Hw/wvnk9L7DUUoZS
tNUJasuPUoAtCHLnsykZ0Qh0Duexb4JfxUb9fY9OAa0Z6t+S7nOgVI3Ia+JWwiiZCrov4rPnsVkR
RWUDaR8/QH/MFv0WcKF1nVwqff7incXw+qT/MamRezpx6J2eOWxavXGq25LWBgHdsGBzw63TgN01
+yKlcK0D4kCcEnpM9qzmxN8YKePAtczEDjMHfsRaYiRv7tfReYaZc1b6ZIwd+M6qxiRXCCailrZG
l/86b07dl1ZQN4XgLgFG/uE4wgEKX0p5Hi4JgjdzCDVGWGyaypC8oww6WWFYsJlWA7t4r1FSv2RV
g1L2KF6ZhkieOPpCFDzrXscD1tLtwubGilKPGjv8ZlNIfksQl/xxZ6HQ8zcVQ9MhXHtn1GbVu4Gb
hNHBqGoSgrqa3SQMuW2dTb2AJGWh4v1VVQpchTbkxAsX/XOF0cRvvVbWjVKrKcLaE1c/y0OooT4P
9melPeNCGzdxKXOoRIARZ/OXzSzLqogt4j+b3wudx1lXQ9BMsmGyQN+Gr04DtEIeHNCrO125oNc3
wO6Z4ElZ9DpRKrN37EwJ+j/qNsjrI+RW2M0y+k9tctWs626WMm3US6s6BdJ/ARIAoYUkTTFm/nSN
Asd1C3uA08auM7iguh0xdHswCeeR47bUC+pcbAlqm281DxQ5LPGzJiPc4kaUJJ7ZD6ZWDN3Ckxqm
HJSoDbtCtln3pwlfWUjWP3dnrgVGDbpsbz84xOOr5tSnsRr2tIjMglG8rwX8A5/ygzL1DYzyYOcD
djzRoImxRxFij/FQ45EYvST2/RjLMyfgQxonlR2QwPU1CB7tCWYrKW1/9FXdFNpCyklt7keCgVlc
LzrCm40+0YLUnnmnwDVqTDR823SPajwPcCu9Z805wSYsgli4xqJBtgBjk7hD0qljqdDioQ9X8hzs
LOr4eklMiEU5qtpJ67hk1hMg99yAUtbvpfmqktD1cnECv5f80z5oNACK3SeQSg2p+BTUezihpiCd
So/1Dq5d9LMTUdBHmZ6F3Vbi91ppAC08fHGnB4dJiwAIg1dTwurYxf2FwjBIkJJH0vti9ky8F81s
Uw5l3mt5Vggsjv/+XmyJm16TQDmpaVVE2j09XuefcLKoNjWimHgnTMbY4RIXrXCyBt4zWXS1YGtR
ES6eMCK3SGbWq9cX+Dv7aKgVYaV+w46EcQYINBftnYk1UM8LPG1IKek2+3lWfnLopfRYmzLnCvTj
u8Fqo/10RRMYWa6sXSVvsBh484jp+hp7HlZMLP9qkJEGsOxStEpEAJjvHGO5BfKLqDQ3G1cfb2yo
pK4o45/yLCYSC91sMJYVuIZI6WnulS67ZL9yeu97xH7YZSIGRapY18j5HjrjncpyxlUsbkVv245P
g82pQJPaqhHiFVBQw8T8dAl081rg2hsjuzVmlaHUUx5pt0g08sKkP4AgDhitJXKiFZ7OXGCMIETk
TiIRn8U0ic6ze/WjlO2+QaXrbovKRvJMaAjx9IrjwvtrE+UuhdjyudApwrLiuayWeRRAksLegO4T
+36yzGIQMgyytSfQha3pnFt0KYWv5z9kxN4N3mLyCM7L25IoWJZvHY023C2nRRdeUdqcEFj5f8LI
+L0rsm+7N+GXC5uV9139XQYXTx95k4vplt+1WL0/wqbmhNql/tqlNdmbAi5Niap7e/RRs7YVBp3K
EIWsy9u50o32Q2Q49RQPiYU4sRJpo03Big5NKPYxKEp4i87noGzTtYhkYtkTwmRflwDCb89uPyoD
60Ap1u7AcOYE4ixpzBgtqki8BPQzhZJKxvL1Droo41Bj7371qDAQdMRy+PLCFy134JA5VzOCEP/p
7+r652BpMOKV6Z2HvXDVryQk/vWzPf8sFc3PHkC2K4n7vyItJBKOTyH2zeiNFZUmPssXNLlZ97Ns
6F+PcUm1mJy5CuChX8f34Klej0Me92otd7TdacwmVxfQ0UXDwywxOV6zwAVCFbiv9Kdb7BFHzGSd
uN9TIHYffz5E9jfUJA5H4+yms1+vErf/09x6Nwz0RAqfBMICzReAMu94iMmmUYZSPwY+yqseAd3L
j+9sbKd19OucKxUKVi8j/vGEW4uBfVBqVFOKr/LqSCsJHhGjce5nVkwlb50FV6unvYW6cPkrsEJF
hqw8qTf0BwdGMe2ilZtX/EQ1pOW8dUfsWmki2ItibokhYOD4WDXvdZHUsjd0VXOw0/neVDrbLMlx
T+szVyt3xfPPepyiARTOpqbbqEJerIuDX1+2jBIKjBr9pYoRxwtywhkGP3NxRI2wqezkeR1KZVuk
G89jSVFYEd890GWCwzSNpCxd9ZFUUkq8wJIQn3EccrhqCPcLIPtVIOyBvwSkQk4P4baC20q53fef
wkezLSvYLR0PpKDdYWl0LwlOjUAWm9q1xs0EnY4wuvhmK0kjr9R4XcJuQWu7xlTSDcRXRQb9/HEn
g7KkdTpK6KR70CIyWhZwT/rVQaPZlkzAk6O8yZMEYXx2FHnbL6VW0wuSHCOb28Im5IMKO8iTvlod
70+0v1WIbOeyYzDIPdTHDlEUgcj+pW+rv8/v3Y5sy/EQyaWm41RT7Q55VFbi6O1gSndQoaWcPFq9
onO9eJfvMqBze1wfxbcF8P+qD+UrZVcPWYy7xpci+qPwM5HSR1pOOvM4RpotRYssNyhosVT/5rlL
cPNFE2V29baqwJuKY59sYfVGfhXjkW8QRgSSMMmwk9sXZN0MIhD8MjdCAq37L2lfKFb/PuSF/j8y
Unjh1t+T9b/NLtDaYx9UiiNDIDJe0fvdHXfFZoj0y8jvFKEd0F6jPBGVnw7FnDKD5cXSgr7DS0s5
ke9R4NXmx0gd4pdhcb1yp2L2ReGO39ZwOo+ffl+9CAtCV2RFqbiik+RvXjlYANvYNVDephFNfoUe
yirIJKMXKeaCxZhwzTDiH2ltpgAfLKCOrjoWvL2qnhFjW6PemUJTo+NGRZ9DO4STZVFsvZ9amftc
5vLyj+VvoETmWh9AiffKZB9jhcLxH6aZrgw5Yd+w1ekHMutOMd+tc8mTrnEWFyMGLWPKZ2/O7bmC
WWnQYXevF8UjHKUrdcu5+Dce8cBJsZyHAwiBeTw0cXJZDhqzEzz8Zu1R5NU3sZM2NIGKLylTgwR+
lUcJ8bj+sYcfgH9wuAAWk3UlYCldwRkfRtTP8ol2bmG2Eq8UytLDRGimcp8DaFa1SRz3q/F8DYYH
aV2aZJxva4CWHOgswkuS8y/+iOYoc/E+XtEYYDYtuyJzUrrMLZaYQi6hpUxdldV3LKB9I7lWo8E5
QGaM7KoEkK4trSGY/Skvs+qXD50p2QUUeljgo/zKnyJhbTL1gKzZ7c0JNbAYd+eVCnSdTBRK8/hN
6mkaxiHupEXY9YZE3Zgq1lGE741wMqMYhnTiM7dz30/IaedfCEwedquG+zgCDxuTCB847b5Gg3vJ
f3aa4MQNz+FWiq/Zdz/F38kRh7Sq4QQRsv9ftAswxjaQoGbWi/YHwQU5QsO9+buNwBAjlz6cIa1D
1fr3YcVN6gOWY8PrF732nyg33r41Fkv9pOcEhJ1YsRDvltuGiGRQBK1U3nMhXrChvnTjgS1sy42H
DeEvtC+F7Mm22CsW5aW0ga/AfK1ajXh7e+fqCvTCHZjHLwZJeOlsyMGyYHvf3UxrYND6cOd+n3IP
E0VRiWnmPTWMhkhMQ1W48QCDQRkE7mJvzja4tT7hl54gSoyUYWwrrk/pa2vCkLrQEe4xEpZmYLwm
PJG9tQ2AOZeGhGY2cyeFDi0tV9UCiWH+MU5HOfcBvO8lqCjVh9lL+4faC1qXhCJ+gXTHJP/MPfMn
3X//zBNDMkfUzeqgS8upXeza6woDi9NomioB73L5d38LDY4T9d7SMbPt07T1XfRXsgJCHpNmtjcI
VBVh/x9ZiU2Hm7IKXE3G6IDCbksqOi+b5QTNBBMG4DEhix68M/y8l/SXH+1M1zbceluOHn6gLQ9w
i3rj5XmY/bhgpw+KHnpkDao+37RT+NSdxkKc3BrBwyM6aH8iv3+baqjPmDGZeQGzt9aMALzAsoA2
eQWGB0V9PzTSeA8DVyl7VIrE4JUKE35TRPhOdZB99FBkREbMtJ1mMsRJWfhsHa8/rthJl14cLYJX
eZX59TPjUyBeVfsfd25zuxGwc4cSCzL2B92FdixqU3bhcoz4MjY0rx7W7HhwpQzIwBAr3kGVEnSa
kVCsUlVVOEBNsBaUjixCCA5E1kK9QGVd1YTf8D5iymqLdkNwNS1hOC/twCn26+rDIl0Ru3CIji2p
Pz54rlY2fkWDbuX1IcNfk6zm6gykQXQ9jQ4PuFKMq6J3cDJufifhRS4qgfc0KXjOHSYBqsTFLtqY
Yy/KDE1YNPMAgO80iCWpStiCr1mU/iiiOewma9OSHQKyGRGh1TAAt+7u9QguOoGqLIb2t1zaTmq0
mrC0LE4JpbpGlgTbTEQfUgOlBDB+mzydQA/elKSEiQCxa4gtpg2QpJhc2OZPSL2KkSlr1nULShCv
wIqaF+tqUZUnC9F91NFV8JjbzS8J8CjmynB5jC19++HWiY9lseJ/6TKGfuds8gcNhKomWzzeq16K
tNwAqCc47ODU6FX+//tgYBDt0MHQsfI+Y0TdVzZg+HfupjsEUgaYG01wWLlsZiQBiVItyEBOCpB9
v/YUHXk7Q5l3OIDL3EdneZ6hXAYfa9MqG/7KQWgAFfZPjSpgR7W+Rh6fz5dXVAXJUk6Ti1jytz82
Di9enUcCY+P0iDnODY8KXPQM81AG/hXM6SsXHmydE0WYHTi28E53AzCK5rzrfBjwGr7HQnB1fgoG
psHWh8XnNsHbgfUewLz2ts5ArSnLM5IXcqzHzJFureC+OhafQ2mZFrhedeTiZIlTZWwx7S8CHfr8
h8OpDLdBpNbBH432Z+jxRbMb/jCtG2t+nc23tuy+m5s5HM9OHnR9CpzEh7RMOwSMF25WqjB84Bq9
sOtX1dKJ9RfvZ8skEPJwOvBvYh0Tl1OVVF8cRfnqUDD0TNSkb0VRdUExiBThekJYkxXsMmDe9fue
KujTPXn8CUvKgxw9bdEuFtT56sS4vsfqDn1lalEWK40ronIGku+hfqWWo05Igf/chkfwZoORkp0d
FzJZdXZhzF4THBt9SriynxEGX1V11WdDQ1CcyAO1fIkj5WffazfVFL8JYiwLm/d/PA6pOPdmLcqe
Wlf8LFmqT0Nt60z+jtJcNbKqNrARTb30aKBn3JuKiWQYCKx3lAmISeWkhGH5uQPzJt9qf6SsKRjp
KOJP0vzFW548hpiyaEnp/bVBFdGZXQoGpdbZIs8DhfPFh22rZSHAa8eliCAzKjmxD1H9RahYnRYX
tsBWAG6ykzfFno/+sEMv9rjHn7oOWTM1YkRS3aQZSW+S0PxolyEq+VFsv8nvdv7PZqVvw7Ar58l0
gOcKcx0Bdqkw64PhQ7mgiVrqoCiKybEvLtLRwGSHEc1bteRxV/E5b5kalI/9pfNyruaYDJojQKL5
31lTXqueDL15K6m3EvxBA5uJo0hKwqYQkhvc0es12oFZDL4tG84SivKkrXE8aL30eFUNPdrHNKg7
kc50f42FAn78Ox6wS5OH8fGX6U3UT4mHqHKil9phzpTTYfvhVir3vc33KBcSx/FaBg7WEeCVJiuq
sw39bKZf4sygTafb4p8x15NpL0Xr7BHLN3ALegV2oz4ZvyfCej7S9brzng1MtHz+3vLdNDKJmrot
OUwEUJ0mpdn4QCTUzm/hTG21801/ffaccfBr80HE6NGuS7cyNQXGVIklvK47duI2ZjVI0YrM6hYN
kGVR5FLkDGWR1U8QLYty92oBH3otV3XMR5xV5340pyWRXOwFv6EuopM5lX+sOIq519xeWWjOb21l
C75Di4ZY/Ahc4k6Oxy7X0qgHTTF7/yvXXfWU/wNewYT/m/7gktCYvCkM+6bW+IaXJwy1DF1n7bQo
zSge5J7CiBkae+NPLh+rxE+HSxROatTeH3wOCESV8mzk+5qmdOfRIH8U5VDCghPi/UaTASrKfdCi
bVbc2Q7yxH/TsXlx/8pFGYIk0E7HH15V2pIEsQRhRYBwUH5vVOvGsZmnDeFRnasHJdxDh749V11d
quzppbd6S+rKlMuHfsb62Efo8xQsHTIhMhK7HHDmeqGH456znojYtd90EwR9t2Zcziz4NBdOKbNE
0yww9S5VsvmAzHKQOGyw24WZho+4BaOgpIy0BCTSEWIn+1SyZVtGgHdMJ1i9zBMVZD6zbuMZzys0
jkM99rY7vZedx3uyQRrY/JzasLM14N18TW9Cd+r0dNxINow5X+ACpLD5qfCjUBZidbxk2inHEGF7
dU3b3Zxw3pjuQrU495YMNhlSH1qe4UnYdICnXLSZrfDPx0zd+mW71ZOwll08GigOujFej5lYq8zV
8YLN5BMq/aSUuvuPiBx6RrpLisUV94oYWh0xt2P+J4zlNfzQQz/zN2Cy3Og2Fwx4bQsli0swvpjr
JcI16ZhT+VQhn8NqXtSNkFvW0hc7Pr4O+R2Yq3iK3lQjdw2NXG5x3wuisOUx1pM7P/MHg/kB5RfE
BNvYGG7VS8q2Y7Fh1VF9Q7AFYgzhwDQsC4EPc3znGq2ouNzEbqsXhUS4+w3H3NKdwd5qE+H0AW1M
r+gVojtgbrXd9sDtryElfzOcip/yftRhCMg7MucALiMMEptUgMSOEezL/VVH/NSmIDc5UMmemUY5
8Y4KkPez3J2LWJ0elr0pCI9XTBInGv6fMgI4y1PhDCh0eaw3legMTTwgrM/bsyBuufYDBXv5WAWc
MewZY603JPf62h4hEDPHe8GUb0KodeaibJdvFolz2Z6GxnIVqMgovoBNjaqn8kPYDYFueVbcGq32
w4pYW3oCQRFS91BlQ9tOSuVagosvTJknsrKse79qGZoPGEM0hEngVnDo+v8mAqiWOqFOxG3rPUiq
/QKQ53yaNebeUB8W2Dhojx8ZvFKibXiLz4hQBVQ9G7ixKeC15gAyHM0Y/IdXLNQDt26QIobOyHxC
ccNunTsaaXjwvnceCt7g00PJ7/T3+WwVHkx6QDMFtVAEisH4cLXJ5LtJC98Zd4qYkhQ9Eq6TrDZM
CNl2sMjFOfUTN3Zkqg3kCrpUB/AaEi/LWhXcI6BPS8BNWvh/QGKu88CO0NjwP0KxKiKK6HdZmyrJ
LA2KEIa9pR89l3EaGgeloznXDXb0FzH9z8DSkgUSKrtkpNBlhNNjNE5zg0AGN4Y9uSCHD298+riX
qAB6Rq2C4BB/ekGTAuxLSbbOkjxpCY8SvdVWPYD/Qf9pifUOu0EfR64SJC5KzbkOCsz7OKNWn6oP
ZD2gHtAn0UAfwchp7Yrs3Zt3qG6dd+CmJcf0nk8hmuRGHpR75d1xI4Dum7lZd7apRuxUEVjJD/nD
eaH6FJvTYqv5d2hDnNbGqKUMxPMFJsm2BoZkSjoJWQvOqmBKA6jp5dTfvdsS/UumAocEZ6bgx8xi
UfD42lGF5hQgGIQEmGvt+4r3VFlQUrVxYU3FZPv+yr53SWYexN66I9JMRjmzxLcLTWdOKebQO1pO
EJCXXFdHWBbNDw6QBz7Nu1/QF0d1JqJe51RGQZ/cZ0413Q4KHN/ALcfcSzUjgPWLSGX+7ePFep1B
FH2t+IOfWHIMxnk2Oe1T/4ZhoPiWGxP/iRsBohjuQmuQwbSbTvjQVUO3qdJlp5VVHMRFxzNTQywv
rqNKf6djULP2S8dzYyzjzpR1G4SpcN9IhXgIIUifODkwaAyoeQA/m2OQe1nRCvlkE3ffgvSlYvC7
CpY+B1yBoNwuu5PRvrIrV1pTtDm8szTo0DQDsDZkXfYcB64WEKwfMb+0VypJ2LSIVDIJdzNwWT51
t9qLDIA9bS2LosTu2mq6FxyDYw9TdeMA/dQynZ/50kBVnWuwkpN1tNIHfcIw7M8gH89auZxTloGw
DVeqGK8OJwno9XIdxm36/4VDEHHyIfsF5UQNSNmC6tXJgaorJ83hGGHUUg6TKRWxv1y15TqnMwkW
1nhZVSuGIHRHJ6cc5Vk9okPX5AebXswHNp8XfjyNwiHya+NaJ0OQWT+2imm0qZkaw33G0diGrjd2
bSXiDQH/do+6TsRk6OEABCunBxec/2pU26d7+ZSl1urZbhLGW/WuDaKUE7SmqDBbJ7bdbnsuOZdF
bnP3fCwQGRXYinwQTaNs6OBYGA1PNmA2TAcC100g3Y61eyKrg0b3iInntD6DduUHijro445IOCEj
64JiMFBtCoo9A1gDk6fXt0Y3kQeIgWjiCgdsKVxNcJQqLw71JyMRf1jRbqP6mYUe3CbklD8ZFVN7
Sv8piapYBFMKIInNUpXgE3M4crswfS6pwYM63yqFT/B0imuiAQhfRX1CSny0GX10NnGYAgPtXqNr
q4E0R9Sd0OdtbsYtw05JbChNk1n02fVcUF5Udsw8mj8XIib9Wl42LLjOznUeSh1fXxDMQxMylcNZ
VMay21tLzEw94lDNB4NczaAk70+hWa0qQgOqYwZ5fK9FiboKuFxZdXEf+Y2xPZaOdRN/zM68ni7V
pNcsZMF3Q8sXuUmwkjQG6b2cAjUNrCljZIQusljOxWlazdCYJp5FIB3DBfaZyuEBB4Oj0EOexRRu
Py859tTEKNxNindB/FuTzwxJqILsQL5P0/vEBTsd1xCwpYzV+IOavYSJQ43aylb6EdXjtoMYiqYi
48LLcmlOOXKbXk1DoMkPUo7iFR6/prKqH4hXLxN07uAdKVanDAMMJi9k81l8sW/BmACvEk186KVo
EbE2m6rtsLcr5ac1Q+PBOoGy/llem8FU8UdQf4U0G92CGMAEjkuPzlTTKbfuXr7IcO85yD3ByPMu
tmUzWxUzuRD2mhrUNVUZ3zn6YvCpjw277oaGqg8TyepSB0bUaso49/XhydofGfqDznJyU12m2M8H
lACfrHt8Ggm55DGv357mST7ULMvm35d/dk3Lojn9fhphAZFi2ZbvsSs/PtxRTrzBbiP+QIUqtvt9
ZZSfwx1zqgQJEI3TSerugjYMNFq0YzWV+3tnXTuwkCMoT7bVuo8fBghsCkSpGhaxQJ6TKOQma5A/
2BURa4XnWaFilF+kRxjKBt8C4QAJ6c0SEz99vkBDy1yzMdKyHvFqjzfC+wD3prIFdz8wbXv33llU
dVwh5V5DXURFStTZSg+q3mEGfrOtuQKKDbbWwDPI9nNACA876Hum7PE57dZ0BxNvIRwm+H4Y/qxB
4rNqWByl+PDAgEnnVAXkS6DLxGCTQ89u8BoZ3ARESYiybJczMevs9TZiJE/gjltmq2CeNWBNDvV2
cThy74EwegshLLy79SwlNy/hRxnqkEtTBRRiK7ygp+0mzeeYsHVX8eB2mjXZ7idyYvfif9xCAFGj
fevqvr+Dl1Dd0P8QZjw90jTvnaeBQjbxnMb8+IdLOjoWOK+Pl/6/0vKOnhLKA/whQ4pU5MgI/C9m
4ARGzM5G7mEUKLkVGQM7yTr9ob9w/trLAYoyceeVfQlgN26HkQkIbB7O3RRRCRFHX3vzwgghmsiu
2PgG58PkFFSANCKxaFjkRHVTGtt8pK9V15mvo4QgtXLFDFZSPzhyHzyULGdYZ+1rnddwU8tjTzKC
cpCP8O3JxSc6vI2Njno8m4v+g3BRXHXkrKwMnqlt1n2Y9i8T8CPfGQCDQ6VIRW0+BCOT90RPQ8ji
jE9md/wWhM2m2F/WBXltUGPWi2o4/ZHiO2XERArakupkUwH2fcQkCx7FDKBku4qvSCrQJJzxxyUB
Bls3Kso/UaKB02Itib6UXB43whvqxIJIFigt2mVg7xlPFW/vyAYZ22k6c4CcClVlFdMEwQ7608yr
Ud5PImrr63i+ESjkrAGU1BF7nDK3PpquGUIPBWtNKVtaaQolLWcNPrZ1OQpWale14oeIKRd7NzAE
5ei58fFfgcd3bjBZgLcAXrowXZCi6izuJaHQqGz5Qj4oWbmTi3fgT0zWR8/IuJHRIPTo9Uz+wIn/
oDi73lMfzK+BRC0UfkDHFf/Mf9nO3jdpNXOx6BtJG9xr9XgMA0H3s3SWDNf5TolhIvwx1hClBhU3
tPB50lXxJepm8fQHJnGKaVvr6yg1UGesmsx+R+hJXKoGfZLV4KTDp4secTW8qi2jHQIv8JKOdyjP
1bMDEFoTz1060LTgr5zmM6FWzuHuyLlCoOKhF4WdgO2sO3oomYE+gLTwVDh/7qoUTLcHwjll06vG
1ebSseSlyTWs4z3+wqP9xWSh0B5su/EyeATFr8M2eDhZygXnvachXpYjn+SftnJfddP0rr/q+Vq9
uZvHPmrgGi3DQFYGoJZ8JkqiDQclxGvnKS2orV6/IpxqUv6xM1aV0F8FtcJPi39EzMPuHKkJCeDR
p8W8N+Fo+163qdvJUedo3NkYdQtN+nbt8LOUbIO5QMiNFogqwFNK4kHQadjBZZHj+bV+ON51QaG3
iCAeOU3Dfm41mVRu43lsVfwE+5inmqD53Jacx0KuBT7pPoOcKmZdnyspzVGtde5M6ObuHAGxCDBW
rPxVE8Ef3CW/Um/PY67ibyoSgHY/LlhORCOseTVR/v28Vlatwk2kyrOuo8quXBlgcn9JfSBVmweM
fBI7V/O3fyV37swotaIwq/pjjA8y2wH3TE3cCXXw0xUPsQbwmAh7KtdDm9/lZjH2IIAd2+ozGkjQ
1gTEhpCKiH+72ZHy5fmpEB9yEVpwXG+dRpOd+nNhU7Lob87pcMsbT+i945Oz4FkNyEb9bGQIDVgd
wpDvMwfWCgJhJ5yEic0lI1oplrFKobCUyE24mqsgHYpKCc1Hijuq5vQCrJow9V3Wyq+bCXYpkl1U
iU7uYeypfJgHmg1xqi/ZCs/KJfehf7/v+5gdd9ZeQgLwKT7t+BWR9zedauMPuRR0ucRVlYv7tjgz
F++JU/S9A1v0wC9U+5WDT7OQ/KhBBiPn9+lCGA8dNHEMyVu2CZI9KBT7LKjkskgzi0SGEfvlN7YS
uP2uxgBzIcnc8/2FzSChD6Oq2BCRfhUHVGC1BvA1pPREaVhXcOcW97AG9wBXb4rqUg+RhAWCtQAG
yV11B9zHqAIluGh+K+xkkTGQt3qG/YoGDB6MzP9HFiDvuqX2PgPM7fU3B96q2LU836xXGJjdBLYq
59VKayh73+5Hq7gNKGetgX2NaTnQ55xa9YvqJ1+utW0hOTXsJONQ75JElXPlzjktFEeI2CbF8Kks
B70RJnEI0K7GZ4m4M4yT1FnZI6ANceeSrVTm4w3R9RZ4zdUjq7WQuEKydZ9+TYh0pCRndZlwjgGP
kcCyvSqpAsO6eNi4XjiJVDvpNhtS44Ere2Vk0NoVE0KJNPJKV+N/tLtzDoJHQrOywwBxwvXDEmxN
79lo1JACocMv3ddXPDrdlJCAko9Hxeu88b/eP7FG9vT3vJzpfj7I6JR7C86LS83ZSpmCveLJcUXl
LfkTSsOSLcdoY6ZQrrUR2IgUncd+Ve0sQ1djeqsnk6BPLtrRtQpE9LJnZ7I/f87DoGFsQ6dPJ9xN
QSTAj7jNoml11HxicS4YhvI6GULNq6yT3if39ehcUFMrhpJlsze1+415psvAvISFiW2ciPWyZRVh
JmGxI5x7zBP1NeLWH1yCNthDtd8VtoqKuAH6sC5oQ193rScVYD7Z0QA/tE6DFAqhVy7vb/ZWYsHG
FT0oYppNn3vTddRknRKGacPnjRLYAJf22zICpLmASW2TQe7CuFzLJzUYBauU5nU9gvq2Ee99nixn
BcQyGL7Q/AFJw7HKzeh36dcxkDd0TtMBN2U+o/QjBqCamKtJXf/aaw7taBU0fYcqAWfXAx5AsZBC
If7eaKbG1WYtpKkmDGhCaO4cvAfMWmWyqvoLx8u+5ckssrxAidREiaD2f0kWsMLsnR10xAP6g1+4
jPL/86apirwsGca84o4KKrJh7vJ70d5G66IYlqqKPc98/MBxGnO5XfubPvocESLw0GVPinTQn3nD
VDaEK/x2dl6B/3z2KG8ytB+ziG92lLti1bxmlzd7vN8ioB2L6+8igN/7l57jyh5fBZzvG9sSrzt3
vdYyw7OaLt6TcfKJFul6tWOxrcGxdaFJWi2sjUYg4F1KJaP3bwB5J4fhBF2Q8kF2aJZJxYP6111d
vsRcapkCqeOb6CwUxyy1yYPNQSFV764EHsGJlcPM3MQcjvw/2XBrXdumey0ne5pjkrugKIxo1aeq
VxXRkeYlLOwwbBUK3FXM+e6xplDFoM8uxVOfrtOEqvGIZ2bsexydi4ip+povEd0Ki06tRBibxVM2
oeWkrQdRC4/Tt9ro4jwb+e8FYD5thtbeihbsdp7Oc/HR4tUfVFn4QhluomrIjuXG9xdGSfi4eDQK
Sq3+M/zp9JmRX62YA4UQKGVxa4EF5bTf2pGC0nJwoK3fwcyu5FRhtESnTYqL4evKNS7aH/oeHzD9
ZiikmX9ep8ytJ5wGX6lXydMhMa8LbRCTJn1UJyeaRE16oFoNaXcHa16/q65WsT8beJfGo3oxVJBY
bqI6hX9/QAkfflpNDsC8D1G7WioEC1tEyPeoQ2FsRGa3gKOpPvRe4Ux3uChMTh8GBwDXdpTznAW1
ioE2sKbBlHoZ5XAyUYGPdDmA9KC6rbWd7Ux7SIriJzyX3qpMxBpHSX/NnNrBsbA3i6hHeZnt0ma1
UTBUFBoJo6BmgyneYsm3+dS0HUzLeMwsWNBcKiT1KEH6B+X+d2PhLLgGsKbVAF/i2elNo3mViBkM
WNyas8p/dMxTMF6dgyxAA2+iFfkFEZKC7iZvF9S8FKnF6otGf082H8pjIHiRLfyiZXifmLLeDM3O
tUeJv3W23ZtK26qhWDJuk2DsS7Ub44f7ZxCNbCokWiHwucMlza6A31qxiA4X/8Oo3EMICuj9NRZh
pl/exCGkiidsbzwCMfVXJ8yzKrPtAepoZJw1iTsGhE32cke+u72Zz03s8XXiYn/X+WtzzlueJtOq
EoyBQ9fX3Dk/37EzkA5i8dTGEBdths1mKhdQOSt3WWbc9nHcfHk+LTZ4Kor+c/5wlIvtERdMPKrv
mwhsaLo7rhDoDRjNz0i/YL/SbsuAsO7nj9CuAVfnoNCxkDMLwkhQIWENbwMIZXQp6ln0GyhoVsrP
cqWZWX9VSY8nb+pyylxuzVFMTbmhmUzqbjt5DxU407hfCwuRXBHOHoox8LQ7ctkGhsl3ycHrhL0w
PRcn3u6dOsLQkaFAHtI2ZFy2omjj0DRP4WDT0YJJQIBjo42YrBPC5NxunuN41s3qC17u1qXCAy8r
HKWkHbFAKFs8of8jupqCfCypQ6nxmG761GzQZFRQohs5AxFTqpq6dMB0hY3OMOlu+9w5V9LFj0Ra
DazhZtd1f+mlbXsMCFohota4wWEhf/v8XAQZ3kJktCnmGT8Is252PmYj3AZsmL2nbZ7qVTdDoyoY
fZofTEtLzbrboNgKUvce8H5n6J01axq7x79/W185ON7O5oycaHw0GcMU9wh4f1rj/gXXik0I5aZS
EmTLNqoMxKibgNWg507n6PPlhnLmCxVL79pIaYY3Me7Z2CjZsj4th1QaXmPKy7BQiudEUZ5fSZkC
zgikeUkMNN3bYH+vmlxSHlKujJUBisVxnRja5EtBZTabvLwAcwTNeH6DBoRSYLkUB2upXjaLsZvf
Gxk87PM1CYZchOAMcvEEEasuiSfd4kql0I0L8vxXGSBNV7ZrsnYnU9/seTM544WOegbIsyZBc7E7
kT2NEso7helSOYXckfvtfd2070UJEostTURupqmhK/8Wk02q7N/4y6Z0Fyowke2ILwF9QAPNdZnl
/nphaWcCc0I9ahgjr/GR2McaivHvWmx2a8HrFatYhY7LDg7fODj02RwlXkQ6eww3W5LTS0v1KjKz
n6c0QtlJgiKGdppDUZTaYAge2WLcyZUbSITtY3iuMHJwD875arneo09v4VOBlweuc3WYEFc3/4Pv
oCcMaDXJo9S1/4JiSDSrup41xaPIzz5fG3NGlg7aIE2qpA5+nLCvhbrZbiDp1esl+zxOB1Yi1tMh
JmmNn07p2WbJKFwiwKArE0CokT4tMo7Tymgq1nmFOn3+F6aNQW1SO5XPBdDqLzCibx1Ek292jNNW
X5RJM0P4yYRm7WjOR8mekdmBWglNldLGziEgTagzvxSHv8KaiIU5eciY67tEYEiXJ73P+JzD6ubP
OspvVg8DnYyDr8zypJb589XE9aadf09YYs/pqHGeav8elZcV1J8TJ9fnrjlcGXU17TGNtJU5zTmC
nbQ34qraD5uBuN9EjA3XnIFBInKtVz+4v1aY/McPpwJPygVDn4cvEsu8Je+pqORlKdMChn+PRW5t
e1rULXz1x8y65Iy3e07icRS2LFKxrfzbJpCv+wGor7NqmzQUduQNxI13630rmLOr1FXPSDkermf+
9lyA2rh/i7y2Y6xsEND9SYZU92I5V//nloBQFpgX2qVrEoD5BgjDiqmjZbEauefQyQv7yXm5kPdg
0JWNP8dnX6ov67b/ai6V7ePjYv2o2E1RfJoF4ftMKyK/znUSrD0liDBWLkzvDqgJaPcumgpJdXgD
QlWutH+0avIy8dJ4kPH/XHJoboExNL466pCg4UaQMo0tnvUKqCuTUjMJakmSQBUpfMfL0rJdrIkR
c8jJIk7pgNMk26bGU/CEAKPezo0z5lIRgtrWlVRgbhobw9TehSe53kEO6JI98LD6TMpvZgN8BVaT
LItUEShIpvib6/Z6Rr5y3kBXfMm+DkSo6Ad0SLyG484sL4CYu1cKlzTb2wP96DUzwIxcYIA5MnOq
2FXE7qZEB3C6k7k+WaohA1Nvq3j+cctYlBSLn23rDwv4wWIrvdauZXwd6luKJUR98tAF9/fTkzaH
ZtM3IvomcLDtEUoxhnpsQX+wxNNpL05Xfl59pBPgBotQwZyYZj5exb2hEK6gbGTzaFkSLDCcoCT+
qZYokbhGsFD/1Br97MagEt1O2J5YaF1jL89M/I8m35a3dcZSa2FL5ijAo9b0XgXwC4ztGgdkygjZ
oqDQAGRUSG4xYBEqrZeFqJq1u3Bh+BCmq4ls2GdcvxEFxzNeyXWf8UkkVXKrxtSZ8yrRMDOKu8Jb
37aOC4JUuj1yV1XEGVlOwSpOKReKnMIs9JT4+p42yqLEFvQLoXE3QD90CmRJ7taEj19Iclat5o5e
5NquoCW3mbLtazqoCZ4Jg9Z7YFnIf+W6MioY8G6Z8HFuwo1/uTfrDG6RioDStb5EfDhnP/WXmXlg
CPWnklJk02bzJRkfrXErHG6aKTcGt96z1RpTMnpXnGwMLevAPv2FCrDIdeNaYKJKS5jNG+h0BVFf
QPXuTSHiCe+Lf8lJ/R/Ls7pFydDVFy4dZVhqAEakLhG5eBcg93SU88VadZXb3NadSkf4sS7qpLie
vU02CLDp1UA1atyD4Vi2gHqE2o6QG/M6I44ONwI4ni32aP7S4Z8BrxkyKXVKIX7QBtUPh9xhvBd7
fWuM2iy6gOUo2CrosSMQY939q6nq3x65SjYQ1MqfqaICeBzeAm8ANolBwNT4qo/GlTN8i/YPjQjk
fPAtD0f/drQ7S7VKVRpoj0ntKoVlhINp8Plx5JRxicOuzacOs3LF6cyiJNOgMZww765d3kEwDDIC
QUZJTDjYi0TtokfUu6FAuN1cpDDqmrB9YsZlEsI8YdTC5pFSwvlzJMbYkQx8EaRSJIMNlGricLUS
37QW2tLEMCgZNNlWaPQrSxJegxJOO2vsWmTeXucVk0thffbx7vQ6ngvIu8IRga/tN6U76nBJgDxl
/g9Kruu7hITPj3iMvZgYEBaR2SOXu1bWiJ8oXYf2sSwOZI55PGFZ1EbiQ5CJu9VbA4VfYN5LP2QY
YmoovSHFidSSTBfPSyoWztDVsmnNT0R1b1CY9ZQlzMIpVMcQ5sASmhxBbJazTh0HyUwm0uy4Oen3
afwNOHyW2gtB3KE9fnqH4gZwQ33eyIvzIjFFyC+bjmkWBcawitv2aWaIec+LVhwwbv0Ao1d75X1/
dghdu830+7aq/oyOzvIqShDl9Fd6MxPgfAVkgPJtT23o9Fz4Jcgkmt8Gg8V2d66JQfWb6FgV1Osl
g6HF6Ba77Qp2i24rmF6PTh7420kTIa4Inng+r0cGj+kbRFJIp+++/lOe0TVZhwWshL+IBaIojEoU
hF4Y3HX95BFbB+49e22EqOTWvm8u+UjczegDm2nu/TtNYwBIGW+uuqqkafoWH5VUbLv3sEIVaA0f
jxTnTRmx4TO6DWIRys9tCSiA8jgh4EFsI/NbXXWsDbqyOaatzvJhcmCoebkwFNWa/W1EG+0kno/S
APvc+v8hKc1VvCUfFpy5r8NRMtDMZyeoH4wMymrmC45qCXZF97GaeNQslSKggp6op7YL7anZ52Ie
5r+Kr62dVUrfbHYLRCDiMHHIC81rWAU242zapPA/6N6p5rurvrLnVv1awJvWgRE1VWCfkFUrkhg0
61Zq92TLZF1Y228Qt5LZgTJ5nru/953J8J5oTL7fYADr51bwDpsrlt0QPX8BCLjdMGfNStaTRnyI
Kuu1gyvZz8znrCebBOgnV2BY4deqildVtHa5ye/chs79E8hBcq2DtqZeUNW//ES/dvsKYWcmlCYf
Vm5QFDDlYmonRO4JUCki5DS1pLHh1F++V+r09qNC41hUhDCgDd/viYZZSkQDIbqngoH7QOyR7eTN
DqafORbEX16saSNHWpTA3PuKop1W6IetqWzq2kJLr2mjy8KhQnm/zZJxFfmj3x2J7XJfbgykTX17
UlGh3DlX9tAhIAba6p7zBbH0giaDaObwU1ESiDH7rwXIoeGvWUpNejgg9pmhZ/ug9Om/LUem7lMb
WVUNoXZIS5iZGfqFB3K1liyy6Tg32J1mS4fmUbeRoiyHetsBeb8UtpSjXPmQrKpU0jGWDwUNmZFK
PWxeWAsPZ8RT+SpzfYoP89SKiq+gZY5xBGVaF5FevoqzXaYJZGgTAwCW56GfqVc45jFwpFoLivaJ
6LdxrB/M1h4Y19rJZx1Uj70PieaumYMQxoawA+Ip4iJPqDNrAhV1pH8t5mDA2sDgBIO0jmp0/RGu
6wYhutD+62NBXERiUs4ypaujWxwBLQ0zDD0tr/FgbMPN/36syRA3a20NbCBm4DTpVhHI80+D444z
lG3nyf3SycCAKJtac0QiKk8ohf8N/syZhBENV2UzkMpvOz7BbLYBzv5KwmJksMGg/RkgSdqrG5PW
zfgm4JVGKqrTvi/tA6GGKVg0kmdGb1inthsFqYEqDCV1ROJC1t1k4G+1SBA96IYqTf1FneIbf+GJ
6h406QwUpcafHPNKvyahQEjBJiFhqQn/jNQ1mSC4k1oL7Bq7N8nwnqnREvHJvrHsSvV17HeNtphl
TFIbH01RHjbhNkWFNV6i7AVrgT9FxvqjhPj34wAT7FAif3WyyfZnSL3R3l9C/0ZZVAz7HYmadWa1
vaClLRXnfDvuXShsyNjD+UskgrJp+SFXCebnIMPcI4Z/X3N+vqyw/ztkRrjvB5HDqWYfAX3F5wXY
PXcjgIRlTcuCktR0bVgAGvF8KQp0ftrGE8UDlGNdoeyCNUXg1gkOWJb4mB/m9GXqyn/idobMwl2+
0ZYOvv4APZeqk86tAJnNAUgqa68KLALlpEmKhmVh0JverdK/uEGBOgMqhqhwJGm6a4oHvjaKmzHC
XGhHEMfqNsmJsqAi0gYnYBV+BrNxP4KcKQJZWpNK366fvkrASutKbBjtgw3bIBMH/F5ozZdxlrP+
JZJGsuOfmW2CbO/1+vMXH3bgXEoToyUzEjBqDEh4kZJEYf5JtKf9rwB3gyOE4l4odNHr0cxHXYWx
mAQZ7Xpq27Nkl7umsHNIC98zbZYyrhC3h6bAiuHEIEyffCGRpT8SWj5f2a2ijtdloW9Zb+gSBSgT
4w8mab63uNeXgtzkzcCNMelMmciuYWGst0L0e6oPcIDKRFJXOCxVUd6oiU0RjS/2X+1o9JU9y5+/
14UpDKCwLm3C59pHQTDADWl5/y3rdAwIJXogGXgnamLLdhS6YKPTWgiWiaku1ueOD/+T0cCUPxkR
uZvFU+WSskyRC5IvPPV3/aF18zyIvPtlrnsUhU3o9PVdwfemVw8CJDtjs9KPHneo5UxPlqHl6Cmh
7/UOF7mfZ7C1L27OhPWYs8fDGXk1GOCgApRdBgOk2Hbq8rf38blh5ZZQq2VQS2055PHbmeCm5s9S
BDZovq8MEllA+rcpaB3dEwpHckmq5XzPXggp7NyXQTXnjC/4qZuj87+w0URvgESLv5FpvFjhukYe
RZxsegQiJPuA340P2xNKTzZjjkwkqoRa3pjoF4Jj0oRsz+yAkrCg5hAGlynh73JrxkRS93KSpoK0
5QMgrm0USGvPB61scH6GQI1PX98ar62b3BAwcdtQbb0Xs/MQOpYtxTn1uNUKk5ppBJqOg7g96ulC
Zp28VAShFOE4WeID2jOkbVpgY49wbSiOCAsReichqysyA1OyQ0EBuwEpZUyS5hnRFyQ9wJ+ov5u3
USWdmpggIARPcyb2hxs1AXERL0sUrfKDKpKZKXZ17Erfe/faZVpjLJQqyfp1wBE+JC5I/7vQgMXa
SFPeVAKIhzP2+qKXL/w62YQGyKyhpRNV6jnm0kIbv+l+WkCsOeXlGY0LJdv61nNo0uCxhnOVxexo
HdZRMJvKUUt0/djC+L4ahw0Bvies6Z+RpH6F7a9HpoFfx7M5eN8njZqbGthHHeVyhVQWT/+FQ29v
dLzPqNIb3+AHZzECKqnF/GkKge/6CWAszGwM7Srq5hzhpSyuxDOQ2BXt8I9sMDfFXdk5h0AzESXF
Pvx8pkp9fDX0eIpnMMytyBEr5inlbDXi/5g1wApYXe/nMp3VOcJBq5VhaDw4ozXs50GzB+0mApVc
WRTVe1lntPqvTe1EJVsjHzGotgm/vBNfxC/IXA7GNsW7PTGYLYCDFu8Da4iM2ZGXGz/m5X6MI2vQ
dveVFJv2Gm3Ejv5M4N66VkNmRjZdpJXFNH5wHRfhijtX9J9tiTZBeuRs8VAbhrDJ4JDM3haQDy43
hUTh2x3vceJBznu/+3mF6FFEjWa1WUmV/wDVL2uy3cUeoCbd2c+C2Sdo4HH+KcQiUO3CJWyaOYji
+2SGH0Sdh0MCyc3HyQe7oBDfBMax71KZXxGoAwzr4SlJruKngNPBpp2ECLfcWqcnboSzMouHQu14
FG8h3gqa59ARjOYvxIdwVzyKrpSDTF6zBAoNG3GM9TTOfDQpVzYkjBeD5/H3in0+ARpRrrjO8RSw
fIbl2LZB2yfxUO3YvQz4rf+0PbH3YbS8ciO0z/LvrnQ5FIZ8f4YtQqhguopWb2kPWLAHigqon+Qy
bAzw+NBhYBXSnk+cY4CT4ceETWE1k8UDs+qgv/cNrcGg6JpDJvnHSlwXkcYz3oSp7Ro+37WFXddG
fuUdAApZ4fyliVrBkPvAwN6u5YbCD00kpvoM+P/MDsJ76BZh0/EWgh+cjk01rsvP5Q0G69BnMrpr
5EC8RdTT/qazvxa/QVcqzQsn51osvR7LAPU980vEZ024U7t6Q0tKDHdSsyEHuariXgZDkppMMvfI
9GlYAMX6y4VzbLnXBQxwGYF63uC50xxPw2a8y8L705FOHaZYxEl2tEhN2U0kQLsmKLRw3L3oi1yG
FRABKYLXfj/9X7nfwoJsGWa4r8i429hbPor70jk2wN8TvqEHvA2vRLEq8Spx9EbaDhYL8m6N2+BY
TaRSVel2WGCreXn0/eIncLSBoVfZtB3xccWnjbwtLNmRR32uvZgW0fW8mhaYJNgKP0whmtO/a8vc
c0PPMYqImr748GyWmm1Yr98DEFJVnVerZ89vp+j15vL0cP12IoJWfPR8Vha63N5Rwb3KJaFiINrP
k37aEkg2V0cqKYYsA3NYdoFa7LtVI4bPOIlkv6e2P9fFx4GN2UR3vP2qx6vQwAa7BC/hMbj7Edxi
8AYPFLy4iKgNzDdAFczOkQWPqukJUoGRQHJIDCzk4Gckl507aa6o7szgE7Dt+N8rM6xhvVof4jL1
HvCO+6/5Gb1SOIVcbMvkL8eNP7UNIfWF4yt0RtY6gJjafQEeCx2eV1FyDeSqqv7M9BwczN82ZsNm
CUFGb9ge/10Ikxsou4ciiMP0YdvH9SuKkejMt6tcCdIUK2K2j5qWFgosQzYFVIpTNIBK8C1elr0q
zXaJ+DElt7CcWjQPnR4OQ4gyNBN4XzxSVHN/aRTNxMFRmzeGhHLUV0M1t9nYW552NR0H9fH/BsGP
QpMIHv9DpNlFilQRBUA16mx79IcfTAxyiTQmwrpNzZzWnh0WJyDYdPSwremkLYGmmHKWJyDjsZTm
ZncAZaZkFeFB2vCHytkNcxWfOgSiR/1lfb5sAUF2JtQbzXtPJs8As7U9/ndUaIUE3Xk5WWYK2eJB
5AWgla4o0wmwgJvOcLyZeO+7p12X7ze3FFeiOqXr68QDjx0rm/5mLhABQ5fSj48qhCMMkvBZnkut
CwBhHr3Z7GEuX8YsKRnd/zhglVfwvRsBo+Z4Js7vVz/XcW/oHInWkiWhYa07Mg7CGqnYWw08qoxM
ZNMCO4pzKFqEfUzFwt7opttX3ioNFPuD6o5tG7L8t/2obg/t9F7HK+U1vjSYy7D4wGJ90IMQ62uS
XkIFZu76r1u7j4CvXorEkSzvlm0uEwnZ3cMu3gNKGrPI4l2Ep2fROwQTmyTbT4myTylLvoia0N5W
TTucd2dONGWBbIpLb0eaKMTdTjzDy8ejHjCYBJkV1cis9eHfOUrTHnKWXO27L214qpLE446sduXW
cVVdW8JITRC3/QROc52eXORE0xCQe7NX7NHgMamxeFbo48kIGI14vPfXUJ/Ib+ynLp8iXKvAOXNI
DnZgBpx9Qf/caVvYo2SZPcjPdhY3v6e1OY+TsqlYZo1SKb94OGwSFad524Vyyi3R75KDeGLOHEZW
yRkA3uxrHKmZkH6cm6HgIydHUyOdbG52Eno6YuoikWzx9gKkhBGaoLb/J1HCwy/23QiXIkAa1LfX
M8w1SkJ7OrzA8HhxDTfJ++qXOLXYJyfR9VgYW23T0xeTLSGLtKRyj3EK+JStyEVIYFYtnAGzgZn1
JKeIbAvxkS/Q2HgZAxt4Uar4AkOi1KJ3pCsRkotJQH08wuVBYhcS62hpcH/ULksAyw+ome3/Bdia
JxDCtVortFxcbj9DU/3meoQmTsNcMNQmuToSloAAY/WBQJVCgGjpse0SqJU3s7V3NGigqSjMd92h
YNxHqSW/w4HTqEZRjDm+/Pha42p+Kw0hq6UR/R8s35G+sDIZco0Ktg9fBFxfaJO6kXdLgJ35pHJE
7Nlwxg3sgT0X7XxPM4pQSuE5H/kq+96DzlUpMEtay6c/lAqciXyU8asw80rXjnG78sErDtTbHfQI
c9gI+FI1AF26ua2UK0asniCLO0kfiCsz4uDG1Hx3LMoEfOYs3nQrMGXyXfJ9DNNZNpBHLi/ol+p5
TANs/w1cpsA8ItES0RRQBkU6S4kLvAuUplAEYtG50foAs+8oDN6JbIevcY/4lk8unZPweAcpuGQe
n8XwrkLbM4mT4IjbWxW1T2c6/2hB7e6yBVb4WK2k+K4t/oEWQSKtUXIX6+aWSVsazIek1H0AKBsw
ZlY0fQg+PR+cecMTNPNcAUhJPsr/gKyNHYfHnaE+vGMSyJ+m93dnuroyNO79RUrD1rny8llC8YBm
3dTkLbdIywQcep3i8/OOc0LKXEfXv2LEaMBwyC0O/JCrDqQewAt9S86eHFseDUgs6RpKAXnUVePZ
mtcqMynSx+UQg2F567zJNcHbvwdmiJzyL3kaxz6l4saZzaM853X+XlBC5dUy/RIQPHab6tXb8205
gp2iRFULfXlEm2RfVL3HviX2Aj71wVg81UCAD76y6+Xz55zfdFwvq8W0dZMDES20AClRGcKY007Z
s40tpipzbly3xGbuse++/qkvS4LL6LulwmtcXG5HEPPEedcCMaXZcX1pjMu1lCV/tx03cutxe7FC
uYUvpX8aHcxVjbHVlGqHnZ439pDIT4oyQukKXqGs3ZeJRtmKKEiD4PhunOcIMk6ndRPYIypOfbu9
dElQdbo/IBCFAkvCjy6agxG+8nPFlyaeyl26F2Ww4HPFABZ3cH12fauGwH0oTPMLlZtFcQTSYSIB
E1pyjnARFA4yUzKyLwhJlyGbz9wLk5V1G0vHrlSAdAEjnPZzHeQYcYaT7AXCgnevKZi1M+1veOUs
Jwz6xSSRb9JyLI59jOwuSluawr4B25BeBQ+vx062Djq7cGlSh+p4NzSPvCkifYkttfgYXjtbPch2
mlvrIwyl8VDHxIIRxzUzmzWvFtluMVAmAmhNsiQDsFfCoRZ9+RsehUA5vw18MNMYM288YPe8D9tR
dGck6C0ab7Pjgna1ZU8CmfO3wYFx/0c0+ZzgdhiljabcWWUv6khSAcLRa9lpHUBDOkZLs9ogbic5
FLtyQHKEo4Elvszx63AFbSy0vJiwe1iiEJO0BR9IUaNAwaZRCaCkjhA4NWdihT9WU+LDhgEZeawY
kldgHwKjMOH2vYte2SB5fHF/pemtaNqXyrvmdIvZ9aYfQmIsBW0J9NU9+SYW7mpqe6TVjc52K0bB
Ia8eGzsy3xl8Y4h+xNP3VVFal36BLglQSosUmnjzMgZttXxCrF1zeewSi9E5d35LeW9J9nvAjvEJ
eZ8FcWCAc4b6J/WrzLVC0d9IgSgyBqsUMP91BdtXDe7tvFYNrts4mNviuKhW4KKvzSlwi4EIf9vt
CG6B73qixwBn6nkhYAI2iRzB96AGXr2z/vuzSlnp7c7kEgqCV6/Ur8bhfyJ83IDzJOMVrOrP4SnW
jIj+NDE25TH4apyUhhUKxe33K2YlIVDlOSTBLRhaiK63Mv26tXVOeFBo72ZNzmvwJ7llZWYFdpKl
LvBMIcR16Srtuk1Ow6HCtbnFZOxZsyQbf2xV8KZvMmU1Y7T1JQa1sVZ6p+MqXO0A6mGcMNIrjPeq
t0F96rND491EAcElLTQwjtAyxJPhY6GDY5YunyVNpthMI0UiZ/VJGgBpi8O8oZlNLlsuY9jhwcgj
AxU27tJuUycio4/jJJsvXXhJq8e+pXIdYZYwv2Utd7Q+uDyyqWXRRyVTl4C+Aw+ORorwrQg4UeyD
SG1hB48vow+/OUIzX36WdVFd6HDVGCnh6lxU7qbQZQxnxQVGYs2ZZavJh56RYA/GycKNsICFAHLF
kP1K9ifoGxtN1LIcTNw3ICvmnRvO2hbpnf4g9d7wnBhcEtF/1caPXM9tm2R3MI2OoYSe0xZOatYn
5WfyfmfkRDP1QffDkpnTasIgZtKNOedbsi3t0uy9XzhNuoRwR7pAgtZPdM3ZPHPN7NSGEJqRJFtD
lFDWQFSvTHUx0/EUp4CvVXkJmHjPR39VZvZOQAx364Yp0+FFnJcBy9NqPDQPocwVRK/iOp2gXqCK
tFOi7ZO81YqjeYzEVzv/MR02SZLfJlSM8T6U7bkXAsEUb9cUyGYbH2wKtiLNU50mlrCNSWNu8J5b
fJq7iDVqg0FXmzqp1/JAsAfdJOmSdzIeuM6C6SuR+LSZUHmHvaDjYZxdOuX5wSLrYgko60ZYBSmN
sE7kWRwQn5RyVu6/tycw2GrcBkpE2SZb9iXe28aaw4pjxuIFywNIUSVj4NjbjeZ3xmAvHMOh2ONq
w4aQ4OusPJ6L+z3sK6u3gZ/xCmWFJpT0k1Qhi/dPSiw3jVX5m+D8rlDUfGkZWqz+x02Mm2fl4rPX
ZzNY2u0jzkNpFjFaQD0VBEDRt8GPBoukkhe6/kM04hFngJiBN+XEuHznHPYx/5JOnXW+g7XDz3Ng
C/+Fzu3vDl/VhN+VVR4u3845uP5q9ZoqsiFwqjFwyNq22ZHZ7Fe+YJQNh6Yd+CeLUdtBy+sYYEF8
4ni5C5Kvg/aDXiaJzuPcoKHnm7KhOUtkNDo28WIx0q/8J6giXsL11sHTPwgSA/XsV03aREIVbNLq
ZxpQa49iyF3UV5rcnX6dttBD5H/74JP6YEenvZM53+HUvM/z/hOc3P9YXPrcce7G8+EcURQetW+f
BGtSawlciytcV/E0loZdRC9bMABEFihssR0VzVNVrytN/f8lFMRbRjfBr57f8KM11y286v7basIj
WkHuEWU0/j1HuIeKsasF1sh9Yq4jbYOevEZhL0u2h/S4XIOmdKhp3UPROxapw8oINzWkoZFw6AR2
448YhSAVQXHph7j2FQ0CQLOcyI1w7QUpKYnaK96RIpPo7J1FwXlXXk1mtLAOFrGDReGxLYKYhwr4
uF6oWVu1q5u7hvr6tyO1C0uSmuxRDmTLTtC5VPZ2X3/26/ugxj34jqD9MiXEALMdvvyK4HcJ3JRo
BTofJ3MPRdQAAHb4DYw5sPmXox9oS04X0giIYtKoLkY1cFNC6cglOzz5WRbnfpXqcfcRm8rA5pwC
/+0zq3lR9nUrrAkih1RF2Xq2Ts6oFOZX61GLWtNEIrqHmWv1TswQgsl33uE2HbLFj1s2bsyDgp+K
c1Tx5g78OrWWtD1uN/NmHkpXwq/L8frycVyYGDM9QtIyhATJXT2s0O/YPUCZ/crZ40kWXZJwhC0q
GqZUMzXB/PjMCkmD4ov2vFgCHNR1+axQBVG0mVRKbKowvaiZIzcxnhCPJoQ8pPlvDjgNq0iVcNQM
MbNXzedG7StzV4SccKVwUDahM0+ndFFe+Mea+bf7jHRVtIJuX/lBlmQVsC2dVqJbDEF6E80FgqeI
DYSpay+YVl97oYw81dCtveIxDwEVPK+DTAF0EEaWSheyFDQG93om2SICiU/GQ4CVhzLMqPBl8h4S
L339L09E/CvVnzdORTfPxKBUvtuATZ/HIqg/Tio2MXH/s/r1gF1ikO8gxGsJci5YmvebtKTxjPmP
26ab3ChjXJDeoCxeMvDXL9Lhcg5yiGI20TigX1Mgd92ST2L5rdVTeZciENBttVsSPznu8yXcSq8P
bBsweyEQBrhwwGaYfTpDRX9A3eVAIAnAoIrChLV1jf0mxqvhxHgz0nFQdjys29thz+uB53/KBeVi
DF2NBtuKsSWv21hMz2MK6trhdT1x+zSRFw6ESwJRMHkhjFtgersJaC0jEZ5nMzhCmkbRbUeO4iIJ
7h8v0tpUjVX1NBiVJbl9esnKnRH6AO7tTVHQKwqePGB0DwV/LB27Zpx4xNVYtClAQv0t03Ay3gKj
EoqjPcV9GifdKVqbr3+zOFw55J1O6F+hsBvvSialuA7+Adt9gBd+o+jbQ+DleMgg9XiuecG/Hno1
IKIxZGA4pG4wHRRz69/mmqm8ydYXG3weBdLLgzEDOXMzKLe7PVJNtA4NrVdt4Dla/+ycuNKHfK0A
78EyFR4CSUd3NK7oz3k0Opls8xVE1ETZEkZFtb2KU42D4EwrhdcxivP+Cn/4LkDsTFf34CuJ/izF
08ycSzkmATS7RRamDEOJeBNAvfZDyG7GRDPLERpLwTSDbJ6lYo+DDusX2qEwgfsvZbrDjnNJlzH2
RfCyq5IDxFRUWQzMYRyJoqoT9o4L9ZvTklwp9O8kcOdlx5ult87ybiToK2SxiRUhOnScsELjqzZY
G+vgWZH9EZ3XA/bgLCJEIGENBHxkLYzOx5XXiyADDKStsVXh7HCFxfNMFbaMm+fFrIowGJ+1GIG+
xi164+e/GawRmtGJDfSFmSCd6AucjgeFTLvnqLGuTFfsmcVWjek9Dlsl3lOQNGEX290DIOdLkH0F
tH1YfoK3IKeK2jFtnXEF3+3HfEKAc+ELNPpN7kWee5qslZc8mX8uoP0eYQlQbRAEvMwmwyd8UJsn
viQmT4Ym70bKpwxP/R9+nwt0/B80v4ZNDr7wswZeuUGf/pYzgRUAF6PeoGJPi70Y+kqalsQz3C6Z
1Kta9cqNW1HVjY7Yz/Ti5QpHd2i2OG6K/1Iz1naK3WokwbM3KUrV+kHhmeQBeRZFbDLGtSHxMpm9
XxjRGgsTSn99ML+OpqNzEVlzpg4Y8rJcB1MbijkUXV6fIWdt1cIiKvWa8VIITy69uZ0krlYJBDCX
WRKL8iUXQr0KltYDVZiEQ9fedDmh7lRO8YNqKxwsSbnC6ufsR8bEWq37omKCAUJV2MXp71496q56
nfNMErePlnD1SE/0A0qygrsarPUSVchlabmU6pdYl/xcu/Blr7OPLBfcsywhsOsw8j+WSQhAMoBJ
2D2Cw1Tv8b1cFbqYcz1GyvmXCxXuPuk4tHKeCugBfkNBOi9h1bqd7/+4iQ+qCRKgujQDuEXI3hfM
828kj3YDppnIIa3JUdHsesX8EKAIgux8O0INWFj4Wh5omQZWPiveNbdtZFDs4ybyQQQv+nRtCpgx
6tcTn5qxKDOV1nATmjJEYF2fg4CJKT5mLRUNAAFjg1bKTZoq+2YYFRYmGJev1OsszyAeXlDd3RJV
WJQ/LYPS7EuTohdXqvD5cTMCC2p/4DFbVruetI8eUOu9LI/5ONYeywJOK2Kb+nnvPihEVoHqAh+a
8ZOk/Ii9/DGCFIV83rczg1grq76sGLVyXCx8maISvQTVmnOEymyorNMQDDa29MBoprxWi6u8WOwD
r3hWqB8gCsvIpllCTeEL1tAPAStDUm3dv1vbXdo4dPezLkG1KIvwfkmbWYFHH4BDCO7eBWzqCaxH
UZIMxJ/xQJNsXHaU9lOKDpx8NfC1pdCG8MnH+03xE+dBWt+87sBFlMlvsR9qo+G8M8Pz+uJ/lrzA
CgVCdIOUtOjOqZsfObjJUdZUxXEGZckj0wurM42nzmZospdQF5IdB3yYOB4752HZsY4Ss+Fbx2ZF
rTbBuxoJYFMbMJSdK75gXTGyDlX0UP93HrFCuH5pEUrHbQvGC/ZAeJSaP61cBSkJwnFaPunYknyq
uiT8+R1DK3GKlfplwkFGeHdoxycVtn1WVvqBRMWwfDlVcnKhQ6k2IimtNe87P2DlRpdoBBP4F35c
tD5oDfuIpKNij0OgZymBHj2AzLHGu9/ztDpaILm2Z6muDihbOT6/AZaP6VcqkoRl8p0OJv8aIGlt
QE/hsgVbIJDEAyoiaSHZLU9AuxFmEL330z6YZIvje4iEWiYMrmE+xBzLWLQ6F/wIpj4ZauUkdWNb
OrfAggPbBPgg4018tVRRVmcCYS1RQ+wpRfqF2szzZsH0UvCMZe9Ia4ShBk32wX1sequSv0YcjFYm
gXmeS6EZtMpieJbfIFsHuNH/Gbv7+F+xOW/7z1+dQyiVHyu28KEkTqiCBT6yJHf6oM569SJ+Kpjy
XpuHCmFVB1As5gjT+7T/7RdjRV31ICeHhH3fu+lUqB/X1NGAqPJ70PvRLuOAJ2J/T7A3jIGK0SFi
fg5eh3TKZWZlPc/prLVtNvpc8anS9GBzc9fvnQM7KZpDGp+JJxVxb/HbKLTXv/qpixScYlvQE9Mr
XxObVhR3K9f/kZwDfcMNNgypZQBaYZ31m2Fp9VtkZujYqPmhf8rWX7qxtSw9wSQlQBR4xSjcQ5HM
KDyrUciAhwXgamaiN+jkUip3m5XuLfMZSZefYuZJy93me/ac8qAwwLRtcMo4CThlZhouKbQt8wiu
+MLY0EOx499E8++aC1rvntRNr+FxwDL3m6tDrdK4MKQPxbxok58VZbxe3EimnQiw70Rzt3N7wIT+
Jb8/Mr8PD4FGjd+T7VY7HZ2YBU4u+a84FTH46VkJZZAaG8BcYcGQ2q14haQF1i+uwsDDI/Y7wxWP
0tguhH78i6XHkXfeipeBm+XBeezmMu2ZWkFl0joTud9kZMRpOdgejZHUFewJheO/taT28sz0qOtm
CGqVvkMOL9+shCF54p9bynYxJHRgYQQsa8JKWVNFbHUyfFoAu95YtW4kb5Ef1O5+qI310rhee+ah
kk22f/0kJK0DuEv8O+8t6YgILfWUr/G6GQ00dUZes+rb1lHHaGfOZAw1jWNukCvVTBVuwiSsbnmu
CVUHqzhsB0klP3dgPnFFzXAixSFHZXTsGOtvILRECwubzDLX4zVnEdfe/qkxUvHj40kd23tlBxnc
mcjerLVzfuoX4nlfCF4JuDt9cVAbyZ9qL9+AfwUYV/VhR1cwGbqDTJ3adnG2aVZbWV9PU+RqAUwg
eFBEQS9XFCbspTxiYBIF4FdIna1UGScywKQZaKRxpR+sbKeXQBfTsZBSrZYKojZUzfaJ5vIpaQUG
2DW/iZgAkmjyISRIebc03wGk/rq+YIUqNqVzBRK+ZjJ3eNk9b5Gs7eMQcxR+uavgZwEVhMWf/sf1
WH/7lgVsNhx09RevOV8BSLwxykw3sXTQoWNC7PImuVffCPlPOtB5fcC7YIAmLNI+ad0PauM1OgoI
wAyBEFfF9hOLuJtL2A8+RVGQkEloOOByfhyQ7eWj1MVtiR8cQKeKaCSYkvnmPq9YsghCtB0oTmMj
Wte1chT8+SIgyFoL5TqH/ZUA6KOI2xDrVihh2grwZF6uWHh+QKElXms1zh+ulFHM44/jg0gIrRMn
P0J/tVfQ+D8nU8pbh7Y9xHanKplxXghvk6Gn2+s6B7actnwZWhuTmulnd/Yvt270V278D4RzIsL7
Kf42LcLBjz85RUOc7zxJqt20qxXWwJx59ZeJ37b6aUKFYEfTN21xGZQjWFSRlkC4BsnL8YN7t7/m
wZAWrzRqn4Saegokn4+8L00xc4x5yPXTZefg2T7HxaETudTT+RNd50sKF5S44eTBnUuUHMa1uSYF
6tKGa0GfG2wh8ecUeKbYa7Sjorbylw8AuN3MDaZuKnLweVr7bwBFEYhMgBPO9UosLNCepLdoriMA
9/Wc/BaTfgfMw67La1i7+3h/KaH9t3ApGPZNhs0V1s+0/t2LIQIRdp/tgEDZ2F5W0jlloP5EXQJa
TqttVNP/I3USJt/tS0mddqgoYqIJ/mzle4tB/bi0sDrjEuKnKb4P+CGcp0OeJhZTuLGwzppUKsyN
lHTeq/h/rlrI01uTXmm0UCu7zAV2Odg84IcDZfJycWuizXumKtsKvLJ5fLSFc4XA91s5TENn64xt
8RPI2iMThYhEVyfSbkU3cCZ5PGfki5606+yKq3APPHvbnja7k4ijpaBw+5rv9TXiGuy9632tD2vS
hKOjUVLLp12nHJSJriKGnzsLbgNYEgEnMR+UqBAY7y42x1w6oIwbtcsT3aFccba9ErsonqnmSky1
knyvvcuZNCd6ughOUCajZPEJi5h/01ULhlHwp/880l6vQaHpCw1jYZ1EiUfWWyV4p1O1yimIddot
OvDtGNdqXRGkkEIjn74Us8eNsMSs7PmvVfjXngWn0bz0V7lAlpBzjP2VKuZJHyxN5AQ57OVuvPo2
H8RzI1EwcO1uWHPtatwH0y9jv++kxMoARaZuqKzybPIIfUZ1ZmF0ROIkHRa6CvBhF4kGXRaq30r8
MusP5P8cjHwc1VZZz4VKKewThU0m7EIPyxaLzshZgRjtmYcZDaVxLLZzBwLcomj+4PffdX5EnjX1
x95vFwYq1gnbiWEitn/hwAyLEV46pEMQ3pkH0Y3TfFAHA/4vB/9NbK1phxyZAVLLHeUCXi94Eb9l
SaXg95mwyOW+t+x600+BxxX4Jxa3A35aBOlGJUevyJiMjoAoSPDXFNMr8tFnz+nZI9W2R0eOm+YI
rOyMW1YNo3el3LKec4FplFPePJos8LrjQQpFmuQTTmTYGMDkGG94wYn07ZA2FolwHo06WNj/ebBo
sYBFCdYqvO3w7OJEaCzk0whtXchrQbabbQ/UyNbgeSV+AivDqo7cbK5qzyQw6TW7uNbBbatGxiy/
NqzMe3gLumDeHzuT9lyZjP25ccjLkLURguM6rJIaVZWD9AO/Z7G9jOjpvnUFCYLXaKCDaJ64OzW1
jBzp2TWa94q+7lznw6xV4CuBOE1P10KOEYrT4/cBAJJpYCZF4nwvsT4H7TEJg/5LzFY3C2/CO1La
RQ8GnSsCOORYjRdl5StuKrgB+HCQt8v8cSOXqMOcS+PXc4D5EX1/rnb0yyXjcQJE8jW4GwfuNs8F
mVFvMF2Qz+VBY2E679plvPWfByzNFbFck2G5f1BIIqsbVPk1qHufIoQF+CY1oxUr3Gs3ppiabGG1
2yDmQs4HkZvnZbZQ94NO6FvZvG+mw2u4C8R6FrRb8TM6Z2pcTa+dpOg5I46J58u6iz9FFKNjdIZw
MI5Clm/oBk2fYf+mLhUFTwxOooRonIbLvuEd9atLr/w42jrQO+2BSjH2L3xUGEYZ01n8EmOrPyHy
oBl7iBxgGvLTFg8bWq5NrWaAUa1gAlWTRF6eP2nSCyZjxHfEEbIS6u+QDIBQ+dcdI9CcwRa7/dzf
52k67WgJxrYWjGQIWFl/Ju8AjqS6moy58OGvhv4hUZSVRzlzEstbo6ylhjPl2soIVkg4LVc6uYc5
fA4ZCRucOXpqRDDJzwmIC6AypjS30+koko7FMwUv0YRpHeOXyZ3VMoW/7BfJ0y9/cyqDjfm5dFFw
hPXzZvZItUSNMWiq8ySIzYqGPwYibvjq8lr6uz8veRzVtn78VZnTvBs92wHhEPyEloI4TS3KU6SH
6s87DqMqypBQElV//0DYCn/fD/k59LzKZtCEuzhNSyrPtUtPIeCm3vZ3wi7akvgQkG9WNrKGm1SD
vCwL3gT769lekRd2kSWPe9mLnGs/IHdTmtv3j301cy6mFk7/GT6jg/cAYtFBHLwY5MX1XeIF1k+o
t17aoTuaZW1Tiv1jC3V09jsk/Bdak6BIkZfBZ4RTr4uEouSiqfHZXfAW1Fmr/E3RLIVy+UV3Nu8+
Z4EAcVrvxhvSU7bItU/iTa2RVR1VQg7vZwkEQtCoCeCI2vce1oG0Vt0nN2oecSrK5G8SUk8PdjAV
zl09xEZwYcgwfFDcTCdCB7WRTPWYgRukYORyn8uE9xkLpy0IHx+mVWrsBexFvzgJL2kROQpCH4DK
/E9MJFcRZfVv1t3qk/r14UxNLVbou105AyxUxI/pMKGxuxOHcZlMF1hv1M8gdUvLk/f/XAtHfw0e
ZxRNdPyNm8Zk0PBfHuDZKRmR6iO3SV6lybiWsvv63erMfkZtsZG6t5RrfzsNIrasYT6Yh+8YEMye
tcmWgTkbeldN4rj3fAIucGuHbnHnqkReRVdpIaOkmG2eoNGvMRqkKi/UKKNSoroGxWY0JH8NLsQC
r1Ogl47rf7jh7a23OSTmKHysIcudGJ6zsyaPQnOSgv3XOVJg17L0wzZeC4eHbkwE/Im7NzuFi3ML
51qqJjL+gcv60fU5GdHLz2F4Xe9rOkR2HTqJFhAH8F8d2FWyOMY5tMOOM5uegh2F+WSFHB1pHJsh
0ON8LuKft3suDs3Hd71hpQz15j2l2ypKxwkzqKUfwzC8wYjJAsWnkvUeFiYNDKFoV5/GPrWFmW6s
EBchm01u3RSn9/qxr7l+J2LGID1WdmBY0h9GZ718+Io8b0nFlKGAAx79E7sF+3WrCfoAKMhZ/4hs
4qt+xArx5em1nSMSrBjUBkok+j+SN9bPSFAzQsr1SEI7BKPKeGc6u0FGDkNZTGFEdI0jm0TCaMJy
3gdQI19lkHsB4FH7Vh0Z5iuFfPwlCqUpihiv74wM8PTL7oeVJSvi0eTe5RDEzjhlefxYG0R8OckW
wuMgfy2ctvpGdeT8vwEULooYEM7OA+2WFOn2RvGS8mjLMo1uVAYclzxnc7c9I7AOFsvxc6vdGuUB
BDdK23Vr1nk4c3XBQrTgKMuPMDkfp7lL1GeTRrkJUie8HrHUX/n6lAtle08bQrSiwZXBJCLRjDPn
IdrW/4MzKo3Hx1PAJS29H9TyguaZx1ri20F7qq69/LFLgeiATaTa/OIpNSKZHb/NssvXYEPkr/wH
vKtFK8kIdZV4mH6AFgArPa/khTdw2aLLx1nsVhViO8WwWkCx3QrrBPuOLo6GpCHgY//KRp55p/an
SfYSvjCutTyloVlxX8RSrAWd5iGit6UQrpMAx1SkpkA+O4bDfHhgXWfWFa29RTkAnVkezkE5l46q
panYFzdL1gGlGPxTKTn6e3M9eQBvFgKOTrCW0SdqnC0Y5z2rdXntforY6xBI440/2c5y02KMwLSP
mkni2xNJ3qJol+egL1by6/yzQNHf9h98qwH5z2q/o0j6PBTMMGN6NbvhOXsIX2uHFDZvAUt04aws
oKTLcMCMRHDVswOVhKD839RaZOXqpJPFAY82QRTBNu2J7gRCO9czhlWJiyFhYNxcrS7VIIeWffHG
3DFRpHODZykTYxC/YvN1FprVRp3SL1kJeZcn9kbDwWp1d9vIJs+F3DXIgwSJo6P9slPHrg5EaAfh
ALAUUER4CRJ2mnfMcDY+1bdYVlVTY+DEX+0qhhXl6qPKIx9lXQU13Ojd7CPJUznf6tOfneit0sK2
u9t0sh3IVw+Yxr0b9QbAZgrlepsz0mH7zVhyJoJUA9yJg/ILGND8m0hprwlBSCpYyh6g7CbUsB9j
doS984zyOijlicuSEk3XkJyjx2IGMHkONyodb9PfzYSYYrvImP5j0KmsbrAouEgcr52XTBDH2I1x
SUZN7/Nrol0m/t/DiQUoF45EH3h/v7K8jGfY0wPH6lKiugLuUiHUTwUvq+QTNWXtlL3XFx+cTJaC
F5HYmIj/I7A55AuzNuAHpA8r/7RvUO1UjT6qv+6tGrF5ynbST3+Dd+nYAiRQWZbBDqq44CY69Y9O
nfeF9mB3ozNhQh4HzxZNyLUBT6ZcjheAsx8m1QcasdO+cFKDxUY8kjAOoocNR3u6vhZDqcbPOouE
GKXcqk35F8nLGUaje5AQ1pnqFEBy1vJ9lhlXUFBROjdZFeInrNHVraGbZ4DXqb+BXlpgowMbIW0D
6Qt1rTBj8XlNg/r6eXgAujt4fMEMN5Biwl2mB/8/m1hMrku43ZhPynYkT35cNWKnfijwH21NfIKI
0OYZecZkdtoS2hkj1wdykTAHmjpJoaMIeN0SWHuyyqIsBGWQCDbEZVfWsr3piwcTHOAvs+ewAyfg
W34P3z0mGjSoOzcqx38ttYN+uegzQj4BWbcapz2pvYWbwHryrolK4yZERgT5+befSRzPXri79FyO
e0HfTuvvR5QP/9d8jKd6K+aFihIbNMC3Eq6lfPT7txKRFIAXCoQhx2F9+4xIYzsc7M/mAi2oBfnV
ysA6EruFF+wuzsZ8qfJp1OGXaN6edMCfo3RxzsX5k84otAmAQyCYHQ53bnUD2zqGvupaEj647vZL
bWwQVk9WZfGqNgkjC1sdYc0yf4lP0kC5PKOQ57gpNh7X90t/gUapjh8Ag3yrhZlKdah8S11yhwQ5
OEdtqyzaBJXGikYfnLlKRbCY9lGSeuXN7niQ6x7+cTubkcWxJ1FuD7pXVCdXopWxjqq7KOu5su7s
o5Dgkv1xM3Z5mKehZMSkCTCx8tPU5mDXFoOtOec5Tr6RVv4QDwNPCwIcGezElQmlIDcm8r04tNuy
gCisxZVZXOiu99t7WCr727nkg3RfMLRQdZznTGbY4ClXrbFLLABOTf++aJusSfoZBoidK1HY0wvF
sRqW6gObM9nWZ3EW//m1YThH+rjxf4h/5+EnJoV7Ona5epsCwVACgjmImyWKGBcN4xrr+bvzUwU2
Sb/YLfVIC7lTCpcIXSmRsFU0JaLAm1g6HbW9IOvtphrRFf533n6RU7S4jBVbTX5l2mCOM09DSZVj
GvwIe9H7OuQUuNQfSQRlJBFvYHmrcrTXU4IeLv3pzg3ql0jmIG0iZnq4rxYuvbueLGxkdrg5NMUN
AM3k60/WzIV/lNACMuRzcwmp/+66nY/M2SP4XhDlPJT8yN54eMIURXFYYb1gghFot/jOZUZtDJf1
bUoWUWlH8AP0rKXooQG86FsSXYjGtBJ4C4vElJFe3S1pcxRR+IF3vfa4TW5V6rXplvzr9nJnTbOZ
i3R4orLEJzhu7b2LwJF79BA7ymwXk8FsEDqDDnFZFsK/dv2hdSjvWhSaFeBKXATmffQdhXObDGoa
cYRBH0zRIm9TQGIXHpXNQSRRb2AFMdbyy6ZCmnbnMeR2X55oG6YoAClVOyyhDI+AvCYDJ1DEc/ym
xOuM+jddz9EUw9Qo625CDyDh3CRy/KKFFXynJPw9GAX/ieFaMBXvLoOh1UK8r10oKEoXqwzchrPO
ZjV0LdRPR4c/FxvukDGV27BlVMWL/fvim2EZgiD4rU6ez1dZq8s2vog9BjuecgcLJqA42wLioZii
QW5Hcbh3lhahhTgcLXtKLYmxFPXQZtajzlOorFtKmmv1FHNeltZ1GcswJMJJ10JVPAyTpWnokf/x
ok2lfK2tsKOqv6WaNy7xKAqoLQc3jby7rZPECzP1uUENxtywxKNMAipTBUEDCm7jThln0rWfOKuC
WMxAnyIf0KY+Lo26P4ABQ0Ae2vxqrjx4l9HCA4kQ4eI9cCnBIrBHJCxgSN5COePzz9Q23Szow4yF
IeiDR1OvFsdppFv9bdq0TRFijuOS5opqXFz6OJcBP5wbaNDWDBriCVgyVANkuhNfYRoEQaD+EK98
L/eR8xQ/aK3aoxhD3bfedBx7dRwm57kkW6cCX5gfeFtJKzOED0wT4l4kLKQnGfkW1bpt8DhPBwUS
zZYp8UhJ7V764iQtnJYhL0F6yaqnlF8MRyUKljxWdE3I4B0mAZeHjJktvfYkS9axid2pjm1W4kVy
JX5GjlWLNQZEWzdOWGqVwq+dHYeHOVNFMdyOnISPV68DrqQKpXRP4vvVNT91mLaCxC+JR7z/YX75
uc9c26mos6m+mNNLbpuwVhTylJVnx13tq/l56rq7ioX4b4MWvfZLX/aiknHPOcARtvh8rg2EsIAE
RybeF/Qp3xIlrD0NC95K4GEPEAfce0dcnJPx+qLUQ2AqrB6qOQRk+CTSA3KgLukzu2OiGULr7Nok
J1mHwbv2A0tpVvTcAxwcA3Uo/ZHxKVDT5RqojUsX+sr5m+dM7ux3QMbqafGxsspPsKjSC7gUrX1t
UAGy6V1Rsrm8zFLpwfvV2TvMhlH+1hbFHc9BLdmSfzAZ7O3gKQ6Ss+aTlFDkKrteDJtfXhlpqln6
u0UBuNbKv12VUtFXdaN+NpuNaHlgIafFh8TAKaymEkvk9teUBoVU7o1gYMtUMeKLmiv4HsrERalj
Mf3pl2afkKM2aClZq3BSLYpmlnspVWsBnp1SHVI12iXl9uotFGoOPDQAynjEoN9S058zAFBRkElj
s10e0g0DZWLtxroBjOOmVEeXZUrXb7VZcByevJHvzZS6r1ATzhLJyewJNSpb6CTre0MUwo5a0afa
jk5kts2gkdHJ/3cheDow7mKaQUy1ddJljL8ZlR7vc2eSV8/8vLXSpPoJH6pqWwZstvY1jpuWtSUy
sQQA8wKWUjUg3yGbOzJBxNANUwYS5eYP/X4YAcS9HEoypTwaTZb1u62D3hiS8nUX68NKayLfUapr
VT0lsAr6e3GQvhplFp6NOV+gYT6JEn5PzwhSyNgJVuQLJQOT53Nff/hN2jC5vyA2zs2fMbbxR/qS
SBlXDCl1PFhrlzd9MMD7vZnhD58Jg4xOoiUeTy+xOGfP/oeuzApQOTYolyItqxEOxJXkdpCduzFu
gG+fiDWcVXNsQoghrk8b/X04XVcx15XJqu+vhQv4C7CIsq6Aw8g9bV2NETjNKVTZsPzMMTY3tuwB
lTakIsvnDfJxk1oZ3vnZ+rHiO8YdBYBfH6anHXYqHf/lGK0S+ZlW3B9U26P1bZGMdKgCyeZWQLNp
O2rVobX/6MnJAXwKbh/Ewj03r8AimM2nXOFar+rJqlWbb5zhWm+fsPkwqRAxQCsr2WX1RtyG8W2t
jb9MfbK8c3tx1P9B8A+VJdzw8RaAYMZkGJzKerUBTmFvCJRMtulHBLaxyFt05lSjYSzZ8H0JCqxu
CbOtn9YuoPrkaUVdruOI6d7qhY3CTXQYa4AdUbHzGahADmtEIH1aWyb8JU2nYcutpsJh8q2vLkgL
478jEdE/GyVrFh7WRoXhTeQysN4UPx2Y1MktTu1Bm25Oxg9PM5mCpWf9Q+QzWd3Mi3jRS6OyVdQF
RYq3JsMntKsXvtFcPSBXZ2iez1qjE/y4yOPEoYb5m4pqcgqh2SsieCIJ46j97SZPcm0a3p+ZF5Wy
FnXg6w+FM96P2/luZV9Gk9fGqe0nFiyUnyidYyAl7aNAW+a5859+G6Z+FDmXQ3l2Yvg3fQ1KDlls
F6N2pVVuG0H6jd5PzHmRkZoB7DDOkka1u5+Seu5OWCQWt8P+PWOTXWw5nRzpSqG3c7lEGSBRR7on
bKQindWZwhIieQKeRsfMNJKS6vEfqNGrb+C9S/aQj3LAb45LjLOvzXfgeoE4a3wPVYj7xvUPpyje
pc+3fihjSJ4SRVMoxvBuIBT0pNCcmwQacY3xF5iARHg8jixS1CbjBmxm9m7xX7JE3N27F1gccqQo
I2W1LpiXxlnSloyiFmkMT+SkmxkVdfzZYsLkMtrY9T23FHvopqWQUZ4JKT4rcMb6eZD3rp15M2aJ
maJUYNgOUBhmTYX7MJR450tlyhfP5Q1PVaEy1LNt61BJsfjnawOAN/52f3iU4bWA+/8l8FwhAaVc
qgVRfTXt9W/jor8tw5UhuWMqFRAtZtjbqFjwQRZXlwgd4Eir/DcMjdOYEhVyIwxFjDLGZGYeyF0L
DXwrxbAA3FD1GfeHFhYouJ8NhSHHFhzmGH7+ymV+f4LdRkMz65lQ8m6/GaxSu07yNQKN+ofpETCP
e4dYJBtWEeRjsLfwxAYO0eOUmz6zToeGuszoAkkGrF966Dt8oIqXzDPbcw5cNWEoO8pTUohA8KeP
D72Sffy1VMDk66ygB8jhEihnRoAwaqP/vv5ZFpqiZD7LG2VmkhgB/89l1LVkcbbgtgh+ilEnyF0a
hj7yaSF+gJqdWIMAmwsSzX39vrjOFd4MwL+AHI5mBr+r/SRXK1QUYPEkKOVTBwkdLpzXTmD7hKF6
Z+QLQ2/kHDLG9bK1jEpAf+vhp6O8nTXaWRroLQnB8IMj5droQ2ZjcuTVPI9oGAzqStBj2VbM6x5Z
SEl56d2gSK5cDz+B+BOtZzq5wvRvyGTDGiIeruVOBLTo88hNjNQ/CsDFzWnkHiSJEiFxtV863f71
V2dl6t+x2wSCZNeip4vrWVWVX+N+XcPmxROcWb0sDveWjPWn/XtPhuqN3Z3P9SSlWyTEVn7ia6J3
1sbJVFegraxvSvBnqfUlUNCR8faHTjhUoqmXKxilaTZuPKzRM4qD/Z9SeKREW4hPYZ5S8SKEDNzS
NkuWr4UZ1TUvc9jctrnZHHHz2K5YMLJVjANc/MhykI+6JJ2NNUJMPTrA+H5FHSiEw/21GdSApjAJ
UjjeO8RRJc0f3qohhBHNpQzBkNvSii7En1+e2CjuSDfDWFp2ttYJY8/amx9eMWBWd02MK3hYRVIj
XzF5T39OxbaxIWgx3WQ1b5UepLy2HkkuqXNogHrkgKh9yIOhuQCa/HWE9SvPBZcTCmCCiUmA53zr
eZRtSb+gLZrI2RwObTtGJ2MTwSRHcwxPxnEkmUlfDpqGnddg0ibVibz3XrP/UhDGV47BojFj5W7F
554UqMzHqZnoju1wTRAcO+I9EuWIT3QwOGD/+V0VP3w2mIDjmX7ULC1+p60Tmj1Mq5BA2Wa1nlnS
hRPzjWhFOx0jkPDescqEchkun7qsvz01soVA5o9hltPIR8rg+df8UiFz4GuLa0vsksLmz27UXvkm
VWqIk0AtWUuZjtQMx4P0b7soAzSdhAZnlws8Ljb38Cjrz0q94lITfFBGsItM1I1IRkVhKUz6cZYw
GvwL71t74pr3G9Xal0iZIk+kDbsVX7TyLjl071xXBDUV6XdyWH3HzirQ7qfKAGgW9VAZlZJxLkuL
4P0nNcqw6iRRBwyNHXGSCK7h8wdpewxPN89H7ebbXtNZhKRuhD5vGfyzjBdE8JcnoCkRCKQCr1Ny
Vpt5x+MpE1L2XBlGumJb1boYeLsd+VjmIbL2BpHzGfPf8giwWNWvjnu+NsiTVGwTr+2c2VtIU9EF
N8/8OEVYas/EJW8sFNipszJ8+ZLIGC7x9KJfc5I61Hg2quUTKs/k+m03xnzJxYwYSuZ2QHV2GGGk
GG3vudchl4TecsuHRYJDqZi5T3U+SsbdM/bHN5pHf2LW2+JK1+QDvHWlrT+pw0FUJ6DMJxTu/Gn1
NcKZ5OybabFW7orMNfhM7t7onaIbM3QiQZWct4Zqqc8cJM6oEiYnSBiyCw0MjMFY37BvhlPpW8Do
w5XOuiw8CuyJdkYk4c8KeNtFbLE7Ua89c+NOWl37u/bxUnekD6xSVdDX42C4cx+kkhLu5IBm34j9
69quiaUAYye1iWJrrV2WhjrFApChrNhtCvN3iQtIMEWV8RsdMBHt4+0EhTx2s7gtDelu2aMX17QK
GCj+jjyzq4AlAUYLXadMqVIVEFS0pH/cFITYde8vuoO9SLdWc/SC99zc7M9wgkDthV6KWwtgbS59
1IjSgydRA5LoyhEKPTtY09Pu1X62hwn02bd11V6x83GUiSUSmoPjejF4VRl/we84YO3Sy3fZOrSS
pc1SB0CcNmbEBrCkC/yXXl+l4U9o5IfDa4NUcWw2/zz9dYt354YzQVPiZ8M396XLQdfvmQiA4aLr
hgPHWoAwaEKsJ6ypN3/ja2r5NgJFUA6ecgpoeT6TwMloRXV1IqUjTfQHtX88fc36Ls5sSDQfaszD
dUM1m0B40kjQe6WAgLzcpCtoegGok7YWmSZokIT3roSLmvpLb3GannP4J6fpaddrZxjNmv8kuIJz
BdYOd2/0sIkSSIUozSZSmrNUyfnnQio/8cbisB4Ltz0JnmKaYxcH4c13YluMObZXBmE+SYu/Jqvc
GMwZA7MJEXf/B0hfL1DAtqHLeBhE+hATGIPOZYZRQZbBfiMHbdmCXhXC5f1FUnWtnAd+L9BDsQGb
jjWmZk5zifUZ0QIoX/PtiQNbJqrNP5fRUtg9JTqLlLi78sxdCTENbAMJUUgsEqFgyd7TKZiUFi+s
VA/7bfBuGCM/MYfM93Mjjm68iZlDBQUBg1TbSSQoLHd26hXgHzwEAUIalFhnrop8OBqjTyRRs5w1
1FT7RXaNp1Y0N6zJqpQNvRtKskf6I2yqFytr0B52Lu1iGM0MMpEZk/CKhgmou0MhtyzDZYivXA1p
sPg/f+f0opC2IetjBVhd8e3ppMZtQGc0Gb5gEZ32qnmsI1VEXUF/zAc8j8VOvHE1E2UQcSwb7hiF
QRVneVbuBZuPc7+5/YnnyFHbC684exkyook/bEAzwMbp6jeRhG5e7Gw5qoIm8crrqw91gBZ9HixC
n0Tg3kaL/WASAYDLcikan01r95ToDhu1JXzrDNTNrjKJrcCWwdorD8p1mdSf5ZgL3hCCpD9iRu/I
7js763hqYFxELPsWspf844PXLEbzLdkKwZfWcu/+TtS/fp8ZIx9x/VjynMMjCgrfgeDfhrE7HWCJ
1wY2kjvR6l1mbV9ktq8qkNOhVtAlzAxiXspth1WuXVkStWPHyNRBq1ORAnFdSzBofAkO5Q9eAgEV
PeF0TtDn4/CQeFJvtWdLmLTpaDLWigMwaqiLJVOGPuuiXkLOwu6c681N5LWeU7zpCkY0kkjIeXAu
tRDJrRr64xHqrKuq/ny/KaxnzRZOEbJEMDBsR3ZveDZlx5nLiD96Q9SwtgTaUQsc3uFswpv3GVNR
Jo62cuFr7xBn3psGgo4OgfVIzDinNHvALQzOm+S8HWvvhPJ8AUwUwCyRkAgmL+IZX6gEjBsKGW4s
4VcskpDXguxS0mHSj2C42h9ZfTsb6OKRi1ufi0RBroE/Ek8ZZGxq74i3NupQWIhrdm3PZV0dVl8j
tX7EYDrk706rOos0RsDDNgb2cimAOByDVfARnwOxjsvqP5QX2z9gK3uB5QdZmXFErU+Rc2rqodGz
Ny3TmUDlxss5+q1ZehSYtkPg9qC91rDzc9bqj3ZKdP9ZxKB1CJtwdxrTHg5HbBUPiATKI3OlrpMC
kM3ZsDWlvNgitMRmehODr6HZYWppRUpqlKmwHyxQad4C6uixMfXOYJLdxJRsrRSLOC1QkT8+t68K
mBdD1ePHQMKrRtSjv8mi2tlM3tKW2cEXQYfFnvp1ELkf11lyhBI3AjEm3GXBpz2UOXw//vYucd8m
dQO+ZpB0KgzGGAJW0qxNw538qLLjQ93Fwa6f6Tdj2hrAxrVVUCfmYn7dOUSkyUv2wg4JONvHyO/z
1ruUnEUGW/iFGaSaKw0Z+YEhMhpsMvNlngBNM9TQz0VEAMV0kR1YkgFO1EVk/c1mXsUXTBRaxj/T
6lzYeGBaVJ6ceNDmhcSJa5mdx2Kxp4bk0QIwSZN+f8h+vGyLWHj/z1o04EnVJOXYb8/xjWY8DgLp
rdPN6SaDhpaNX2Tk8t8ulaDAmEnit1rSTzRk3tEQvUOOhIKCaUA5bQL4vcoyyotiTj60CY1FR4yw
BYxXVuOuHEvSIfTo9z2P0OC1qan5nEalhaMJeUOsfdcTL5h9Zy36pa+Cj8FVD7DslgCD4G5GOnuK
qKKlvPaowNMPbPrjWg5hmIHA7D7zk3TQRvBxopPKK+t0tivuKkjogI6t51e6QAvw5h7RI0QV3e6m
NmpBz7QxQrb1yJb/M8JCSQdeRPur7FdnAgCEK3/d+vV3kkeSHD6SWzYjVWpj5Jpsasvqmx5iZxM5
0iYIVcYJJhEbO0Tcs1FssRgxx+FrfwtIW1zrXVpY6yGKcdk4xWuZ1XKJ3LL6L9s0dzcb3LDZxIh3
gGDRfHbI8kjlc0smE5F6Xmd2xX9yUyQf6pVNVH8dLNqX2aDDl6W7AG/PKolOmGvzMhVBYX9DobrL
Is9AqaTcYcuOZrBJnJv8kTRAg+JTEsHhWLzFO07709mRaaUDAkECT38xBdyMpY+rqXSC6yVgVqeH
XFgMIo23L8U+BYCujOjn1liCtNLw/lvCemfkHWPWaEl/aJ+9SK6BeCmksEQ2iz9h7y3bNQfgUejm
4N8CJxprYCoIzZBiHD2BhmB9XEfF9i8nNZrt/2yTObD2oQosGHyeMp3TXgnjAJGpfU8G3jiBN/R3
zojpKGoW15Yv8cLoKiEIVsh3KpcSHMl2LFAZHW5P1M4DleURacoyFmxcHarTKtW+w075OUBXkpsJ
tGRa1aKPf88v5xNeO+CvaB7YfknNA1JBWaBsuOphRK50/veHWh+ctFZiHiTuTEDT5YzEUY8EpTRM
CJINHgfH9LL0yvsKz0vQnPd9jbFScLs26K9YI4pTG6OgKIpS4YULJEQw/93lAymp6jT/CnDcfORW
PTGj0PpMhJBZnBW++/SvnFeg5Cqf0YafIlSMUhAx+gL0IcWJNcKFn2Kl/0n7Cg+CIdZlfcdxFiTy
Ly++smwRAKfbsDjdke1RXqWIPM3//eOHn73n7tT81w8fkrjlsebqQLUa9z/hWCU34h7cq5SjuSXm
fzyxEkmoa8OIXt9hBvxGz0rGRAazN/UuBnni+OvK3P+96z6dsK+cchB5hjpnDmgFz7LoUoSQuxSx
owCPbLWo/OSEwWfm9RGul6KYCaQ+lUCkz06kc31ZZ/NSb0092hfhGVImn/11h3Gywk19Lv2lyo0Q
FCiLok944MzSdz6C6HM25uyWIak/ku8rJv7efl6YRXzSCZCIu0nwq6fHqzz7eECQbVH9BJWJwXff
3epCTBnLVKZQspK1zCVeNBkJgkH1+WImr0x7mSgzPbTljyI18l0oiOth2Y+9917pLA+nJSW+FBlj
RDESi8ItgpsWfZo+1aEeiIopdP9fGghZFPc9e2217gO5VyjP3qap94sHwAHaiEemrsYsOYRLni5O
QzEYVEnQmUrIngYXAqAu0iE3VECi5bgi9iYnGgpmWcG29O6zMbzDbMdHTSYUmRLcsBtBbNuiqYDJ
PCWviRzatA6qrVL99k5h47PeBRqaHDsI6mHucS1ncizjcEzZrlBScM53I8Tfcab34w6YQlEvnIY4
XsoIC+R/yl63EUU5wr1W/2N78xvkugXUWg/RvwG72nRBNheNmkB0oQp8dfo05NPa4tHhyFc8C6fA
Y3RQbmPX3KLTncKBFrwTWpBwicHoxdoPHare/yKlJNeAoheuWHyu87k2lmDtFniFY2Sd8PA0b3EX
XdE0HTTEFLkH0ngQsUGrNfBWk27xBLV1eR4fyr3VN08PjdvKbspmz4hFfAMAZSJE9T1XhEFsDhLx
FsYvwE/HuiYf15bPJa1WxQFAF6ePmMZuNqZGSKVh0J25Wf/ScNDmSoYubZIBHmm2ceEKd+oh98Sq
2Iog9fSq7VWlF20zZcay+7p2g/tYZIZKgMeyYInC37uhxG340gvOcCMg23nwzpj006+AeQKh16hf
vDTA2CpSt13P1cN5rkS53FiaBBup6GDG8PmQvP4HZTbelXMQ5SIJHn/3mQ+3uU+at0Mjf6rnPFGl
zUxwFIusaBg5dI1pzdgVD8XU7F1hHC0t06jrnN8TsR9KsIa4eaOAO838tOTeIu0DDcigz81xkGpB
0x+MecABawwTY/tARXRs5jDbR996FGbQO4Afxke1uIK72NHSB4teR8E9ZaRT2t+FmR2C3ckXy94m
2zpEouRquBzZ3p+hcVBsIFAuVgTMrTb9Q/vUEOv+2+Kw7Vq+7D25jbOJXbrxuFbuzbE1nh4jcEtt
RYd7G5fBCiY//ngT7j8nDV1pV/l0HcwTBBKrLUO6nVrf/RKXEXo3WdoKbZdt6KOhN14brELE+GDn
BJrIGpfwyd4bpaB23Rsgvu1Tw45gsV03jZyNwQ6ingPgv58fpnmA9o4V4jxBrcDNc1ZlITGdY9UA
gHjvtLXj8WFo+j3Qflmk7gOHYz2KHL9KOhEZnKnRCSdAuk6igTlJiu/kod4tpUTaNlMsu2zcb9zA
1vho5ByXkWqIpqeuzBYwhaIGYCal/ceziDsKLW41+aHHuTUFmeoNZbfEXit6pBY4RbsQn1/pogcZ
k2MDifabT4Z64JPRo+rBcWZQhi/Qji1nOIb5ayt2vKsXGuT0jp5kanCSSpZa+N25bq+TzsBZrxOE
6fcoxVPSAHQML3KgocVCB5kzfevuf1XPjBLnaax5hUYYrDYJdHkMevBTqDnYE3KgggWZ7PIWik1C
sIxxZQTLD9MiXKcGsRmtv2h0KEdB3A/BsKm+IAobB6AuBrinARybgwBlcXu6em/8qgo0kFIdq3tU
UHVJN+mn4yzcSTEoPDDeCvtRfizaCQzhSQW0BhAWZku/crhmQYR7jjo77LZTYpNrZhuZ6wuMtxqV
TFygUK6wu1oRLOTQrsc5r7hpECyKWbbsvvoc0Z9cZay2nsm+K9UXzbnZMGrGybSF9IFGIw69TYed
N14daNTzbks/J2PcHya2sUCOcfsxBwkNi7Lpg3RZjxQBzANSBs297oTaW90vXn9wOpcBZyReiPeq
r77QNK1FTpeQb+tQPqWbfkIyMyVaybTRslQ3oa1TICCpEkb38rZGxTBFId5ibC726oq3RUH5A7jp
EVWCwyEOx6SpAdj/1rcBPN1+jtybFRDzbeccD06jBZ4Zr1NJC0nlLK0LbOqd4stC9q5DeDlUDD4E
z4rizm2n+IAOBe1cz4GDbDYyENU85/RsDrB1mUCSId7XGuQGlT09pLS+OwrrmQgkEQtJai6j+LgA
KRU+RHbN4JupMTzK/AWzicibY39DtUXwCj/WbEa8vT6xnAanjrT7uol2w0BVVa4MNI0c7/FZTL9Y
eP7VW4GjxB0cmRevSasq5b7Uqf4j3BJVH708/Z3/uBt/3XDZmUBQjA0nEgjrs7axdZgBI0CbSgnU
oJ6AzAjgbLT8oRxl4RPyuMCGBXLP2DfZwvyAPFcmppc8T4KBUGA8AsR3q5mHLm/45aUuZW8jwSQF
1y12PO5LICzA/keW17dFCqBT05MuawngE0XBCBhI/YiS8Bsk9MpzTBclDie338vxtF5ubBPtERqW
l6TvJvytt+wNmqqAzjyC0irPEnD34AgMR0IfR/qdxV3FhYikcgM2Sai3wKL+VUyW3hFU5di7eFmr
lrTG9SskTpuQ4SMjCGig6FvUwEVF40AvP/4u2eilqH3TnO3vYvwQG2LSjp4J3bQ6WBu0Q/pF6hef
9c5kxce5W9tCF4K+I1CXnn8voBRBz9XUwYzLyW9DXoktfEymMLTkmkazoCs1Bm4sKC1X6+ehK3DE
KOZsdMTKAxee0hOxEoSXUgN+gkKMFaj89UOG7eSErQWq1e1YXQYxRme6P65mvhk3UceVajUlXkQe
J7Hfhpf/q+OLXzQcDTyTBO2gaw+RSn8rJnhYysVByquYiR/3dEH6kxYgONPRFBBLBtCPO+dk416w
t4tD5JgsLjWi+Vl5gtQgghptsh5/eA7Tq/RUGBQZoPft5vG0DnXNnCSeWXYWoft7gltGrNvTCUw6
PfZVaXrJ/eUmIjpE4NHerkWrs3KRkfrFqVPhPkv74y77s/3T1DTJn1cuMOJJorxKx0h/1HVNG8XD
KgHRAYHZTScf2/KHUCj6I+1Yxk/jQORdlQHaEk4i0kL66Lmox31AdGavEIYkMNH70ebJusUTWd7s
BtUR5EvBoEayYnCfVorFNnZHpXsX6sGWzEAkTwrdaFAseFsiAwCrjocIIxN3KyzSnvptF+SXGdFB
ilFlcRcpYlOIM4VKdig5cwn8vz+SWGSaYp8dA6EYD5qmEuuo60Uby6Md42CsM0o0YPt9EWrPmc3j
MuQRE34MsXbTM6zfGshvI5JKy2zp6nmtSAVzagUL8nCYKmTTCZlZ1w8MYg419ycTNO220SMAA4Yg
tICC+zpxq7YZ5CqljGYre2m0hm0oaJwvnZuAtQ/PoROnAAtLKuk5zu3oX8O0tkGYHxxC0w/dVaq7
JihIky1RfeEVrDYLRGCJ434CkvYYilLXZh9TqYlirJlH72kQOFYN4Z5fc6EK2Ore1B7jhn7UFp58
Bc8XGTecAHWllqWZM6vAMZomnR0e3/ykS+45MpdUrUWNeBckW2mcLIv+UA3Lsq7YoTZq1A4GFMcY
cTAPG2JkAQtBktDRLBwAbxUS8iVhvMELXy26q/sHMOv4OlLEivw2N/Hpq0zJOYy+mlE4PWnex0a3
rXzCtSQXXLjVL0nolz2pt2gTt9IYDzY3ChY1hjdF/nYQeknrIvgufixLwnQ8KxAOfSlZwgMklePJ
KgYkXJBExhqkNWkn2ySCT9arXdBD3dw3jl1wofuX2LgoKbg2PmUZ1gdkNE6x6qyJbL8IOGT/KwdV
MuIjSndTk/sSNoLAQJU5BLezgOgnfvdg6bcSxlDODgpH3ig2HsJ+TZo37I4uNxZ9IVZSDuKYqhH4
/WCaYpxQ5lweMR3RGfevZcRyiUSbSYqeNH1g1KGntx7TgD/L+7lHViYicC6b1Hjxvi/TDcQIAr7x
nuZCO7axPb3LJZt2Omm1+tcPCM6bC9kJVUthqX+ZMq748Aqx5GPRJQLlJnGbMQTiejBvrH6XGPEE
jnK/lq8nbElB9orY72qHvqihKRMkIzyQU5FZ5NJsXZkUcXrj7iENj/z5/SCbuWfRrNn5NDK/WQpP
Q1cQL8nt2SjG2DoWP5Id/OcQeJB9JDR/NW4aL+37G5VOMz6TPb3IRH1/3jsYQevdOSKXdW7bvLxI
GFOorSpSYA3M7+tkTcwgePvC6SkTYGyX3xqHa94aFG8reoZN6H8UI6uttcoaUjo0ENRoixFEkpcO
JkgiIe/s7dU1dfGYu1Lsq9FlUd6NZhdJ8Qi3+n0ivn7KyskS0e+jXij/lcn7SEI72N+FQXkxgQ5n
70SofiWgfBy41AqkLonO4/J51wXwmN0ZaPItWRbeYPDAFnazRqAb02brlG8QiBsf2v33wtDiO39l
2W+7uCNrjU/M5B5qOlHUu08TlWNj8QyhfdURw6WXL/v+FbanQAyk1JCid+pSU+pUhpfQgUxiHMA8
NlaKmqu99DW7DiNf+co4g1zqoLPq79gooJTWQ/br+cqOkfyZFfhplH+oVNJkcz95jpk5lBiIpWtl
M3t+6OiimftMXjRa30Z6PvL4E4N4Y+Uoo7yml3br3dgNAB53Iq1TkdzXsmzyFFsrc5Hwz4I5mNPc
Vl2/h0DZ9iEOjhkDztJgW8o4dnxBolUT9OLBdD2J3bzOjbt1YpsbenZIWHYVrTiONVSAzgZOBqfK
GXjwi4Bufe8SUAo1zgq4ghqST3Kz7I0Gq3shMpmyTEHAWsa3nFi91EjUd1/f7YCz52rFRLJ2lCx1
PUZigdI7FwYu1f7zXapIBQAhkqUsXpzadcbOtiWdB7kbITI/DOOAV7fGCt+3egpxlt+qQQo4HvDD
nnShdeRiq8Wiz/3InOcpM6fsxRn1r8DgC/PZ9/yDXz7kQ2zL96FYLIY+0WyU9/gRVlRFZgwGEg5e
EYOtazuvn9lpaO4AB0ex+ZlvCB+EWTik8ZzT+WbBDLaT9OK1dcCTu/rEOw/AmxfUU1F6VvjCeheU
e76cAsIf94eTvdeu9OcIrdjqW9N/QOzjTPBoebD9YORDr9cLIaz+G+4HRZWVUZPVPMS1S7aayPxw
kmsbqwndWjoGfZCWWPl2oOuNlPv/MP4GQfsQ3vJRgBDnAzLgInvjZiN8ynUTXy0zPzBrphLBH1WP
Netutx8Qf6IrNRvJP26hDLuOTQF2UDleikPQzH7XjktVlZS3BLoipgF4OdO6SgFVNWw+m10Y7SdU
Gth36NNvu1K/3A2N78GOjhYhXDzGB98A6r/mdgk7V+RiPMqgD0QfXn+5RqneEE/LnPWYVs9lfwxK
1WsWq0iV990NBUjASFvnWSuKhlgAxx4xEyjie/dbJweE90kVloxkZUqCgR83L3eIf2YqPoQQ/cy4
ieguwlK++PK40DKhkt6zFu9z2sF32YDpO9NrpHQgUu+RT2wYWzaq5+yFQ6JzC16nUzgNqa6GqLwT
rNvgJ8vcRbGeXnTeMmptOAWjuxI4/v54Y+j4HxR7Avkmw6WJTIGcH3OvakKyo379qItzAKkZaiKE
c5dxc1bgpTgtcgmDknU7Li2TiMM1SkXfG609rYO1A2m0TCi9gwKgsqWrnSqMZ2vZ/smtWEC2Hh48
elZshWN2oLdZ6j7TawMmTIw4LB7RtFrhmPQMvUfc1Meqyuir1Ny7LSxfeboHxbogC50Ie0fSxUVh
i7EckDgLMP+pNeVZLATiS4GxhBMVmV969wHJXBUvM01SS55iXL08IV03GvcdVE7to8gFGiNGnVu4
PI1m7ISE2gB4I3BG0rirDhDXJ7O18c7m7prtj2ahqHCyNhCgt2lZcHa6+aQ0L9kLcCGc9+I0Rs72
EKauv0U1l2GVn3fR5v9uDJD4aLobNrgs5x9CxuyhDe75q8O30JfTJMDgy9Q9nrmlZIxGp3/CJm6m
sLXl3WiIUB2FBNkGr4TMADAN4v23A9KhAiI+2JSix4QGf37cx0/RRTYDKb1MGg9ghdnH7Ke5Rf2F
xJMOc2+PEvDylWWgE56TvYxbb4Z2Cx9Z92/EoXm2xmI+jfBKWVsFf8lVZbECT6JewWvbdd+C5IKu
D+KiXtZqlEvJ3VjfUdzREMEaYPfpp3msOCJzI5AZo9vBVn+iIhuYmfZK+as07w3gKdi6qCin8aEo
10lLibuK3l781szswZ7IJ6hErOHUi/hbc5B+FKdK5WEN3hJRisafj8YSUI9iJi0QFPAr0lcvRsMl
S+MSg5TAEYQUgc2MYkwPo4fHUGCxaT0Rl8Temt/G+TlTK4TBo6aauGBjJiDutLpz9nUVo87ZqFWx
4SORQWEozJavvlg1UUng7T+FGe30z3vkuSwCtm+qeO8GIkln/neNM4+fd9bDwnpf/2VxhzYfBP+P
AsRkn9bLubaEOaE7Wfce9VhAEolsrNnkb74X/RhQXf40xmogTUtOamj1yTOiLMnTd4IzpaMTvOyY
z+h01x9f1skcjaibgd9gyAnI031Ml3YxWerzH/8n9yF0pqj6NkpeE2Dw2ervyzO19fm2W6ogzYHD
7LOJQ3O9pbZM/FQKM85DIyrzFAKE/DfuMpDgD3gneA5N6hmjsE44PQoe99YfP6p6dlaf7BQGHvSC
YmjJ/2UJcxOegD6PocwsI9bsLqYrhYX2AhH0ynkM/lgUnwZ/cxiS/+djswlUUo0w9dJ+i14+78n/
O5SV7bNPgNFsd0yIzIymGvTJrCGaM/Fq8RXAwWHUKFL32s5g/JZeNgcReaOqrC8ROZ8t5Xici7CW
AdHR5jqCuzTmY/JVOwcdst5C7+8RLBkGgOCqPf/NJI+k80LYu95kDixk5JCiMyavZwuYSYgPRnVO
t4ZZrbv4Ue1yzkXuP/N+UqkVIqBfxgx5rM4NIBb6K9vj8+GhSQnnLv+KH5fp8CxPhe+C/ZsspZMU
qNWIYDOq3opoJevv6Jbr9lKkkw2It3nqu+WPfHDo0nwlt0NOjH+/lWUA2p7GbPJuy3uv7kPu/CpC
h56H6EBRrI5QDmp5/0rmyVrMVFSuyiDxmqUWe1+pIhkvdtdXUqTR0v0ryLW+5ayjkM7MDNezZRey
A89jwA297pmSeB0aNE2vUM8WCxelkFNC+YCaBD0/FA81p8/pghcFxM/29iaXQSwGhmCW2F4Xi/5C
q3jOWElZmKuyn0bTYrahAice7Czyd9NTQx+gwQiSnuM08Gg+EisBu0f2EiB6PqAJMagwo4bMzEiG
f1nGwcnPkfozCyFYzP1cOVd144LztyZhZOf4u+zk1vPdz54Ym+BfOwVTewFox9N98YTptza4uNtn
9tGAEDPKSOqohFCUBPok6Tq83N7PgG99L4G93T8+6UHXKxJ3GtoLpBA//YOKUGywe8xCCSaooBIc
9xP/nto5dh+GwLiOUhs8ZsrqFPKLshpuOw3oYSxSktHMxHmu4vpCf8QO/GZzPanMSYU/BlAEVuQ0
dXudsHg/0fE+eNvT1+1OadVAVrYbImUtgEA5zVW6fcunhlg26nc5h8bkkOh25mznFHyZj4Te7YG8
ivHIqwlvkq8Ua/Ukn1VLhi/rZm8AaLY7qq62V8HVakRnjdxctPij/Qhwmdqngx8PGUhRYzEibXoy
XpsF6A9YgLJiF8VdqYErKYuL+wRIWZ+5vzzOoyb11cqZ8hY9chqmWRFqAxYFzC6sKA5ai8wtnVtB
3pNG14WgHPs5bi3dngZszHzWNxSjqLLmhnF+8GiS+psHi44L+RXAZhkVDwMBtSWxar8Mw2nyplK+
oKvgETHQ0GDgtuM8IV1tLXrsEC1i45K2jem/hTXJkRtyDUNq6Pl0B+Y9G79xiUDZr/XVixl6bThd
9CM1oPOV2TArUIGoGrqq+KH3U4552CSNxTOECLqzSdG+GaOd06plmD5bZmgr4+pCh0fYXrLmekI/
t4ltZctkMNt2MDyI+gSZGPCnckfyE4/tZmzgxEXZ2efcpEerUR7hG7C3cSpAQkVhoPOKrm28EnVs
dP01VpG91lDKlAM2myNto84eGC6iFWM+Km+8RjRlmTPt1aBsXkQmG6Gge7GAX7HFcYMlgR5V4xnA
7H/dgUTD/HuIMNnrdXQyJfSPGkhTFxJCN6xC1GTSY3ZkdcSWQkoVdOzMiH6r4lAp6Qp9iCBYS/i0
pLUtjYJTHn/cjUsZ4opjF0MjTMSzWcBDh7BdBG1bbWt7j6DY2j6HQueg+aw40KKwARatIxK6KgZY
hmS7tL7BRk9Mzx6BaCq1T+6Grszgvp4g0KaUjJvNkxPYfZ8xNTsg/v6bi50NyzQZLncdcTu+zetZ
I5LDriP0rbvqS0JZ8ctczPUDA9obRYLQln252ieuwHvLBTekMEkLdy/qBcQ/FFqG9lDb1CGHOuzf
DpcyzVq8k8RulXbtUOI3Q22sImgpTnz63Qa43EcDryE4Y2FQQwEqbVxqr4xfDYhktmc/Fi87rJKA
IBSi4IMjllU5vyxsZkOdtYXdgsXxaQnQ52YeJuSOrI0I70PzNuJnZDbaDzm5Z7jIVyQpv6OOMO27
3/fRjy/DUdfqBL0YzPrlgIfLQ9Vj8sAC7y3MXNoa6CDvTnGL2wVzihtf3tlaMYAry9zFEk1nVzz7
qypJPsQV0+WnnFPKOzEsKXfy2D2D+zOAp1UuxWCs1Vbjw3dqYD3cgXeRKKLdPK8N5DKTeVORMu24
4lMfsBQ4104DWWAMBx/tAwG23GxxgvgWcLXgE0DAz8Mki/oHeH6AUZYtp6itDlKVhbGVFHrrAs4w
Yf4ALdsMWslcLUnspFAdUZ2aIWEWhph3U0r5/5uGwbQQ/QD1nu4DC7/vFHwvEYMr8fQJuLyRtI6N
jThpB26oEOZNWfqevRh25q9+44E8IHi2fUWFBLWExMSKEkX5oNWL9jnulQFdQhpK84QI3pE43spK
gBr0S227n7PPxiJco0dv0lXGSBXUjFiL+H0yBeBI9DB8S+GM4Qlo65xt5fqO4wPJaHSUMyiOIr4x
QDnsz4fGe9NTrp1hbbNuzqNW49/mNmaJj9fMHkXP16BLRLXUfQy9hCCdQl+0Q2lJJRuEes9dNyZs
aovLRPQ7abMC6fnTiUbTxzBSkYkI1itIkuEHoub9z5E+xAtqD0F6PO2H4t1mEihaVSZdxWApqvbR
UYV7mBmeE/wKUS+cetMCT+DKNVMbeld59dAXOhs4jTyD1Yks61zDhrJnIVaVfNTWv2pxXq1byLBc
JhUWaT7S91wiMt9czkXCttm978qeoZZPyPbVgc2ttIDa1HmDrfwDtp7K/d9O9SD8boYCityYUDCX
xGV/z6rNGyyC5xOCR4AdvQKCj65qZoUhEbwieKs/oMO1ls30dm//aEIrPf3KVsYbj8CPZajiftIl
/m6doYUNKaq8TAna0slxtSONAkAwQqkpmSLt1REAVWFK0bA3GKAY/QCuP8QEiv3/ulPb+7ZIno+z
GJK61Tkobs4Ag3Qb1GTM26PUlqHuO6HZE69fBMeyGwEWHvIJcDdRJ7vkk1umXFJ0xJefqPWm4zoy
ghDpxNAC4Soc2/sglygp5YYhU51t9nr6929vxiGGV2dIVK+jy8aH4ixn/3fPMG7GlJFTRPdljYxi
g7an+wfGCoOQab5bah0kaH5r6yg77ITlrQN93KV2JNZqskupfyhFz8V2UL7ENk0+gffXTsf3G8xL
qwePqRvF/dJV1lF+8OB9vt/aZx0O8C4W0JcN3ryby0cFI/m2dfz1Pcya7sesTyxap7gw048VJHkK
Ec3U3OMci85UAXDTRuNAKOiJtvh8Km2l75sLBlnH6/HuY4hfgj0qz+axL3JzJxQrDsfvO5xLDafW
DAZw2ExGEarEoaHDGdggvbT6w7PMmZwMngXCDPGFPHcZgfhLDmrPjWzIuTjgacW7qeuVX3so/1gM
0CUcYnUZscwtBZJmneC4rf5zqOG+jBlHvy16GvCJ5kgiIQEbjJVtOkz38aUere95E75G1T8tHjIp
y1KckO+/M6dTFtpkVqGccA35OpqThvDgAebeg8+OehKi7xtVo+KSPy3pLQGDlqOuw0otJxOUtoyR
8C/jHCsmTiRT4dZ450BiDESyk8fSaZdFatbdKQQhurUu5/R2X4PBgixsQkCcl2AWT8n1y8CfKAan
y+ZvSRZuadnjdjHRsVlevbTncoqjkI89/F7yZmH9/iVGKmq1eBO08/A8PHjHEowEuv+QP7ggA/C7
WR9ZeS4/3S7EVhYN9adMgFTDwF0JZTTAEyHFG/NuH2dvelwt1RG5Nf6mI/pMxlONmyNLRuOW0VpU
J26ukcLM/YE8HmEtwbBlCcAtUxBsRvQduh+wqQ4ydnk20TvEQ0ioMWzB4ULzAiYMMEMm6Lg0+mN2
RDfx4vdPn8TPQ5zRas6OmNGLCqz9VzQvUvqzbxnY8J8XB+k3ZPm1vwVKHMsvyHW8XbBJw1/TnxGN
hLv9bAaao/Jq5FaG0jXT46qEp3ChXDmDqZVSYGrH+STFN5TVcy3RPZaUfPMVzBZ/bA3NA26zw294
0oexNxvwVFsSesX7rHq9ShfYsX9Q0ZiFj+rm+HivxYiM916G2fkKE3UjtO+ka2ENTozbytxklvHk
BY2CaRUMOpcf2HlcF29DQF5va2qMtXT+dRyM5bxFQnj2pPEoTZP7xZfG5jWtJh8H6KRUqjRSIwmU
Jg5TMLEvb4n/RUip0RmbsAT9bLanIHGj3aohlvlfz2RAjYdSzuvYmejA/z9bz0+tVQ/0Bl22IFe3
ZOuAbpieRyFWS6DmKGlRD5dgS9UmFhLeYatH4we8/5rC1PV1V0YOMPRpNZuuwlz9GXENervGUiGT
xWvzesjMKrvmN3cjCu5dhBxAT3FY1Wl9MbZ38tDXSYqSdIJ8KYWV+QttfN+8E3Sg1GjykX/3Et9q
fgjuqKbM99/r3bn50yUWuRxMAVFsIV14qxqZQBtWCVxSfE3LKSTUx82ntK3mS1VeV/fuJQSo3Q+n
rPDniDQddIlLeet2YYmyqyKshUsdWmCcneTr6jPkTmdYF7OPqZxaFO8rxnT7SDaiMPFJrnr/RsDw
OuShpdSlU8pdquM2BgJEtIAlfz/6RMsRmt17wGoqYoVakKL8mOyrRe08+wxTgQVNJV38kmOg58jM
o9dH7zmmz5PIW7cPq12AIRUFmtdTg6oYgkezgPyCxxBjgUjGElOGDsTUT135rBcu/7wShIoU62wC
BuF+iBCKqdvAtbnB2zVn3LMwPGf1vlx8yLsCHfTRut3oPZ2LAn+Abqvwp8BuIypRFVvnNc4LSwkU
1L7IQlnh5BktO7wHRCnv2uiss/HxJPZKEDjJNUojXMhVEoTGsCxesQtMdHiTTPcZrrdb1yOb8r3f
oK6+dCVdg3ieiH0gKSJubLlIi9wUfiWUxQho5ooObLzQEczBl+Z96GZ62k8jQov97G0WjBER1j4G
c61zWdBRXOm4HvqldYYs42Rjj6Enbj3ZpslHiukm8aQEIB8fnvvFUquQPykRroxzvdch9SEH2qUs
v0NvY0MrywW7fYrT4B9BHOE5baN7lIiBPTvOlG8rc1lYkJyhknsGiocCL+bZkW2ZnDeYlg1OZJ1O
Yaz2nAfWqY0HLwZSaqd2qRfFZkjrgGjZ6eWdpz+aCQ6chk9JRJ/fT8K40ChVGrDnzph4HXiRAnym
Qv4fxGz8ERwIhEuuqhWVBJ2kuypAx2NnmmdoD8SEBo4hnPStxxS0EfzHgzjfTXPnN37/0eMwKeaz
bQhyOjIBU9FFfhC7wOny8B0RRkXiYjCVLlffKOovs4bKsdhu0I9hD6y0yvqxc5J6AACblyKc5zl/
tLWnzn2H8DX29kuK+0YuiHJgQZw8GRdxmqCV87uFpZVCeVbtaDcuL4dnSEue6rywHxYQwxTXHA/G
rayZtl+FvQWdDxiyuvA7nXPcN+9KHSLZE2pOKC6KOeBZUZfx9QGW2gVx1/M16leehY0d+emVp33F
OZW8Oe21/ZnLT5qCfYQ1paTTU51tvnepQrpvwBPs2ld/rvwnYv8MnHKuyXAcYpnwfFl46am2gUXQ
Yt66b+8GLIemwpSQSeF0CdQrJ7I5cfluqDf8ztJ5OGX9fwZq3UckCYvmH5CGz4x+hn8G5J9Ulv/X
Pvgybq5EinJe6vJTEZCeRB+7UmJTbU3yoTdwkE5btycJW78Vkgc2hfyz4TITiLfLWE7i+3PKlszk
KTJ5WsHDVGFpLNe6uZ2hEtjwLziE0nEOmXzmNo8OhSRbHLTcMecrzlmJ5JrtyxAXP7sVV56gYTAV
fxyKTkc54SB4HklwWh0kht5Yra59ew2EnvzT6h8lO0eSdz5WPJHzoO/bEMgY/GQtHHrYS3C4127n
aZrazWu3rZbWgPuEvodQoED7lWA9gbLv6sWTJcKJRm7fr/z7vpN80MQcuDuoP25Gmr4YlvxLGNf6
/smApBDQuYoX0bdsEYMEnDsgI0i2YbYxOiTZxD9PxH+J9gaZd/6ckPAzkOCzzZM2t9va/EavLggZ
opkqNn0hO+qqOnswcaPaNydLw9gv3oUsSOQ8OjqgtS38YhjIe4lehDli3o+KYHp85M40jR+dR4SI
Oqo+nfSJuLj+86wZb+kB5ODzP5rPHarijSqDhWzsf5IlKteixZ21ucPOXHHsYd6DQY5HoMi6NG9a
T5axq9VzvqggaOl9Z9DckoqmWjKDfozE0m9iLDCRfQauvxW4j68zQIJyAghvgUetK3vOp9xaTXRG
2mjmCaKMn8ZaQBfLXn/FZduKtfjeoBlp39ryUGNtbV5sTkdmXmRrEPy2FGU1m1FgQFXP4EJ+w9/l
w2g7Cbgb9EW7zlG8u2eK04AGLDWX04cGQSjeun44HiFRXG1u6JLULy7LvZUzTVWJjufjMghiqDAj
pRqpIfPMuQQx0v63iNCwf7kyDe6QA8cRQOPQOQNgzE+zpBu7hTNfXvFiq2imryrareQC6/TnOFkb
8JwpV8AeBc8lqyUCNe2Zxy2uPTGjS1d+dZOOdlf8oJaQB7ua1uGKBNMSflq38GnHEa0cXWAU97wp
q9H4F5npGM1Spx1M56dHM2YiUknaYWjJANCie3LSUQLufshOm7ePvBe3xAJAiSJoO6b2wPGPn6fI
sTiIcgXNE+mgoM9VQXNW205AqVXp6w1lN41rGLLPBchqtdNfIGXsPzEUC+myQ4MQBWavYn7gissW
l6FGmb4zH9BRqcfx8XxvSJ1UEejmckV+Bx6cs5SDUGQb518KtsXc3+v0J3+x9Bcc65gVOkfVEYao
jFN08G8tXCZXdZYo8OpmIy2RXmZeuNunA4slso/LAZLFtG4McP+v+zPQ214lZKcLEPE+ihV835Dj
YCyWtvaEAE68vAwGCdbFlVFIBseQc7U2chKV1Z+gaLgnIn27yGjnwcpURrFUI10UStqONYnPhKcn
IccEYRZmYDlonTe7FgT9xv/rAXtOhUWGT7vEp/e5HO2/T0C5AR1+ElbV62QCOscNkMoFQO2ThbCd
asfdTWcixxUV7vZDHeVqY1gkXx4RDbxIn2E7yst59LfqvoCw3Ms/g994f82WFsz7124P5xLWh3i8
2Ne11AxWU0ubg+cPC8W4XtAOl7L5HbspDiXhsT3cW7Qf9OZw/zqHxHEP7ICecN0QgrQr/gN+Iy+c
necNStFt5s4/6TpaxGhwTLOhkUQCY0QvtXDvWBzRYwQ/dTz33AAFDdsTwfuAz0Fy9iVekQSYU9Mf
T/tyySLAiftHMmBAcL42Pl325Bfy2mp3YrQn7/IBhhIm4+0xKdHJMDdPO/bLpQbm91tt0pzPeml/
1gcL3kwgyKXmf84MrwCEvOp+mcf/TFNuFOLDda0UMc6wYkkS2UVM0GAHsahB2oL/k+T8V0gp5MvQ
PLzHcVmTCxaHEvA8OJzHVGZiirUvds0e7GYJfLGphF66euDjCpV7tpEm/pAZDlVV6MvPRxVlEGPg
4q1iFq59+nj9XXYALv6FP7PkP0tF69AJwjdtiGtcxkJK/IkphZsgpsDqKV7SYIlUhuutPLhCWGsM
R+gRphLl9KsB2vUf7WWmeQNjto7UHOgvRRYPfzrOm8HJ1Uw99fqAAbH581LaDPriKtP8odlsqdSU
Tx1ppu9mx7us6Y1yOYsGFPZFbmVCoRkRxo3xTJ6SyzTCGcoOdUBXkAMRviwoPnXt9UG3SqwDV8dD
0RBGCGBh4YB7SRaoUvZfMYWJewbBfg7OFuKe/bTeH9JlsFdj+U8Stzy4puyw10vcApXnkoKky4Ey
2ow3sWHMXPgmqf2bYVKZmnDBqbWwKwsCLcZGaVqnXpH+k9t0jJonZcfP2/CMfle137EZy49EW7T6
SxU/E7RqnT1y4Wn702qv+DlxsHKUM8Bs/J99JG7wAqMeBwE80LLpYqX7FGAjw/fquLNd1W/IZO6y
TYVasA4Qi4VxmXMxuGDhmV5a5zRSGO+enicJ7/6SAARAo6UiMrefacUeax+9Xul7dp7Cvjxsh8zb
vYE6kVGbni2df7qPu0wuERc6eSC2MV1mspDxqd8whRYaacqhGUify/iFkw4D+Ol6CJKqMXodfCIW
a7an9myd48Vqwjs1LVMyYa9HXDObpMGcacPBptsv/QMs8d7ZUanzjcSjT3kln6x/BUUve2q0c9xg
CgKaNaHp8JUP1seHNrEiT/7PlBjjmMfk1ZhfhtlHUYmozO+NqGXlrYV10BOrDqegVSh4SG8M8nB7
JCje62tKUlgVQWOfH6z6k22YeqRl63N0m3sZkaf2Ck/ndMRpMogsWGbmCMUjHVvGc8ZSVh/JVxco
LT7qalFYMX4FMAVFno7reQPR6uh9ZKxVhJGfZjTYr1Cd6ja24UhyX/Kq2ePr7znk3/5ZtXjaf31H
W0/oe7I/3zUF8cuse6fcs8mrh3s2Kh74yCKhvulBbk01PaKYySJdjCk0EYgTmlhqEUeBXjV7x5/l
7JcEGTI4HPgExTHpXtocyPr/jrQ5NxU0LZZdFSXoXH3NsD1KhK8y72S7y846x2KfmN4T3yg2hlDu
LyLhHr2//Zv02QjFXXKAsF/x1m9l88jdHt6qGBEMS7XqDYf9+J82xvA9mKebseGSr8z3J1HGyG84
LJzkms6VPr577LZrhrNXuncxaAucgwuf7XOzZ4m14uZ0HYgx4vy5fKpVEiJiTMRVaivwkMpmnXAJ
XRc5c0jISG5Ei63oeVGBhyrPIj1uzWV2MUSwyGj7RYf2dh/vBM3zh+KmQGJqOOb9ogDC9WPMCbgw
t8MuOaOkqBrNHyIcZKlf7ewlFUcYXTokMjGbL5ICfXr105IAiRb3vHlSoQERD7FLG8ULhZtum5nV
ig9bVEJgUXjMGnuCfrRdjwm9p6ZMFn65rOF8FP4BR3p092YmVHWIN8qjiSVrrRMEayA5Fhpmhy0I
Qk43tvji7lEBNv88qxWvglHm8gzYYqFAFYDqL2CrGEo2Ml+tXN5oXx8GyGXZSYpUU2YEzBl4eTGw
w+axCuwGwEin6HmySXQiTbbjIMsh8APYcV2vqzgYkZDhByyJuxA8hQ7i3TnIIJPj7x/rfK2JS2qT
Qs//UDmowLvYm7RYDPCN00GyW2jAxlOvnYGgImeoykKB4DRGi4Z2k7YhtEhzCmY3pOg8NGqVyphr
5rwc45FvmlDts0yQonJfrRQaTD8Y/fdC63I2N/Oc0QVoA6P3d7cLHw63zt45awLZvr618wLrTKt+
AR5UJfmGucfxPCwajjVn4zk7Ll5T/ZU6ikqtt0RR20n3K4JIMVSFgzPALblQXq9+CwN/neYkEpFK
jUi/s9n2yJxfGSmJuqV4zGUFHqdA+JJgQYp9cK504+Ek6wa1OyFH/TQkq7uTnNQUMXoOdzgHEOB4
GyzD2J9nKBOWnGLtTZpNSldXjRHTdRY0yQMyRZlsnQWppmCsqlQjn/K6HH/tapC6QdXXQcZwWfBq
HurwkIulP1NNvkkgzqkoRPOo5bkiCmDak+Fm8xLZemCWXO5Cjyro58U/lGHH9HTmqRPr8KoXp17+
xY2KPS99+tBqW9ISr2xgrdqf9NoaolbPLEMj6MhgibbnxwDFb+yPyNXJUkp/dP8OTxXgL6rDFb4G
38Ww3bgm1kmh98NK6UvW8SzcAeUcMNzZCXQAXB6pdNY4pjH9mMFbq9SZaCZQAt9DyNq58TFLPAdb
LpmqqYtxl1WJeK5tNqwNydJmt6PMqVy3Ey/HTMPxmmEWs6bXrkZwwkvse87RlxC0PnTCf7qe5eyo
5I08YbCm7C3FHcrz9PVNOZP/k410GwQsqmsOb9lHqxb7f0dcfH5XZw0MGswiU0UoH5+A0wJP7cy7
b8Dzbs7Ij/fKQhZN8vlGgLAWmHf3+740MXOXfvOlsPtIjVXQFceEPgUft/2NWVUSfMFLhYH2sId6
UknkMJM9eYDaZKSkOEUDSRoAtDWXeZyclVrU/bLJLAYH5LfB8R0Lx7Zb+ZEtpvR6FIiGcXp+9INj
Vt0ve0wM231vvufrZ0II1OuzUCrJqbovLNkLhFY3MBv6ZPAY4qPwT7gzV1qLp6k9eT48mIv6CHYG
lvcgb1dVX1x3SfHP9Gqel018rv8FwjBj0L2SXhKb/J/vZJT/XmucKluwDIx33Oc58v49k6shUVKr
sIzPbKgCS/xSlMJpEUOi62JW5flxB+9d9mSDJSN1R0mc+21si4b17fy8dBgtfaZbWjdptHz5AUma
gHEHpOSizg+YB+GT1hmFOSc65jOdzicp3eSG5cpCip/FozZ2oRoD+UZlsn9jnl2GdND05xJzTVpJ
QTZt6ze66TiNRfpByksE7o0mgWfDYbBoM5Y6WWbRO5Lphh0w60qHoGVgCod2x9iCnWL/YCBh2zAo
N1boiQ8BK2tDJDZ2arfgOrLuZbBZQAjhouVAECqMn3pxPx/lt3Mtu4ClXq79i91tQ0Xo7T6ed65d
jmLVq/lHZGioZbi29Uwz6FU2Y9bGPT7gr7ffiBkM4gFIT3GbLH3tLaVXTc0J0v626arrelkLYnnc
ROL1NKQds1s451WtAhue+9az3KItLN9q7G+d/kULhgCDxpf7RJH/qUbWf8N9c9BU3LtUK4+qF8+7
6Lvygx8Fexjy0UYAnRMDCO3yDuTDAzhtu16DxXENO9hPvjZmHTkZ/O/Y1l7aV1DoNhr51FPB/EFg
U9aaUcrRRuResxXuaJBAJ0uG64F5CswhxDTnTnatlbBN/36MyoNy80LDhQWTMiHO7knCmzZwvjcw
utkgMfT58JZ6fLCb7MRqVq6YyZpsO0KLCT4zkXzYBOHkB/retMn3fuFxHAay+ForjnI/3zH+M7uK
EbWbKBp3zwg97+s5F1q7syH98OGkLt8E6pP74YVMykUh2yLaRs2iYGhi0KYLbjx7AZLNpgHCW39g
q4JVvz3l9jSRtFRKeAAW4oHMcoIWKai0frOuX43LQzsl9gRr756oE+aGTEu5IoZK+cfNSx4RhHgt
hFm80C4OEDy1pAtGqRRDidB+E88yHO4aoBOAeEhW2dYteJhuVV89swtncWeGh6wrD18dGpd5SHpc
/bd4B/D/TZiWO6CmwmiIgUcmtKVWWluOs4E2VFFjT8LqRysjw4ib1KoDEpDUUyZ9NPUr1vTdrKrP
EpFTdJ8YTIpZ13LIyllb+ReV/KuEUAkSrtkZ5/g034oD6aCBBCE9GK8ZxBxZQHWPx0AB+IEcgUtN
58ov8WMoo1qKfG3ZVgMLNS9RLhhziinuTwdMv6bHDxrjXWucsrO91qNErT4fKw/G4k/plEODa7ni
rC9HFOy4Z0EbPoFahZ1MO6qZ1VunU/uiBvVZxEZitJzMlp+CNNHIXrjlygscbBl4D8zDlfm0ONUq
S4b/1b+0yQt2a5NCxxRDBMNTI3n6JxgLW0CFQrEtm5rbaCcfddg3D3NJvYLWGYGXv2yjqFyrCpPT
ahfCrfP0gwh98hnxDkqxkuTm79ufj1GipXcaayuFOOYBKOcwVYwH9npojPowNZ9SwFbPEITlQ+R7
KTsl0VWY+qEUiPynt22pzv+5vCWoBTKlohk9rpa+A9rQJZiicHDSa0gg3E+3CuBYpJ+ppP8Tzeg6
YXuV8cqc5tFKKC3CyPc7pYuyYHBEz7eSQzCdbzatpLkTLPDg1kAk/w/liNNu+ojhzUk3A8mviKQe
vll1jsgsGKPGd+up3o0Oe/eII7DEhoJzFV3zDy9HZHqn1SXMRedvFhxW3Bj1eak0eSz6mjWbLhNb
4Tdp7cTUf0rFGJZgyd7hTxpZIYvySr/omiG05tQXCzKUEUuLaWrkRhQIqAhstll+cGpmN/qshBWz
vKzt+u5WrfedWd6M66u0hC0kEGYS9tF0R4/styvsLLZim0uqr3eQZyNZe0VtUV6aVu/agtXUV1U7
Eul4qIzb3mh5fZOaFdE9FD05sbMs3H29rmxGw5ZHJaqabnsoawKie7dQ0IbDtB6Pduaqb6ZTFf81
GmmNXOG5SaUgdkTQnn1W1qMqS7tLtLkfcZYmPxH7neQN++g1IZIgFL8n7Yyumhs2XGq97CuByNtB
EuAJVrjVKTqgT7Lz+JbUEeSBFpMxHGxv0VUzgGpZdHO8SJJaFIPnrTPcOlyhvwQj+X2fFOESAkYm
mBW1DYBAvuHa22ythDZWBvkNhjN0uD1SFjrDunDQKSxQeU79CbRZnVO9IqB0gvy3gh1D8M5uCkY5
wlXQkEa1jWskbVluYlqyw5Sc5YGLDodkgQptEf5Hy9wtZRbYYAa2awLUPW3lkpre/kykSEL5hEs2
QWjhG0+APKQInA6l3yV5xHU3wsHSJQdEMF1Sjv/w4d6aiHapZXb90+l2kCvGtfWw1FyY+ycHMGEg
cztl5RqinIfZwkGdhyw5zXerqkV/75GNulQuSvvtS3OMc4qgYUxRqHZLshXphuAoZXDTmRMKx+WF
Bu1sEJN4h4YUFqcvPUJdU6RXfd88oq5vIHLE4iczvFMtJvHi4gT7xnKNpEmlAUhxi/1iugnBu/OE
k9p7WWsPsy2ZQ2+bkU16skY1rg09Z+qPXKWBYhqnmL5zq34o/ZOO2IMrsYEjqiLF0NejmDDBdLAz
3EBNychjJ3nqjDPOROYhfRO1a5V209BlAFxWirhclpoEArJYMNTWJ6RIERO7VVW+znPBo9WyVVD4
keTF98UtGv6Lm6W73Ns3Ais/RlSZV0eqCIi+yVbqAafo2dF06carn537BskSLZ78omv02md1UIUG
DXD4hrFzz47TfeNQzK/ZJxQNoh1dV5KQ3MSb97HWroVhmDg7Q/0ToCNdMHW26iK//5of5VcCq/pd
Kd/6WQVsD5MapWmCo3Fg1pzIBoRfIUrYHJICwBWlOl1UPr6zWdFPg3AjIScWmEVDOg2UP0+lwzSu
pLAWgXrwHd6/nYVPy8bjLVp7cIEeGnAeT2dVj41mSQJ6zLTf3bK8Rj/V/9GpDo0YJbCaXmEFhs4k
zbKNCAlRnpPbLchF3ryFgiJuWw0ryB1+92VZglH3zklZsjQFwWvlzL/RDh60sNBihjgX/k6LlAfa
F+NeS75FO7+nZa/MPVpKAxZ5+F5xaznnWjNo3+YP47XQVMcH9EgJm10sjzFp5l3jbXkDGGF1rB2f
xUSW/Gjp8UuPqBOijMqkI0Z/TgXH7OM4a1NKkubseiTOOYsmrzPCtpFt0yHU73aTt+ABo7iBwH0/
zwH3VwY0K5Ybi7of6hbrbneUdkN3j+GH7G/r29b8cAAGNTYTHIPDbttwup1jh53xSWYstueE7WE7
G47AUbOaM3vrGsO5m+A9nw52iCeX8Wtqrl4KunBe52d4VYOarAd3uM977SDgaoQjItPZ9CKBPcDS
wCFojoEolrITM9CN3TU0QowZi6uA5bt0jGpXWcUxO8IFOG27ZaVmLcRD56bJ1RuXHwBleFq8gIjA
g9pmmMXWioKOVGe/Nhv0rKmToEDBAmB0VhEwEnf4uK+XJ9WGWclMFgLWAXhsfmRUkvxFTXnB9bqM
nUn4LpQypJJ+RLVX8EuYcGz8GJKjmaLGYB9f/cgZebhaGcpLesd+eggBts8ub9O5YORh1hriyBkV
tQHoI6Zo09TDd6p24c/CiSNnfps4uIHrsHFYdNeqOdojFBE6mfggMfaQuXAM+vyf1h0dR332dHL1
5t+Hnm/t9sscEXxnmGyea0pBm+049bMvUS0yqgfP3BGqJSqDRfmwlc8JLJCl9NxUNhibIYu5ZXP6
HRwM+Zm4T+KjxUD43a55SpiDZwadjQsnsB253XshDFSrdxDNLdm/Lc8uvgvd3IVGFNT+uXbKzKhp
5GiQomz6Z2s84z3K84Q2th1DmYYpNwr1zgIua9dzijNPANZuShmnuZj6ckn4+r485KV3ZOYNK9AS
byvfjJMw8jsIfwmwBJD16Hc+MKKAMhAMdoZGmrGJNkxIobM4lrBjdPwAy1Y9v+qYdw5aLh7Krq+Y
AZyLS7bNN7hx+yfYTtb7dAWmSkrLuwdU0MwKXVk4nG1vSHFXObYEAVcie/tpcZLG+XKWixfLwBFi
mkuN8ETc03qCmifnxT957rDGIOSAqNTEkdgsFNJmf0F5h4dxo+xEUB7Ik5Zu74jWJW9vsd2Tbype
hPcy2NM6M4T06s33LOMDie972yAOT2zGgoukVNgX5ljPqjLEgjk7XTtcxWbWx0FkLRDxt22+W52X
q/Mqw8fmn7Q5a0aZuSxIHQRMsU5h33RWZqY8HERv72YOKXR/t3aWNC2tZ5Ts7XoSDapWuvwVjMVg
GF6rvFIrsAeIz7Wr8ep6cGDG08YJZIVJd3ndMn2zJcDXY10UOCzH/He+Azp1ygvw4vgxCFOZS9zI
y1F4MAyKto9/HDHgRsT7mF4jCt3Bc99pjo8dnJb0XxRq9+XJGepaHCRG4p1tMIv891urXEXsnjm0
9nEnq6VRXc6ffjBgQGAiQVPzCD2CIbnX+TXNCxI9Q2zqR3LC95oMwC69D2DS7CTZH19+lCv1hUMK
0M6SPE/+ueizS3VUvwLCllhM7UTByK17cthwsOT6Y1CLwe3iHy/kR9PBzU0U2CD2jJnulTZLgO7n
EhLHeeZoC7QNH0FkDwqKS3C73qaSqWbHyEtX1dn3GAVm9aMcNfiujM36ZZfTJ7cgEOVy3fKaS9aM
3EayQC3Z2ULsIz1e8DmUGNHO2dlvZhrwoIU9zFzJEESiWJxIyPitcpsjYmVxKl0FFmJ9Z/vSa/Xa
a1cRjgTqws177ZiHe90OkbqfUgv26csYS/KhdTHuCIzgOHaEm7coIXI7+rgIvsd8vIvDwI8CZjE2
7pCsoUY5D2PfKHDubj+UE2JfJz9RcuXlVAgXF2C1w+7zDMC3jOsX7nI5Tcz6NanzIvwVYhmo6FFc
VJziwVzv4kBp7ShicUoWDzLkZQ9KdPmQOe7sj3ksGsf9MSZehkUy5rW87eRmptin1Oi2i5IfYoq1
tletvjT9uu4G/pZGrxlOvKFTklEgnNewvF/Z1CmcB7TDFvOJOhG9CSxxQ3Z/fIEH4BhjgJdRYVEg
jv0slDBOi9V8fpep4cpTXeGjqP0VwDrGOb0tcfZ/GUb7lawndmswpISfKQWwd1EJ4mTR1oXlcs52
KpJXx+h+Z56plluPSNAm6nwFPIxN75ECUPb5VzRDtD0Nvk38oSpS/zVLfupfcAmp4OuOrNiLrTBz
GfCkUta5MlTDCl7OIC2ZqZD043dKb02ePVl/WVIhDphBgIlWQ5AREBNoHz0ILCx+6+cjtsHbhmZO
08C9YLR8oCAnh3YKqsTsKmAE1m9iSD3Fm7iDuEnnmIlC2pCP8oyWafVKz6FXfVhNcs6tUdPbXOFq
5uDU1sMvQYP3In1dUlj954ZjAPjLrE/eYloua1pWosxQwcA8dLrNWrrd1YZbVenFbRnFIgnFcn7L
QgtqDXDEE03QnledP/X1j27w5At4X1OhREfE4CoY0S05cufazmWkGdC7v7ImOo7h/RW00Qecj/Rp
hwE8F0RMA2zcdSI41kwUvFZo+7iAXSJBKliV8qPkY8HgkJjwcBqsjT60B/AMO49Mp0DH+Qfwvun0
9MzP1C6TPZSTVdwU6b5xhg7uWcUUTztitJsfrHVZpwEIqN+nW9mpmNIDopovboZ5kAKDuUEkzNMz
6fkEXp/vAAL1dYpBQl00WJI6PTiKODTJQPmMR7x7gdkWv4OBhGUdNb3PFJjjSZlxvu/3KMusdpHM
N+guTz9+I9tqa3rKWNoC2xPZatCrYGy3/08rWaOajUM7o7io8sYmgbd5Sq5pDAjzxxI6dwZaBACD
4CHjb41BUgKgawpvXLAD3MHcbyR9yN7vFSz8wsKNWeX+FGj00piIXIiOeTrGPQ4y0z+PF2tko0mr
FPg7M80/8BNJQ/cTwGSwPk9jUSVrrgDf51xqHeroua9z9xsnAbMRk6Er75FfhFx1i1HxEkvIfmq2
sdE1mpDuDELgHsW0iZjNZ2pm6dAvzr+Bgeow306FJdQnDjlhcfyTWaSigTEuCF81PoZVwd7a+8hW
IUFNTG5IXCO2FXD90lCjM5gtGxg//JcuIeVxKAgWIp4iYm8ShfGjtypD/GrFwftJzNcj1o1Hc+Wg
1Al6RVmRLbtg2LBZ6fux3DQ66i3EX5LkrcJJdRpBgTgHGj/WK3gTrN/1GRxeeZP+FwK58J2V9Ffl
YQPgp/PBwyZ9+Westr8Nb0A4wfqb17Hqq1glNG8x6v6H/O09H9C88aYVqS5Y3mTma9vD1+RkH38S
lp+EeWxvfGsICzjMiyx9O90F/Y+JO+6z2xCMAZ6l0i96b+uwLutbmRwo6Q1xbJ2yajQq/mE0g58Q
+9FS+k5lE3xVoNXBW8rmixTwaIqip8QzWZxgpmms9X9qrckkBGl0+1gi2JnA3eBOSUKvRywWtnlY
zj4j9NZjJ2M00ZW+F7UH2FcizmYR7iYzYLBcy32bvrvKDoM0NQoIqwyT3Y1QzptG3IsxT+nae1tU
/eqak0bCU4dzpNEBeZiMuIaSKcTbsjwi5W4yAYPGIq/ASTpIHTis4w+92dMmCzW9Ik6ypcXcNupr
KN4I6VYAaXUIhPXimFUzXAwqIUggyjC19kufsX6bEd+xiBNcd+uQXqqYgUffmVZUByqP8CotuTCd
jfTaogTHaoTQz9H0WOF3HNDsk2Tr6/WrpNDfF1B0hzNjruwnFBMTW7lfWqmoQIepA1krxBvX+0vz
NEOOMrwlbcxmaf7vkboHHK93JKt6MHoo59dENOj8Pk2LjL9vu0TLxtDmmJkzfAzSIHPBcmzD1S6a
vzypA7w+tbY8no1o8rdZPFdEsJSZWwjoaGbRNa/BirP37I6OBz+hZlksqsVCsrcx1Tbw3cs3UdVH
hzqvugsf5nIoPb7RmRJHk8at+nBgeHAZCM3ZLbnevZIXuD2nDPxi4dkDvdG4DKh7pgvSCsM5PJtf
G/4oMaOIipjGcjOzlyGaksdK5DoeWN/L0lCO8ZnqPhX2+OGDtb997D8+bNws1xpRGBQ7gb391Tbs
OUQbbxhpGYsVhsWdcljD1gPAvNUZHLQEyqSsQ8vYrNIySWrlgvwDOPrBUpZp3viehXesjf8u1piZ
LLHUTe51E2reXEM9mMC+QFrWZ9g7ffSAwmS6dJkdIfJEV6H9cerqlETpFfBPn+ansmxrmLNzFPTc
D/Ak1xvvRJCiXQx0rs4MAx03I3ZlKa/Bi1YmoHTJL5LPhahHb+35YyEHm6OIndaHGrm/2paaTuvK
iEFW2H25ATRTgzVxz4VoLGh27s2OYDkkSXv9Njys9me8wRhEo9v04eLdphlDQMbBeTzgtzv0sjam
vla778CdLojbI3iUA1UvdYqXsOa0Y3MVF50abMFVlSBoo0fPX2paMBt2zGZGAPIpOe8j19z7CMpp
Ot5DuvLkmQnsgTPnqLeXA9Ukps6AOHVoLic7Q+GFjMCBsU+qT9ECvddFXUmIycDtZz2/MWa4TFO4
Y9Dc/c4+8pcMjTicL0QQHJzbLi7+A1Laf3UzCELCyFiubSyWvhs5h+qmieFqYyq7JHLrH83qP+GT
M/b+vovn9tvdfT0mN2egLn+dgwsJ+3d6qdLSK+7wpKLvwy24EOQ9CKcTlft76d2yKsyYAihMtHyo
Sb4hbgqHREM3SNP8uTqwJxPSuchFlucQF/y4104q5Fa3+4NLB/8w6PWz4SbUC8JBujR2ExPMjnaB
A1oQoLG1x+8YlgeTd9ehoajm/7GgqIqbFW+R5rewRj9sWgneo6FfcOlj5BAjPUHriRUUH6JgJPOw
GMNsY9hqnPrWZ1oCSJFBgMnYFVIbAVJV9GVohqUPiUh/PFJWk0ZNQ8tbwbcAtLu217uJK5vB2n+o
ylhtEqT3kQ+JFyRPMRgiCArlM0lSV4+FSxd2iC+aK7TGCH0j5Swf5OxPSeDhokoNc9u+8S2AWp3h
Oivkee0s4TV/CmYYP/C5E8ahbzNNsMb1fRItF90i29KBY9NYH/4iu/wfLit6hBWXd8pBOMYWNDQn
bpBXSlUWLrfsPEuzHXAOXhjlFzcHTquHaZoTKuyA1hYmRW7KgpGe3TqIR14uPmMct9Mab/YJVrYv
vuCDWb5PC1HIntyww+7J8XXjUL1BA6eS3lVCt1kIgPXBQ9V+6XOUuRG9bKsmv1er/xlUgGTB189w
msowNiLpYflAoiP6zIusl9KMF6/klwK2pxmibgM1sJAAgN+CcaQtoK3Y2xOoHS9vvGGZszm+8n5/
rDZpOnyMIuwirNP35w56oO34LBS0vZky0oaoHvPYkn+ODv4ecjDFahUab592A5pnl3JTKidKyiuc
FYgyXtxTXoS0V1IQ20XjyH5FaOqh4+jMaYv2EOqip28zf/VusskyQAgBxCw6/SLA0uQRkQnuY6oR
/4j+In3fYYqfT0nN7fMmOpaxKunHAFj+wJSH6vfhPEc+zobxTkzXhW2sE/JoBZ/c6vc6DN0f00+G
Gz4fLi6wgwmHiOUyaVI4BGL35Vw/86s0BiKmbtj4tmFTOyylTsEe0M7eQVkY3tE2Q2ULft+Zx027
ACm5tCyaz+c8T/D8+PEV2yYnkUEiu0SjlLIA0RteNjUxyQIrsS5AYF7XlDb9qkgv1wqvxqfzKSKC
aokTonAI7FdjHGgqDJms31EzSZiRHwvwfB+2+IndQD3WF/4jR4Gu5YNakGrVscVDvR6ztiTCN5eY
dKCA05R0zusl/QJZH9Z0xGvFA3G0IC1z3242VeT415T0RVMx90QnTj1N/DgPzJqgYSeENezs/Vig
PYOsN81kWSAjeoenmBTGavQ0bEEHO/iV7Y3/jcfukBrgbjQVsLS1kuKy9Ck01lbI7fcSFkiwPFN0
Huxbg6masqLwDwgxU1EgBwXmrmKQ7Q+2I04C8ZI9Tfot0ZseYghFmHNuiMynapq/n0ZJVG35jApP
Jn0gT5riWV0QncP+tT8HsYQfJ+LDUCeKLG2Y8rmd0KfU/DREr9iV4sr2yr5gJ+fyMx8lXJmqWVCA
Ianxtb+yv4eYl6ZdX0G4A05dGK/amwuDaxo8ElujPOvFn21PEX4ju3zXLOJk+8oeV1h63Nl/wEQx
CkP1kHWRh5IoTSCxgz30GXTrPXkY7N2ytWA4A+nCjLC99Yc0ME77pd5Yx611r2kz9rDpjIDKWJsO
FVlIDxkQXEOYgVFlVIf0rFpLlOYeEmcoMOEb+le6YPcndodOd9ItTyHEdrRnXxQbwQJQ7gkng6Ie
HV3lSf2U/N8+W/6PLgFK0fSUYaAmxMMLoDVl6OZgffxEpEj5SQ7ipZMK+0WPWKRne6Hv1b09K81R
5+AL0ntY3oE+r9I74OrKSzxOVI/4c/+XLKYYrqD/hVVGZNlcvX5XDvmio7HSO/9feGQwPM21jAm6
j13DnLo2ydFICXzDYJK4MgAcdvtczznSiHEuf6zUsEkCplh03H8vRQX3pIEUGWsSFKdmEVLO2QKu
GdQJa7mF8I5kvpNjdhp43dNhxijF7OiVSZbScu+pz3kiFN3xlY2c94yOX8JBXmXaeZQA/D8UiE3U
Bq/s78Gy96XDqOeiiwgmS+QtNnfhXqJPE1G6h1ta60QIjIonvjtlDrDd3+sn5bX9aoxTb9zfZEB1
nUOixx6hKzrUtj5JAohKilVEMY1uD//9CFNizAJbdn5rF5xUHkPmeAbc36WRiPA2PPLT5LH6yQol
t45W4YKfcJiwNPc074HkIFDz8EQha6jWNpH5Vujb3z0OVounOanEsgq1gTqCj0mURvBhnqCqwQ9S
7E1lO4r/4m+W9CTLGYm1Te3srwl2Hsg0bPuQ/OZRhPc335RUIuWxPwmvInMM2Ub2+sSdpg2T9h7u
65jkAbmiBV/dDF8q6Ml9mBqZGUwMpD54xkq3qhiVZXp/J8Ss8WwQcmfYHQ0mIdQC4PZ79tvcZKHl
oaGnV393Eck7A56/a5rV5FLO368n/dVyIh6wUc8FMmMo2NNPdIBHBqT3svQ7g6NPcT5jWqDzUROS
ePkFngpPxpIsmnCTPNP5AJPAsOyl6t2wxvwbArKJZswThYGjPEQ78FBZXmlFnRuxReAJmzjJ3YIc
KK68ZxK3sRskNv+CEldrx90lGzjDT+r01JPcAYqIc4f51LHrqlocM4p2TRNUDRiNhFm4/8ljKFKa
67dPy5HiZy1wT7l1fMaI3rtykPriL9l7SiTFB+Qhma1sHXB8Rr5sId1ETIdgzKinbPjaZsyBfiAH
Qj24AukdZt8ZjM0oj0ZdmostmjMrev1zRUL3zT7FZ3gHZkIyvXOEeA9AYgGvqdP78Wxy15fpfRsj
UZ734K8oePaCtsP11OnIQat6vzk9crdISQD442Si5ICCBwZM+xPTGcv6hJZCd4WXvNzXSKObgvkV
FXdjuAqSG+Y4BpwkzA5w2Un1qx/T10Yq1YGF6JRe2DFbMt0KM0q6fDhOqJh0ugFC0U4v6m2KuBZS
oofyqEO0ywGIrKLud6DntR/c2CUpH0EhGJVVao6VzMdL1ZUf/yUB5RXuAMNYFGDnGbRJxHKxvKsM
wZ+Of2wdb0Ohws/AFpbMnxrA/erkFNiyf9xGWprK5BpF+JZdLVK6xcOhEbZs34zOwpo0fQUEO9Q3
WfGyITFtjXCJaI2iUrsqO/qPFK3Dgd8DbZa128YKvGiug0y9zZSy9JzWl9BlYDJ5D5308UdVO71U
kEJ6/SsLpMkltIsWnXVHZYgZLBDltjhcSdsTBH3doFPVkb+pLO7gKmhY9QlR4QOEseTGisWZyZsY
REKY3q4mF/aB+XSEosV2yp636VYkTvqHAUUVgPKoWtE+0Wm4dNXZyz52k2c6K8b2adtafOw/pufo
rJoPSWAtPaUjoKO1aI6Sw9CLeaqb/zm0hK82TtR94xTUjx9LbyXClnr7Jh5R54NVu9zqeb2iElg0
yuFsbxgm4CWgHWZ1Y2w91Z2VO/tXy4Ga7SpxGuNuEeSHVdQGV9tlrTFve3RuVXGVE6lfBp7qzqLa
GDiDvu3slnTQ8Ma18TEUoXqHatsxDPdZyHANeZ6jDpRIYx3zAUzUyk8A1AQxCkwWUG8SxomwEMLn
QZgtXfMFpnaVtFNyfDf3Tamj4Wahp0EES3bDO3x/lKEQAmpR2tJRpmtznZdEPJT6FVf3Bgd4k/bB
t8alvc5c+da8r85uO/JPCWu3C9XRqRzwuMTxLp24eqPWso19yOEjHzpucy9XGMpG9+YnbyNeOcDC
pLXp+tgodKW8jpLlghELxLRh7AHnd3PxqKj4ZuAiSq0PnzPavXrgigkJL0VO1YtLhSHQTRdl/TXa
xzRtd8cVijgGj0J6IVa0VLS3ev4RLibPvFwxR32lX5zWgDAxtqfeV013iLbi1v+7YbgVusVrjN3/
lLr4z+qHIn1/9pHQVxU3YJOFhx0cJk4L/4aoUgCEZx7oxTirL09PNvz2vHlL/AiSQuaRMjq5NN82
YEqpa3zFRubhqGrr7Me9LZfKCf4J+C5cnBf0sw4k5urfhv4HN6irC7DDwL9xyR+g1rS3JMQEJR4Y
tfp01f9+ySM9g+mlG+YqbDKLIX4DzU6OuShBiqrftDhGwf4Ax/rKHKKDhr9wq7YMg8w5sqZiPsKm
ip8aU3GtP93pp6TpMUhw4r7VvZxO+jEispLm6F9Ei4z4HpTRyxT1Zom2jMpXykkRfTZrJn7Yl+ZL
RGAZ2rAZT9EZc+8h8a8GzHUwigxAZmbtWZYQWOJw7l8gg8xrZrDTYSE97eIoTqdw1WH3Fmhaujxe
/0JV76Yj3sDD0ERBwGOqUt2ZwABwwi5nngMmkYvckVWz83z88rAYuLIx5AdYVN8evY35Kdjy5Bql
5YYadu8aY7FEXXZg7ujPSeF8RjNx8wY80mpfylwL7t0L8t4TGSBh6YpWlTJZKQ9R47yyJU4WmDzv
iqtDk9uotU8qlz4vI84nZN22iWUS9PiK110n3xltmx0Imu0laqvWjsNyiwirr6u9d+TsyJJU7xTs
rS+5l+PlctzvI8DARLEzSXwuE0LueImooB0ayXu8YX2pDy72eZaDycymFk2di8pv3n+6oApb0bt7
D+523H15ezyGPf8iS5uf0IevHZUfFlYENC1dUgWzx4K5oq1VBcZi3ObTsBTrLT/PiigOMVupaaDT
GAtzDEu1mix8bISX7aI5rLaJnDZGgmus5JyVwibiDwuI1iCFfOmPcCy3HTPmpDaeYU/iz8ej6JYg
b2k5ZfymIq5izG5U40SH7hd9QzUR1OY6gvykCpUAJXMlLg8ose4ZmjB7d3E0uaVoK7cgm2Y+sjRQ
NDEAwQHS1fI7t3gv6B9j/FdpXI+z/YOjJAKr2Tf3JesEHgHFuCahMxSSkLvY6+ngUEgEQJ417e/U
txb4TxIO8PgPwQDj7I8/MJCC+Mu4LHN92DIwCiIUMS1ZFFdQSSOiw2alMIYwwKCTsoxxy60+IjD9
iy3cL9lbCWQrFj/83rzZT9kREM0lSGwh4fLn2RxNzmheLGct7wHglI0q8qwkT0g+uRH/JWi55nde
hON328YTe1meO/1iNkEBvFAvVdgH32so3DCmPRUCWDUGIpK6Yd1DqGOoCAN9aVmll98YggD3qwUW
wMdEuQevRO+b1i+lNbUNkYXL3h3RdbwzMvMtrYdK/O1tDRMBRp1iVDeP0GruULRnS0IfKO4gVGDr
18grFFnQpdgGUXE7iUwYoqotGnIn3tE/Ms9KMfec+cZRFsYzuiaSPkc3IsEBBXptuAQ2JEp/zyJB
4uZWO4jR+0+p7VCnGnUhHFNyPsCdsBtDYa2cv9Lu91nBzuQmpfDPB6/z2yozb+AzE/zmXs5tuCyp
DU1qYFtL0LEBo6V6rk0TMjJoOr5uKMJfb0ngVbd/SzGJxyAV3/7IeZPXFkvRjK64ukNMPnCh6Xyw
QTRjgTVS/KhrySCK+9mhpEukV3lVBuZtMrr6z/jIPcljjbR35XKRRBJYrkGA51oIBI2e47H8XCm5
Uw5DmUepWfuhMaZ2nhzkJYzwNT0rcSlkkTEI9TRetomjC/zg94ScZtHVLUsEDxOWnuUFgT7mEQjr
qf0GJlgBNevjSpxCSkrFR0oiLY3l5GaULxYhxAkK2qBbczGCaPigrLud5WG3FoRGuc6ZJbezBRPI
IloUFYpzw0P54dH81mcaao3P45cOMqxNFb1rrJOBtCduSN4lkHsN0ScTdo5N0R4XEqvYqXpn5z7A
VINW681+tkbiBagj0kJnZCzmbsRxSjPKCDW+TisBaYnPYMoooMPoqPFKN8vsjFNb1JrCp56jiJsk
iRav8wk7IJh+9Zi5xMZqgPpuMkgsZu0FuiWjv0GBASy+WFUEq3upvtTdBuyu60qe0zskfk11IpkD
JbWOED2BIYcizjCg/bmSnjOo7hRGEhpeW4wnW2IukJ4DqAa/hTNk+3nPEBKDMR/XukjID51a9ekZ
8cYSaiRr05WqqhHMJmaZbVygK2gwgwM5X5VtLp6NN1XR67Depiv8SNBZF/GbAh6EfN2keNmmJeaP
/UbYwdjOA5eJ+h//7ar2+uvSaWc6s5P/xnVLQLyfSLI582i9ccl3lFCxBQIkuvj2SmsJVhYgz4CH
5VZWKbeGJM406zbYkLp2VQPHViyeuQEBsc7gDfMSY8JrWVhUjNF6dmqliewz0dDFvwtSneBC11uq
8/yBd6Mr7viAMDIzy+oqSRdWaFjnMnXjes456eFh1tou3cHnueHjTp/q24YkwDjkouiwUO+BeR3W
rG7rNrG0Q9T8RFcu9hKlcjkqfdWabXWHjw+cBlO84d893sPIye41tACc8+0VK5ItsDQsT5X+ddgx
MMc8FIlyyJzgRWLXhYs20mB/0ZYI4DqLoqZNiE51Fvor1xQFVWqewIyb6R9oE+4P0xGEFF8Do5oa
YJiDzrbklDer7ryTaEic+EO84LXhCcnSzNEnqrb6gJDvGJyaK2AhlV+IX2B90aVqZIWounulCOrP
6oUYVmVG/Ul6d5HRWIwKcL0zSfDe201r5GIYHQCtpfWH8b7erR2ROQ+f6PJAL2nlvcWLFCnTrU3M
N/GidUB//jvPGzKIVtdS1ZVQYRk/W0OFGZfNrcWwvdXsKx27Rx9dMG8A2DgdiZ+Z5DhY8twEJGxw
qk6N0OJkPiw/X/ZRH3NZ3da2xRV8NOaVwcZSmYKIjvJiDyXrs3hweNOIDOnlAWtx6dXC8hn140ab
zNYahgb5slRdLz8JoclN3s4kXgpdOezDdBsyVvCP6kWHkNca8+yR134l86zaLEgEpnI3jGOvFgF2
cNG5YQWO8JAoYmwVRKheKMxDV+a8z7QP3skG7DXpHw4cTX5ASHKzGgi0kkwKEisYZq54tCAARdcg
gbUtGN6FtC2JQhcPcd03J+9z5rLBsfrvTrHmK87Jfw9JXwWjwXFdiZPUTsZYq+LwlbjeZMTStW2N
CyhMn7jQinGnIFkeRF3lEWaN8AzxT9PCY064pjjZuc44NSUIuMfqFacgnq+YYv7LUBwolWRsda4a
cDXJTZQFtRSDzrRuGeYoponcM/4umCc7gohWY7tkdATE5CfC5SQawxMpLAFNjR7mPgAFvxGdmwGy
WnT1ulhvIpJN5B3SCFF7RaVF9MVOBoqQPYPpiEKZgGfz4/+PN69o/wAjTMahb6Wn2kH5RU/D+EWo
oNjDKf7fRchIa1KKJwV5wAwnpIMOCgB81DfpGM5FvUUPz4eAr//19Ym8PVS5p71qQbDbHVNamwRQ
KIf+Oa2HulWkwlG4rQ4frDu22g5gtKXQKPCaGGEbws2OSFglgvG3oNnxF6EGgLFr5+4kQQ02S94N
9paIrIy/IcGTnZt+ZqjYL5dpuKGw6tPmqkWKwKqoqGFBuF/fZW0CAgo9is2cFljCVaRTXnv1KQsZ
J9YFBtmH+xbj7DPNgtU5TpVF26i74xdUneZ40bqu+gzmo0SU0FXGLl9NR5bI6u9HgMVRhflafno9
ttZIV+UpSBdj522SYm164/BXItMrUYY8Fvm1ri65+Fd/aT7f9TELprTeKWvl+YqPfBBXiYG5daxD
VaolcFRCKCS5UDJtGHAFri0wfbmVutoGzcQcWIu72pt2HojQh4XcDPPT19LtUd1RwJdUFbdsadM5
7XCYVdhYYK7PRUUVWbyY+G0WlK11iEYIKiNwXvP+C62iAEB1foJbTJhXRxey6WqDPU9kxjA6UnNw
KJGCoqUUQlt5qYxYAsYJOgkHTBAG2XhnHqimIxir75LY6hxq/xUoQMUo2qkjnBp1GCqr21WT1cDC
1jAX2R7Y3no03Yhx0+EX1Ya0itRirvId29t2O80CHRaDtXAllW0MDDcO+9L8gOSuVteMg4Bfybok
R6qTiRnrUibTLDaDHOp71cGNGti6h8Z1HDTlEppnuQPyhKhpgPVUCnIU/ub68FnE3GY56NNz1ZbN
K+6KtXAeIyzqszoMpqwEDeQB1RG1sDquHoQbgSmoX9bVmTjEYtXlHmtQ4R+qeU0m3JIQ24igjyop
3M937qtUx+aTpML3S1bRIjS5dTgvv8Zk+NWdaNLOjFr596pIOCePYkH4mZIVZmfCU0wM8Si5v0Mt
dcKC4OpWJkTuCPASpyYgidoovRyPIDGgEHFA1fCW1WQkUMEeMs8c/SkalUFM4AV6QTiJWAxCsPLD
Eqa3IEA3s6F59dk6mK2UFsq2vrFbTEGVwmrCD4mkmhlmn4e0kUgAi8Uayqr4yE7m2wr1fG6XOHPA
EdQguJ1bnBfD6EFNKwC5ulFJ+m/TKFGK0TZ9CdTJCp0vxxgPSxRTnaZ+YTJWatXE1Ar/FpHUcsbD
BJQjvbxKcXrp6k7isJIabIBT7tJ7CNLqUa/rn4mf/0qoOx1Vq0mQU6RRJLGEPaJTyJzUMwm0hZjT
JQsjL3E9Z5jplE8h0/VjkDYUdGFI0BrW/DL3clBwhpRPL+mMXyUHQsDt9fdIOzonmZ6BIax2eRDt
Bp2amCoOvUNe7OFOMThPlTz6Y0FJbNVxVu2rGiXWDpMjXVGxakYRjjNBe0g2E/iMlPxF0ZDUmYVc
NWDFtyMT+VBiBtP137vOmnOlqvxZd7Ds6+3SFh554nBQrEJX0rSuIkRcWiqaZ97PJqhzn3PXNWlM
lYT9iwCIXnPdw1P0Mka04G0tdjiaXYI4MhHxl8D/kr/iNWx6nC6XFTTz8KCZdApcyGrM18I1SwGh
wIlw58p8nrT61rJmfEx1pGRSu3PWNYBxPYltd1GnFOeA6KBmtNiJDc2WU4BJ6IAja/256De4bg6O
t9QhPcnLW4bsG8B3J7GxeF3A/B/FaIUxc5sDxcgJsozKme6sU/qxJlWR/ThyQ9QEOF27VNwsZDW6
8bNa7trftQQM98+JNeip+B/F/TwXSp50JKUUOjXmcg24Dy0E1zWbtFLgkr62uXejzVS1QXu+ubYM
kgLk2InewN70qy5tXOznQBulA9s0UCgEljx6YPLNI9LWxjTXyGdFJL4dVqftwS3tJYSNiMAWuL/3
pOz9RjeiwRveUeItYlMOKZEWzmHnhtH1Dqou67Iy0/KmK2AdoHOgj+Q+gSotkOh9ZYyQ6EjUWdJ0
Esf6toKXnAUt0kvXvWTy6UhiHDL02G11C8mKc/Z6O3CsdJNJlIjp2zCclvdv061/wywtJvwR6Isw
uVGbBLoEmErWBXlCjOvzE9su+qR4JZl6d7DnBHH9av0VWIUjcL4d8dHpqho5T2u78ip7K3En86D2
BQWvi8F/caw62LJtd4Mpdv2E4EoBXx38VP+K4A8LbCyAK6HIcdkjmfm8MJlys7l9h6b+PXLwkGUP
5x0/rW4eC6ER5XUW0R6BnuMOlROmjQNSCzbOKFi6bmN7aHr7za+1WTqKf7lGSBWS5Xe9xazwNgDM
iONcrdKX1vorjZWlqmxxD3WiPOKgUS3SnSbwdtne/0BhjnYwsAdVSh2ymcvCicsWA/JjJTAp2aI4
Ez1aIPvw7kwVgBt964j9kuttgNMpSI3MZ24VCW5Fl3dgp9w7HdeZHiGCeKJksYEFW4/8D9KvruLs
IhOs1mVurYMe4j1Mi0DMVZWie35tNxtLSCYAIfdoWK+ug1rOtIuaNyayMZ4Nrmc2G0NHCF6+Y8Gd
ASW8HgkI4/8U9iYxukb5pjpjaGBpOne4NgMgkKwFPBXWcYh/KGfUC58IIV6MxG8ECldTNB+pPTlY
itrPo5DGWHcHzMG+dgm18a45A5fnE8IZLrvCU2xie4pRLLElRde6ZPRtOm8rnA2BaL/ktF34fUgV
qvFObi4X35OxM4gUvs8Dn6yxd0iVokDFkCw/lFUxhczKjQbC+hSLYmq8nzEN40Y5PAO6WfuO8jJu
sDKj6lFi1Cr+Lpa6dxIKW6HKXre3VlFHQkDex4UDFfyd/WyGZHrrDujwYIufpmCpTAosGN9X/A7g
ggP15X19N4CyN7p2jtVYw/2zptv0p5JPa0pFENtC1+vgTvhTPLdRv8beza4qwccJbVExYvjB2skq
1IJlioafqvcZli9wT/b9YlaBDvYe67vhrfnnW0Q3Ej6MLz2gsM8crlwz9DDyeWMM73b8efKRkNdj
EpCjYIsgUbpGM+pnNH0KUL6nSQyaIfpDWyXyap93s1Kz6xJlx4CR4PTRr/aNVUkZF71UiYMHBJbA
c9DZOxu3jD5W2TJrZz8uYBqxQNRpHawPun1n0uSBFoV6KpIsknmgJH9PMuGGu9XCqwvELFdEYka0
r9AxOfytRemqjspN2QemV1dPE2WQtdXlUo6y+0ceSxIt3NQsRWT8oLeHIQTCMezGIKl1qAf9oMJc
qyiCL5zY8Dh2J612ch7HHe20SrZ2RMbf/pqnYryqF94FpHXF+WYr+/L3QDbau7CxA19XsG5bR2zt
o4ASWqPMNJMwVijaNV5dSBKqwohAG0+/OL1mAI+1peqmFopEBnn8TcgBBMrNl3KZ4oy2jTzwTvZU
Gw4f1NfGql+vFsmdfEZ+eYwP5/dnE9QPXAO3Z7lyVfVaPYJnYFTrtXb1SujZtMGD9D18xErAwz8X
/ngEscMGStrHFe9S9byQlSN7eZXFZFtoAvElwuK0VPq6bnG+d51eFXR0Irz+5ogrIUFoQQz73xev
S7Mk6PnUnnqxyAavcCqpBoDiQumAUEm5o78QFfaY8jpxaVG5pGZzZg63iPvZsQFvDbY9qlXwxpPm
/fMvJ/ZnMWIBnv3vQ0lOOw62bIY2qUaBi9g0bzCGAN/5RjspopXsmOcq/Axmfg4yndFPl1hpVt79
vsCUe84dPmPmoo2FRBVjiLvAafmUBfpxA1+m6Mz8T6meDXohlqAPTugqsOyXgTzNc0K0qbtzWc2d
BtK8nA0oVVpKfHkyc8P2ptt5LBi/5npo+c3TKLzSAYsHBD6Mcenrs3bvyRKrNduLW/i1r2A26f4N
tDsY1dKSoNHBDwdmSWC8KDpiSEpf/iR1HE+XSOZt05Cbzenr86IwEjfRKXRXUmnCwpZio2fzWk3o
DmHonl9SlNVu8tluCKp1vyx8DKKtDZhwuraKoRjIBrouX4UCwvVVinPLA24iwicn5MfAQAX8xlGI
YD3EaeaJGG5RnnryHxL6mjpBKmmNp9/j3C0r/nzcpLPi91MTbX+lyEKwDQBXJmrb9K92iAeKRxQ3
lwn/hs7hNnEKldSc46NRHmyRuteP7DTtSDbhrJ9DfltdmzmVPsdsjde8Oo6ee1cZXhWW+Ovp2t4P
GR1YPwHgNjtcYt7LUCbkqkyijrg7CBZ7tqhIOyIIIKA/DEwJ2UAGVJtEKCH5iWBkk7K0TXeQ3rh1
UFjYX1ZRuIbn+Qk8qzYFOeKvS36ZJQLT3I4b5aOajz6KIVZTMlVhsh141yPAFRFYxZuSbiABp4Lx
AqGYi6Nrj5ZlIkYI+SpX2M/aFPCCgoC/duVKNMx6GbyIBi9YEiheyng4tcE8QgLYzu6JzXB/xl3S
qf9LNEUpyIAbk17EE4pvjsOxlkysdsOC/ro5E90atSVJ2b5QKtNbrZv2eqEj8TC4Ml40MV+ApmIv
5uE9kh9s0J7uWSTz7gCBbPX0iCBJSh/vzI/6T+CFqXsRIfStHdiw4LkoKKSM4VbyJrvMbT0+INWm
wfbFxQ680k51zIXoW5A2dxTkEoqEnVQ0jIbk1fXdFrI6sshb1XjqDTan2+b0qmsxOLpGPDnrUI5v
MxVc/7GD/IjwTvMGwknDUFlOcQPFGHSdpVKYCgvSB6VJFbd8xTZduT3g1rPzwj3KtekejzoS40gF
Ks/zJx4KY3SPMkhzsR88PVFtfzp4aksTKJtIrdcnw56eJi5myGvrkQ+Vn5St9b/7ztsaBcY/UsRZ
LE9wKqFQr3Izqv2Jw0h2trgy5JgB2tk40mVZE46ANKoJWRG92g8QmivFWRr+LJxIeU9j1STDVxt3
1cXtAhd+BBUrZG3L+S4+eBEhSVonxoTXBIcU60G2onfp59jw2hibH3mnDISFlsa7ZlQR41i8K5OF
ImZsgk4Z3MyZuZ5w7sQY3nSUgaaEQIftZ9Axpe9Ew/hYvVY+f07g+lrqPH6QcCWOuj7E9Jg4RGuM
0m3PhFJ8mnA7qHFoOlcHWvChO06pB4u7lZx/oMqQfHp5g0avqpJVS4zBrXuE/0A0agGJLjIBHOlB
2f6ghHRveqSOq2FCP+cG7fkabAivl7SCFhd011G1o/VqioDlFRsixobtWflMdxpu3rrKnPiv8Hoj
1p5t7TpMOrHkSPpgUtRhjrj+ApjXBbQtqNMYXNWbkUcZ5j17a7EIgCVXFJzRRztYmBfwJD36rCX5
nKQ9s0KwN4/wgZH1olN+WqEbgTu5ezzqsIBtc5K3tTJjRZcCZv1deRYe0H0Ik/5pUQwUfxqrM1e9
yzsSjwR11ReZqULR4jZ418bCrKcKQNWkdV+uRhGe3zY6Mir7SKwNBxNLj0Skweq5CH6OD5JHWZ2N
cGUtLruFlCqXjKenf78lyeyDasfZ998V09aOEtgSmi++L4Pfl+QgxNLe2fsBXFq7y9j/kjDiE8uB
GV2Pra/zYoTUfkDsX75SJzkFmRfMk5NwZiLI7XqkIW10qWV8yjUtwxCQ6PDe8sIaNUY2Jr23Cvjg
Z+wBSe4Wti8p7twcjwmsemyG/a7atGLb6aK9gB3MTIRh8jShYtMndGSJjAKnHncvgqUUGGUaUd+Q
cQtyV+HppW85GYTpkzsAYqsxubcEB37JPGlKZLrZ6F4Nyih1mDZ/WcxD1VHh/Uiryd4Wn3ISuaFk
fogqxMBLAejz1zZVEIha9zGOG57LLzHl8z+SzlrjSyo+tsxgn5k8KMrc+8AAAngW0XQgRykF9tHO
aAz2rqbG8NoqR+Ejmlp9TKSZbAnW9ieQj1FNNMpxv7hRopTPsCWEGYCLFPyrGisZmHGoZ8ydNVdJ
Rlp28Dj9nSa+xrDsCzQ/5J4uMbW6yrQNNufWDdbmlr6dIEHefeT6mdkzS+/zOLPXXtQnaF11laie
e935Weq01Z72HaZr1UVseUgjHRJpT+NJrtHkTyTNc0GQggOpxmXR2T4ITKSfkBru93PqG63hx1pj
yLd/ozxlP0MkxC3Kl0B5vwvlHjdmzcq0DTQPb7qEvmqOjRnqEASLkFaAGN84x78P4irLI0L+VzTf
E+y9AVQ8zIXFOO4HwRmjbyOgr5lVoOJDuLkeLA9iEF11zpGsxaUiJB1XJ1F5Hd9ZnqQIL1pV5Vor
2AIUtznJwqTv2l1suWS40NdgLfeTeO2H0U+aHEM8Xgy9wjY8zIb4cbcm05yAoYImxDF4AqDCjTLv
b/MVHak6K4EMs3snEJe0ydVkzAVnX8n19ltXtcY/+/P0gprUk5rGe3wmqlKHJpzOdHa5cxz0AXvD
pB2XnSmqgG8hsY+cjt4BnFWtpwS+G22Ms3u7HFdCihnr9j/moxzCYa9298mfpz5KrCNE45GNmfnH
V+EcYWG1kYUI60/56Y8pVOuHLER/o7MxV/W9HlYoqWhGo7fr2SvGFEVKdXY88bGkBJPzlMkqto+n
f0KtamJ8KVNDV14d6lT5OPJRrmP1wWHp2kTNkRxrZvle7GAcsLlsyvjogMSD0Ad79W4Hb1dBrNFP
ykuCUh2vaPbfCsRGZqsMNqt5ayVamD4+crjVf5EALeRrSPz8DYDVt/6FAQ9I5NkqLBaG2Swru/Xo
UTVhBjWcfVo0h/6EgbhKp/s5gkMt0IBiCUBzNexwQKvrS6oqug6S/ec5zP8+rxGfuYvH/GisuIpB
63t1YnoVp+wS5aDbUzBVA31+GKkbZ0zgBqo1lXEDD7rt2E7iiXAMmOOXgTSQs3rePZRm9w3Hp4iK
jsILiRZ+i8IaxjqmECXn+FumVDesSAcvkoiX5YZH9cUcn+XBwuhkZtGvfhpbnOjLu/OJ1sGJ9tu2
UiOzE8sJPOufqXWPvco1KdwV4PImU3C+bObTLa2g7fQOiyplgHMwGGRscN9+TNlsvY+mY/2N3paL
Fr+E9rjRxgUj3hubGEVqfO62KpbAhyycW7rq6q408PhhRwuL435nz3JjXtrKGQL4ZDVGhJlEVurr
h/9eFnBXovoQcYhJLf1++RGbGOtKB5ErZmy1Z8pN6vZIdlc7Dhy4VwbzmWlIY5o8vOEkMMWnextY
1T+d62oOm7wP5Hg5cvV0MrT6K2k+lMwPNxVTriUz3FjzycskCWCKy0QUacWRtX0Mqzt7YM685wvy
MnewetlAmdBCvduS9BVW4OXsWvlvcOnsmfhH3VBu+b+WoXnCuG9df4PE/cV/QnCvm9504XgD75+x
8Xt615ex2G1VhCyaymOBemTTMx4HoENS6IyoWOVFwAJXLU0UcWoq2QEZzeeG/0R0ztrqRPKpO98E
+DdkctbMZB9RAuuHplGmIKTNLhHJ3wkd+EEAbPGs4tfJrsPubp9bSUi1R4TjRHqZUGo/EOor5nbJ
/kOBzhlgey4l2Cf1hZw1FTMJ8w1ex5ZNs5euzkJC+W8vyNlZmS5+PJ0rXicUQ35X+TvH2M7a55c9
UbIVF29ej9wrEjafF/pHXVYIxhfCUZ6Fxwv/hm0bjGp+90Vy9i2HjneK8SdM2zJrbUe9j96R9NXi
uCKvG1ZqYGOZvR46SYAn1RdYhd98LpEGb63CDpr/5AXw4uMvaICkCfRH3h2u+5mDaop+tTnOwxSx
G8QnKgBgWDVpsU19oNq9NNXrajsFrWNQZIkNLrJQAlGsKqF9GPO2dlemIJZzH8KP0eouRHaggzBO
f1U8gFA7hl2szYD7g2osdr8RnLG+8giZQu3roJMGqBohqx2KYdhvlPZb84adfLCzT1XDcPwxGX30
VBwzIHaiJWFtraKuSWBVoBgSMzbrSIBkGS6F8UAnnvWp+IUmJC76SpAM/4WZ3adKON92JT+bm+pk
+kjcPYYrn+e0i/wKVkUTEw5eawFseyj1LNbXkOfLRHjIdbCBbmoL0T1B77Q+NlfncLIduhkgwll1
P7262A5QDykwYsd6df1mVt/TP26Y9TcFmG9CYxkZFyVrmn5O7EpHzmsnhblXU7CN4i1VhYWHhydD
m4e55nRccHmha6jsuxNXDCndMSxEM1yVkOLYNr4l59SDnozlRIAmBFT0wIPBUI6uZqSdQOky1ZkS
CkeB8NTVDaN7DzG5Vy2XH5C88NVkfq5/F9OlN3SNrEUr0SeDRg6m6iThCZAXjx5lalxNfKfjbNcF
XrCk9vAmwfzhLwpd1xkLblDieaWchwtk7/BDMzCHEvmx4pk8gAbcbnl2hKUjzZYxUjkWQ3yQhuDu
SKZzlMoQ3wBavR6G/YYhuuZyWzVQUTDmhM+TO7vsqcFSoJCc876lpuUvif85ni7rAxLHHa0GruWe
KrOiL5Gcl6aZL6pT1JTeNrLxuFJqVlTJLzPosdBtZg3trqMHi1JFK26h+pfTxhEvCzYnidoaZ9XB
YBcMN/iP3uv1Q8XLO1zvd+qBHlLaUwGlPpK1sPJw3J5StWaV+ve6itm5BZKsRj85+pCAxwB/dUm/
rSiZh1NCEH9RKH7xU18Xa8MdObYNPDKNEo9d4OFNO8sVvmJhdPb5+Zb5IcuiikT5GsoMrfjJGasX
eiTCNwVjCNL5/FeHj7D2Y6t55gwZ53ybIGvWjpzJ1xA+fJDySgyVht21w3w2OJhEmo8X3f3Sq0SM
0cnK5v7Rh6hKZeG3zzoboQDXMx2an+Cjxfqeo0OVdJ0OmjaN2fV5fJNLp+lIbrw76azbUeb9ZGIL
4t0pTUEr862vz10YRpdoJDK+StcfJbEfJXkbsJgKMZelDfv2NAGYkH1JcpGLGrBjrulMLpvvSP/B
hhUG2QWBilt3zXKvdBk/cO35nPrS2vQMAU8hRaNdM5ukOS9R6MwvXj2hAws7zMg7XmB0DAo/dKR3
qxMli5fHH37+QKiRjEbnivFlUGqBJuDFjngZSwa+CzdAj4Sw3e+CWY+Rq5aEIWWBocVjCJOgCUhs
fABru4PUF6dfbk9HzP0PQHGxAtz1k42Kh8V5Ogcl10lGxmXwYXe0FzfVvZdbuLFcsnf1v9gFfx5g
IgNNAhGYD3JiksTrIdJA4Rcowlxl1twSRc9KdXwoIpaRkAxdZOcvi0u1EMHw/n5uaylOsBeYVlPr
ocfJzdohUyucVDIRJnLq1fNCc2nYxvFC852oSx1zkjJdKkz+d2FxX6tfaWBrI3E+xwu+tCTZgWlr
Y1ItISelz4/WWjIFh5TkoNYxNsOD7GqthC87kB7rC1ZsYGpiutUv2h3lkkAsB+iIm8hT/eXZ9xKc
hJtmH8S1MYmkfdFPlu5g/mMUeEg/Or4CCWgb7hF1WErWEtNvrTX7Gts8mAOhxEEkYNz0raAugdV0
2AbHAW+ojXNrCdOw/r0B75clXaAGjcKnD7wl6W61p5HsZzHhudb1yZUOqnnp8Ffc2evoNRwRW+f2
C0eh2luNX9AScYJOK5fOWq35edna7nQNz8dVLmiKIXDpL1AMj5GYuRACbRNLo9fhI8dIJwnf9amg
V9cAGy3kmiT9DtgwN/MONpo4Axh7/0S4og6UV4FJZDROF0nT95i4yzsClPr9K+PtyY2x0IeCAtA7
/qfZxodnjvEvFan96KJby4/mSgLdy5gNcUUhuzQg91tvezPTNNHo4STveH31/EuuVulvKTtOUcXw
0XkOa/gj7UhoPkIYsS0rXEtrNgvn4edOazDa3lU7uKOfHWY9YQU4An2prsVtLwgbJAFMlhWbtncr
9brAMNcDH72kO/GAq4OkoBKcEy51BTGl9R0hdmewnxUxAVtq3c/bGgiBnYVhLFsmeBBX7hhokz/U
I0de1G4NIcOY9oZ0//1MbXlu112FVVuucNRcyMrbnzl6rPIdj6TQRlBM2pjSXHxkgDg99g1kyoP4
v/M3FpyzaXRviSty2vmB0GRk0ThoPx48PGC5DXiL0Pt+jNoD9tNLBvCvMPSuFWIENMNT45oGrRTO
Ul72BwOCOvi12sm8+0W3npdsMZHOvlPNfGpEQ5S/aZp6qrBQZ/rN2+Q8y6Pfy7AGS16Sxvy56PZp
TXjNKb/9t7wLC+lkmV2nbh8vXt1afsA57B/yfpw0zMm7E0PQJktDB3u92PRHzOSUU6UOer0lVS9m
2X5x7owEERa41RFC39jwBVvnsA6ehep5+LaDY3mo6QoE/tilosD/YDdT8WX6FUZvxTQU3FGr1hQ8
ryGEfaVEwjcetxgBTSBs0lQVsSAxeH8gFBLXH6nNZf4BVctcvcs54pNgYidaIdBoOJkORsZVdUC3
ZxKJQJyD/f8XCNI1uyG0wwkI7j4f43s0nqmvacCrG/0+2m1PYwO87FrFtowyVasHNcHLUvbjPObZ
n3z3AHTDR/UrZY3MNYkjNszNMfbnag1VJVY728+vGoAW0dRwWMsLTrdJHxREI99O18Ij9U/ejfM6
p5G8y+dy2Q8EPi+4NCPRsysvvMxvWoHfriiciE83HepoOop/kPm8k1ipwElC7M4JQogekwX5YR30
/Ue26AqJY87QTIrRJ50xg6zyhWzKg1muqTBOlcMsgRdDsdqf4nqh+2SHanKs9zJ/E2PhubEkXoP+
dcicZLpeRCBzVmQuLtQJbvg4sruNKifbMRtCZJ+vhuglcGe2lBi7qbr04/IHF4jZH6xmtFR0IZtm
pbxSjgfAVIXVOD20+7JDqpu1ej+tOCZA2JvrRdP4RNRMO8lEyj6RtQfpoJoGfuG7niO/0ON9VXFt
vfmelBFBiQmIRuNjaSj8XJ9iUbyZhfwqlBHTWQLn2dh95eO72y8QcwFkjTSXh6jqN4wLSBKsnPtP
EsxWOIOu+K5BavrmRHlmBrelgd8R9h4ofrqINnZVaC3OhO0oTRd4ybIIcNfrFgIEC8slVSOSOoCz
CkkYZLUpqO61TLXLm8UjhbP4qaHYdGB/IRatUoF9VCjxWIxDtoxm0f4wKqYv0gDaKhaEhshrkMyy
iNHBLmTe8Vsb/jdfuCsMLQ51GxBLACGDHg9wEn6qzSMS45Xthr0eONkeBtOWj90DtKYL67RfRwk1
+TNc2lFkp6OUDSibThLblM55RUmTdGdp3oAkdVXwtK7jEPowuOQvip4x2kxEbLcUAiYvhVlF42D4
XQApt9w0oAIRVls4TGiZXe3ksPg0JtAw5cDaBUSzCldW4qChuNbEFLhzpOcXNvoa+yYjdYY4POi+
wQlAG8sILOFLS/ROdo1dFc3wl45SzpMdP1Vabe0rinoWJF2JOzjXnpZf2JVflemVEGn1diI/pdtn
syG2uZe343Q5Aet8XPw0+/mTfqj8ykY1YBIjSsn5hSciGkZBhws3Af7d3TF41vl6PYOvGZhLrLET
kXO9NeKEmTfmAYCVBtfJFytiJhwog5Z0r1o8nMShzUEBGeXQq5QaoXB0HVpIX4fFFd/2axxKlOG0
mD3KllawLy/gmtTkm6s587xBab4AHGtpFL/tgIJVRHswBTuM+iEazzTkmIKrUnoM6dP2CFcj2PQo
u6F1GZALiL3EkxC91n6ttCpA2fSbWgIzXNbqzXSIe1uCggQpuX57moRmJ0AQ1gICMyHqc6vFSsIx
WDqnepREoLGht98f2QuqyTfGZTz6Ad30O425l/ahehZzcZdau4vzv6yhEP5z6Sl2l5ZRvIinADq6
CMsegtR3ixFh9J1WIXUxYA6IHHLpo9sAqUNLORsl9YLQFUmR1rJvwK1GU4ANmCwnCwbonkkwrSrU
YyDumsd8OZiP9PsZuEvc4ER6DaHNfwKcq5b6V500BrpBjEG/cDT/Ps9chnzRrlGc9S2v35iBG30C
rTzILfP1e4oLuunlGEZ/K1iTwAGaHa4SaOvd/tgv2aoBt0b/WLHRMjeReo13F3mESw09eOUKrfbL
XAUbnXCStfF1xK8jnUfKahbku4dbSj4u1bKMH3pOyOIS5k9qaenGBfobtekrhJ429c5Q2T0+zvkI
+aSeGnaPQECksYkRxooSSqB/UEBxjebc+somTo1hZ2zjB+wf1swCyYOvDf+BuPuw5NV2YxMqX0vG
Cc0cZ4W5PiOsUUaZ2f3ukXEyQSxsUvFxSniB1J+QAYPTPYyUHRfLXGz7YrWbgRhYQI8urpTokoeA
gB+0w+xO4DfspemNgrmqyKOTp6UNgN4E7MU51ZiB9ZIqIHa+hpzViKKEcejrCwOej/5+cpdXqk/Q
X39ttCpcT3Jb1MZOrtgQb/0PyxtafrLnm+L1WIDAbH82rAjsci+PNUcGp0QVOQdP7wMK7g5Xm2b/
YN6mDE0+1Zk/YV5qXedM6+cQmC7BS+eU+wTsC9/h8c4rzd6iD7icICq2YBh2rWjKWoQCwIuxugo1
YfaH8JhcMbmmToNembLKnwmGgsM6RKbUucqasr3i0LN4O0cFhoyicp/Vlvkp37QPihRESW/L0RYl
RveKQdOOcB7oqzW8JRY1a0qrko9M2IirJoDBLh88crHasFiW9VH1IWC81g7j6Wte9NQo7VlNIJK0
X9YTi8mN8w/xezmWJyIdEP2sNYMqVprMFlw9wQUiFEfozRB+d3TrmWWhfGAMGoELkp/iEgSMWcEa
Di8TTyOoG8mzLk+GTSH6jcME7xfCL4fijnaeZTRCyeFLgNkW8f3hoeGWnO7rZKQf3aty+woxxd9Q
D5o1P7mm5qgoWtQkbi+R1xMb7R5hExhY/mAiu4kRSmtYNtbeTBbmQ613fBBsSZjNz9/RGDA0HVyG
v53OdLSpauSwWPKAag///5TW9hJ5qZMrvbUAMfDCHeaFEsuQOpSb1MCSXGGKTAe3DjTcpmYwNN0G
4L+irQqwUcoGDyo5xgPk+KL6Gz8HoM5nGeRxOOW6tNXmz09WVA8Sp71HV0zpzY+atEAX0U13XMwy
vlHEWe2sPWwsIxlEe2eZfq/NYZGAWJzZFC72KE+lgJAVeJSu39+Kp8CJ7DZvOlNWlgzN+ZNKaRLv
IBewN37gbG6yP3IEnEgOlWbHq4RJmwGw6L/X7HE+YbWuGK3HT1OH/vqH+VomkcfoNynVX0eoc2Kw
EKJRyGPQzBw2QfdpBtcOGPCNjT92xkUngFhDNrRkuc4CTSyyOl2JqgbOxDAXCdRbwxet3+UG+lfw
i4Ugdy7f4vJCUNbPmw4SolaIOrC59zXfxM0Z8+KEM4ZRKrU4RDsmDK4JzC8tLnmG4z/ue83yls/R
dBh/U6PucA4cFzoKM1gCshhvVy1/P2YhRhxVo/UZZfq+piSBTDMfco/jqOBY4J/v3kDSFIBE+hIy
GVCGnKX7Z+Z4s8qrijmB9htIewMsIFCIXTjaIZwctrGng9weXGL6rzBjrnD+UsyqVOSxbPEX9Z1x
H1JTkDP+lLNBJKwCLLjSbZe3WkdweMfsGF/8h3BTz6YjD2rUFHlc4VobSJ8xcdPWcqURHW8/M8/P
ArIf78RFE4iBxojkR3ZuVNOe7xDU+IkYIDK8D9ojuS/nlqpG92IwfniJzqKkwcxRu9BvNdJ1wrSx
rhHP/OOpm2bTJufuaVaO5tnqqUmhgYbQND7Ni4t27z65W5/V7GXIT+ZZccsroifAjGbgLWEZTP6n
y/r1Rs0NmUy75O0qf/cM6bz8SvdYkz6nvf+Q7XwKfp4/hLBo3Mckc40p+7UXNkZqrlAiTmS6YUm4
EFfpwU5pLPUfEIIyG/z4MYuxDCo4tsTgo4z8zM/72RjrkpaBpcQGev3K8gKwpejH6RD+vAOq/PBG
6DfWueyE0KgUWhHG5PblwbMsg0VXz7RJnz1Ne0bl+EyLs4VdesRzUN6s1OMTVYQx6a2PaK7c/C8N
uCrHqHgiT1XVYWzPSOnfpPyvSC1WUa82GVYmLjitv+IKt393q1Sdh+TB0nnM4eRovp6zpuG2RDEB
9ugiv3EmQGzY4Z3I2kJ0R++2b46X30pInODgfzlgc3c+depILoqC64BrfdgjKkYOh0jvnzL7P4Kr
g2dQwZaZSJNgZfEzstJHkcn1CeozYG4HVW+Kq38K3D+SaxCPG4GevZjeY2p7QKdzzI/IKKmIktQt
TBX+jt/VFN6FkRtfaa392ENtFllYqnAGM6TQBL3DAJ7U3tqOBSG+GR67tUNlJJzK5UaXm1bX3A5+
744aIWMgbm0mLMo/WHOmVXDTWkrzbyHXaleb0uvkowgCnjiqK2rHkv3Es234IuCG3Fgf2+SWhsDk
qzhLQMVGQb/hHWhiRXPnheN7m99hCY8FcklEqhU26Hd1dmqDMuWXBFgwuq1dRBT6o9QlPZgvWtBd
kpvXVOcxW5Q4IsR6qUYPCmJ5K2eF1ISI6FkhZTfeh8+hVAQDFxRApsNAJ3gRFKauPM/FD4nYLfPP
f0Rygk2AOPCWD39P3jH3gmT2h7Frt2d/KElgMDugtUfMtTx6C7vO0XKSLtENsgcIGurclN9DLXDJ
v9SeRMBSsl+c4BeGTUa/oipHjAFFAypLxl1y8XM72PWpR81+i79dUYNHMY/MdFddXXNAIKU0qNO+
gNhVJA8W4G9iKmUU4HwztRasoCc5CLOWXVZSUg/PzqRW4gBpvJzzDVgPYW91i9vey/tBGVPMHnoH
O3JFrFrrKzXGFC3SE/MB4bBXKyYMcR/sIpvgesaQ3PY3fCIjk34rIvlA5Z+mULH2rOM9rdGJqJR+
gOebJdSqdorJ/IZU0KRJQSip7iN6LYTwO9z3r/N2VI0gmMg6xGk/yD1KoraNG20AFc8h8AepG2J9
8xDAPXRIPTVLm7sdyDyRAqGe26IKmaRD43Oqd3TI2Ma8lT43jEDRibUiSfVPbiVQcVRwSxAyGdvj
N/+KTGTUHbL4p/9EnD2kvLwyEDQh8cpeYRSkJKxkUyiL906XdpUp5x4SwX6XqlzKN2n1avwGbPLy
gB7+e/+p+CkByMmdL6YkCtv+DBMwlKi4VL0orQtyRmldbP1mWz7XuGiW+XmGE2zGkKEeSOyQsAye
ihJudxXI1ftLLFVHAsOAn/+DY9p2K45Und3DLZ2/AbrVgYNh2jYJi1R59Jmde7abqtgL1ULjPL1o
KWXZkeviGSuNIZ+8juLQIE8FpTvarlT8LWRknhXO2FR2DM2sSATLNNiwmRzghPK/qmU/a/L4AnwI
Mtjlb/e8aEoQhlgJONgIM0OHZnyr2zP2BhgceJ6ILZyH8bB+iFfWNR+v6IFffcRaqTLdfnCr3Eki
0WiLVym2IaISpVwuz+VoTODw4xgf8Nb7e0AalwYhpl8KAR7x7KvAGhyGwYK1HWfjQIO/5wYtJPEW
aWZ3ZQb8TinU5qOQ4R9o8iW6RMFb+5J4h+769NpgsVVf7uJazcnsol+1whke+eJ2Jj7dZ4IYGXck
U0cxPQjuZl2+T7XHekhIMr9B7U3dZEg8Q1P8jBy8yy9MHOWJk/W7vlwevWr1+xAtSojTw27rfZPp
KAYEVFRHPzxhdTkk5SkyLyuhcf26p2cyUxMS8O5jwUxChmxGmPJ7r4kXwN9QzpWdbbKRKjzoKwes
MOIRmhWsCbpR2qDTOiafwUHCQwUWDafwsx67JGaHsZRTWfq6I7KYAffaX3SKys1o4YxNbyBIwUFy
XcKGFP+dUJWxQtEJ3HupPqGHPT2Et3poGYrEL1O9MfSbFqec5YRFj86gCQpHAZy9M8sbcjZcjy1t
E9U3fK3FFtkD63JetSkE/WM03wHHhgp+LLKaBrtG2y2ctp88aE7+BXavwlIeufL3w+FhY1r2O1JV
kdyU9/nU4VAvEzYpvYnPWVRNvgIYhu+rDNKRdcHUMooA4pGQ4PMfCTLgZG1b1zZ6+kXCzyEmNzY9
iQMMUuuqBe/PTaD0wMbL7xiHJDI+XQHa1bfKk8zlwj1BqRszYPCJBYZV+kVQVq0RtE9LxI7+La9J
NddXt7mkKTt0r+4DLuDc8EngL6zrqd1hFsX29Vg4fIyXKtbnZgRkAwyg8s7UuP85nhnOYzDc6Itv
i/6/C7Ip78X4wKve6y92T1RdPp3OdcA3N+GlzADA6qO2xB7rIg4lTZBEArD/XrrEcKX56FM/CLxb
+ITU3+kA6732qRhSiogAuKO8vtyAxjo7A9phi0TJSklYDUIfleZYO/zyWcITIDzLwezgwwqSmJmg
pqUZzGt8tKAh5PFMnqUikIlQFV7eanh6n3BPeM9xaJ0FUC3KRu2Rh/JK8yr91j4MUyTnFua22uJy
+HUSIiC1i3l6PYfXXL8Faz961CHwTQUSL92AAn3Aoa2MZ1aIr59L2UrleIw6/V8+xBvCblT+oF6E
Mn84CxmDXrVPR4CGLf5o8NLZsiNFyiiHSbL0zmhuwKI/jUeolFmcy9eFgi8zfqz1AQhdd7weJykB
1Ze3kTXbQQNLi+cOGnBkS5atQft7OzhcewbGf2wqXUNlxxGHIC3F4hrx6lMbLIZwqlM1qombQ2Wj
0KtRL+PhUiKA0MsfPFgoGON2lgf6mCMZHOx+WoC1QJbr1uCCW0HsJIjWbKMC3OdjyUWM1TfRKhKa
H73OOzcQhRGO4JD8Bip19rsZXLMpvwQLzj2ZvI+Wz/foDoauy/T9mR20/teqM9UFp1Em1B9Iz1o4
dmnzgwfY2La/7byvB40HJgGnnAz6zLeu6BMmiFdCHAnZp5OSvcyVyUuoRK0SaO2qzj0nYsKBH6xy
PPFXCn0xW/Nl3318DMVIa2ahZIW1APVHLEyKMx1VQMA9F1Lt2R+Fw//BRZVeKAytq0Er19oBe3Xa
RZJnLoHJguUvbWL4z1r8xjbw87mlkp+t81x5FyriOencv0CkgP9s2F9JViPCtAqhZqGdasR9f5b6
1ZiiGgJkxXUGL7u0+ubUHSN49nPW13HUDO5kPHirYzx2T9qK9J//QwCmNVeAsLQL9cbsPg/Wuzb3
xLyZs4BUHW9DpqV3NGTypo4tqJC7mhmRI72EwqxnzxFheVTcuVfMXbTw5O+cGCzW4LxjpND0xR8j
OVU27wGrcrKDAzp3JHGffZPw/5vn1htrr8AnDr5JQOx1EQECDaJxtoxVqqTzdg4NKT5cH5e4jYrP
B2Vd318UlJKYsxbXC3WR/tqgWq7gdMg7WaggGLzdyuYs/4t9LikXFAzDkPTh32lNswUZWPoTkQoZ
LyLmuJw4ynbx2GxpbkE05bk+g6NhzwUwW4YS8bZsDgzqI7Cdkx9VFlh0wAsVLbhBo56Gjgu8uL8x
SwuqM3yjPyVPLv/3kAZppppfd8O46LxxxdiXnSUHhehEQzhXXrMnEtnzUkIyVwj7zDIZ6P3cF9jM
yNktb3EgAUjND7IDbM5g5H8nfj8o4RECPVFhQTZQPRpsdGP7hJLoJCTIJWpHqxAoMAv2PHLaqE8K
bnqoGM4DsnStXS91ffQl1cI1Br3Ub44Y8Tto4cgsJnOIdXgkdldTqQC7Uh9mbgUbdsORbqKghxnA
zD0nho2KSsvs0hm77IbwEP3u7fLZJ9FRBafxH9Ds1qOzaXNB7BkbHAxcAd57MX+UUSFJ0buhchYk
Pj6y3yAmlOxx8p5B1yJ0FXnDvt1qPSwlqyNyPUQ0PHo5EKjC07PdX7IiKQxYb+uAdEWIwUlJAlMk
zzYHjprXTcVGUq2AE/nu5s10e6fiKSraz9Hubn19FqFLLiapKfZZf80dbLrojJpcMQhW7hFXHn5w
Okn9PpWB3JCgHdehqIZIxSPs13x4y/iEv26j91YP/a28848dJrBaHYKJrbdl5cNNuvwuFB4Awd4J
cB0BGYCfkPXi5g57bPIiIQsrb8cYZyq5wUQ12c1zRYrh2i4P5ONTOd86SLUzNkrDaAkk3ymdd3VB
TjNcIGlbAqW+zqrgXXrjnmBXHzMC5yX/jJdGmgbJi8fY8WexT7M7QOTg9Sj2ETKbVBcEpPUBH+b0
XX5GHKvVmvnB3uZXULHeZUEoxK5FZoVA/98I3mxiZbBnD+ytiM67G3hgL/qY8SNaWUJ3gCJ7sVtM
1i/X9FjVdulQnLfNUZfLIK3FsCEYgJ5l6lgkJXZ+ADWmrY1E/7qLy/IJf4SB3pbPpFdz1lgcWyfP
MVEFfckISpah2n78/KZGgOQSo96WDJskyfcW6JfBmNOojXg5QswT86usDaMF48I/RpwDkkyBDKzU
hXzdo/KRzbxW6l3ZIMN2/zJzEBPpUHUAD7FcJr/vn/rwlmMjWC+C3iEp3cCc0p2E7XKFTT5WE+Bt
rZ/Bwiq2rreO0jrJ1uRb24JePMnfgGOygcxXwpsHtlhv0TNDLXLyhcUE9RmdHu2XoKC1o6S7POO7
dwG3vhGw0agytSNeo5206e21tANCnfOu54epjP42k/kDeGCX3atmsBXCVC+59hhFiKvJiZ1bhKds
ENM1q2658dL2tSa5BJ36hNieATsym6dBR0Gtx1xBsPX/b2WQXzy2xHkIAd7NOYTkWlaX7+omNz86
SVub0GcsHFKAvHHOvWPuJ4bQVY1r/H1pZcSRyvO3umHN7xEK0dyR6abBdoS2soBxT9WbgwhcbTDF
1vyo8P1g0WOVTJBawEHdylGOuOek4RbVGH0HTECveOkNMKaUvhX9F0A/DXW8ddSHeJfK1BZXQAaA
wTYj4IZjcYirw3XtI+Ifb6+jPPIvrvWRVypPn2K68nnGEMhxB2ila87SI0ItyNfO3YiyB7T9ZkM0
Ec+iNd2HcR23AqTGVFJfbOtTlck1akR9a/ADa4JLd9lKMt0XZQFNtlpQbu6Cv4XX8DAbh3t5PmeW
CDqVUKbKr6r3PhGu8bnN9ulPYZd4p9smpfMjRXzsyiP6VekHQtImtydTRuuQDp7Hh4SToHyJmmDE
adzj79UPjxDYSQlfDHpHUh7lM5hUWsTW1/c+lh+DlolvmETnXSXLARggwKKShETX3Fzul0z0rmVs
mIG3UIaGZ46GEJXNj5zkl5AtYp691RTxPMpAzcZePzoY5nXKgR1kyBVuLXAcWcYCoJOe8SA21U74
pH+6oiK3O8QnUcR58sLERf2BNEf3QOF5EGFoRBVL6pyy6MO59BY45NSJmPClS9b93FQiQqe4z/rq
xE+2XSFt7dFGWzxi2hM0SSoQqVfcelh2+nEiqBN8FSeZ5aRk8QUdJHfw/3IBfJ+/j3QnBHDQ4fAv
5P8bP2H+MHpnkeIVw1JgHqUBnawFQ0UQC1lmm/nuxxy/8BqUQjEkMGTVAJTng2uLel9JF5DS0iuB
w3uu74y+OIZo8v6knxIoHdwQDNDCbqU9wPKjU3NfN2NIuoPOeGBUSe8HLMUCYo4WWbLoWoyEW4Fa
YKpoMqtBKu/wG/y23uoNmgKl+Kuz6mEElzkhijR/vvrJkhZj69mci/mgDNLOH2lRlUJvBFKpxFYJ
xuXBKliIHg79vsfvxzfL1yZ5KGremKEEnk9sbAa5jGzHVNgYndOgV3vYR99RE/84YN1WJ+M6ke5M
7uXU4z5y4MOKRyEbuq5nTF05vSr5SwNAcjsK5LIBk7eRwyyeqIkGiXNUFXiHcfPNVxi5VokHvuGU
QNTK3hWExDJv6kZJW6bPnM+A91snk6B7ycSE3YqPB7PwaAgowFW8Ex9inCzaTItoeBP5QofL3wF7
qBacjq9Ot+m+NYAMyOsc/xIwPiyjZuoxu254Ju5+/TKOrGVXzgMELbeTRIZezpu5GyRqj+EDEyWo
vayhLvRL/NMr1vpedObMnJjPJus4XiY818jRCHEegqkzAbpLYpemtV1neUI20WOKJDBHU02OYhlj
hjxsLVrRPIBX9tJbh4xSSfI23nBtlhpX9sJPf7nn+6TRuUwqQIIR3/82XYmGNPPDeIlu8iHXOvGe
h600Cm1aBCqvLhXNesIW2THoDmcyv/9r4DuhMIS0vCuekLJCEuQVcMn3X5O9f4KM2aORJ54qrMwl
UrkaJM5SWn7GENQ0Yp90FZNu0w3DP1/MHsndkv5af7CzLvgUYETVUCcSzzTcVvyP92NmR7FvArdG
MKYC/BuzAm0dtfYt0IdOZZjNFrb/U46CFjfWHihXeXsQzyJYSiOUri/g70r4yWf3zuAlbn9JSaom
gSrUL1UMEHijV7QlysYYUpfNJdo/zXISl9JBe7Et8mvpak59s4GNTz5cOa/BoMEZ8oFyzfHZaLla
wwg8rq6S0TgNn0ABY5ikTqdxoJ3ygXbgejRWTk7n0J8L3+NENDfNx0Y4VTl2hoZ+atzZ/pwe4f5x
NLQLMseFD6/E4kCmwwohkJDrWsYeXaLl+Mjy07cIp4zdpO7UNmHfVkjaKBNDMyi3+zB9jRP6PhRH
v0kUpqJ14CVPBeKE1Zet+jIjyR+DabnVVTB1retxNzTzwuyxl71v6S+A5CTOavdjQ+qGnEwbqjmr
JwBFMBpariPNS6UxkOWaIQYxxu/dPWyhJRcuRbq7pYtGODK63zqPfqrgneQuRR3eWmRfZJhDo2Lk
sSjN98xTon36S5eU548kxTuHV0sT2OLIO7iw7JvMrvLNKA2mjUujYAr8VPYTkCAOVCuYGk2/8Qwd
yEEWF5nDAlZAcEFrKZDU83bhVReUE8sYmOsrT7LfaupVyUFxQPMwpUNMxEHny0KDI4FyUBkDhZxW
FjzTUkrOWQPrlJSn6DoEzQxKb/mSf/xYYx+LdNe8/zlsOm/u8MTJret6+8eKuouz/ulSDYTnJP2Z
xwALffJY1ErEbHUEaEPc5f2U9CF3rco4NI0tuQ/xhk98ecuOM8n1ZhbnolAIg/9Hx6NQR2XokpsO
Qsxif2Ehtxcr4gQq3gpLutjZj7k3pOK9EcQ/jR4LzlwLAFil1ZAKm2HVWd8/XGscB8MOLoxr5g8U
XUpyc56z6NjnUzpmeHucFbsrzLB1gwWLhxn/Cm0uw+Y7COFk7KSNaSnv5r6qHlBcs/gfoO7Kz2a3
Hj8SvOqy6Z6w0hg6MDDSMKIxG3T4M0j0v7EzXXt0gXDTIsLc4TrhzamxPoTvcpzNmrLiwdiIDCv2
m3fLe1om0k0/zJIU0DeRxKRb62d/MKEgMko9KK6EQ4hAxgAL/SwMc6GV91MY1F6zKxW3wm6hgX1b
XmR2990MI8ohb5OaFiHyssO0XISWtIOEXiL4frX1suPlTJXQcDjWu2lULSN2Qrea5hsypRZYYAjg
n2PIOdOshzv5nnDBd8oMTc2u+OrGxz6pBFYRO9J2Fvv0BhD+wMvTQOCjgL7xxKbYWYNWPltje8UT
ggyoYUGtvRoX9Fbqra3RlEpL9nW2IPxaLA9dAFP9kosk9uiFEQK5lJ8IlXOehXPWOtxY6leW5ghy
nAPQR9rVCtDxpXW0pk4uV7rtqQJTUZkd+fNMmHLwDGxff/qNyZjIMKeasT5TVusmHCvxDphKf0ES
naja99TNQfL/aB2vftT0MLHWG6/eVP0GPpxVFhogEHwpREQd9t8VdwJ/zhZkABAXsUhERqdHQQIY
piGOouAkJOgBdmLwbZWL/R71MlN07auSglDyok+1V5OlmMxWN0ngpEyQwHxbSA6+CdGuoCI9aXBY
yMopIu4l3s2T/xdkPqDLGhjmr0Ya7BAW4hNiVGDGD2kW3S1get8WBpZpwxkrVI2ary6X2DieMUi4
c/H/6y2TGWmYLLPvV+zO71whom28nkSw/JNmi2UELCxzv3ndhfngwy0iCATs+VwGBXzT+oXFAq6l
Al+OFs20jO0Qa8Kc9yaWCSAsvRQ32nl1lLHOGZ4DzPpiMZgsKLm2KRTsY9XA+HjwToInCmhFUhmS
p3Y4aKnH51/wL8aQVJ4BZAw8cRM59SgaonCSk8cffrNQQf7IkozK11U3gzPhKFO4ByjX3G17s3tu
fVZ3uU8XlbpsfkiveBhLc3PtFW94z/C3yUvi6jhchVnuuP1HbOHp3eOVz1if+0Vrn+KT32IUnTr3
2o7HoepEYUZYl8fR0W7q5P00xWQZf0qHopIKV2EgnlWwuDnegZXbNXAKdJ/JKTnvHGwy+shvQCgW
BruxLvvOf6cc1grb7Wunxlb5AT822BMd8L9g0zV/L65LJWE2iP62u8G6XlW0Lq1Reko90zBq3RKX
fQSpQ8Y5gMOR7pf3GjpaI9L0qCXL67tJPSiZUQGmCpoUcrrEgG4q16hiRC6XR42POv9CeHGWsreZ
n+XJt/yo4Erh169ocNP8Za1wwdJ/8JadrW78V9XzwWEnOhfPeyKBLvbhtgSDV8/Mtc6dAjVWGJGw
lqvYWPVYpRUmtgORKyDRlL21D+ERR0rh+rdE7DW8G/GAot7whx2zbvYMnqd0mD+lDi2gcWOH4oDL
2uhdcfyuvnyw6ZqGY1mmMGGj1dO2LRFQ4GkM6P5hAh7Ueb5vm8KvOGhJonMJiNZuyMp9yaVf88di
TiloP+JvD2woDjiT2Bb359RtaoN7goJVs3ix2B6Sy5tC30E2/XYG5Nw/MYwjZ4TXtMvHgNGfJdKO
Hm/GbVzQ1bN3HuuK3UNfrzCrC4ZsFTqF5A6CgKw387qKXfdW3pKfIlgUQmLkUFiPJYxR1mFTd8+W
/Bb/CLV5DCLWGhulB7yHS9Zwy9kj1D5TigC9xQDrdnihPjbeEawAI2qbiu3RlqoG7qCdov47Iryo
IG+UOhCtcItJs1eO7iS+UpslK/WfcDcO+LEPik8TD7LTSjoayGeQqHMjcdz+nW1RvZYkE5VCoJ73
sqioljCdV81wLGIq6zTvtiJwm+ygAnN9t+CoZwZqfhWzudV9qUxk7k4ijqlYRnBhzXYdjkw+35f9
e8UC0DVxtUeAHBO4T3VombhFrqHQRBMYoSVr7NHKbiXVKS8RZW+PaM/sPOfKxAIXnf1Ut2UB3wkB
C8wQrm+IxbyiBWcHoxVtpVwGmjtKOU0yLWyJ3P/6c01yZI0B3jTGab8lHEXSSJjvmjJP35RuTP99
yBOlSUV/Zfr8cEMcWNPpZPA1wz68Ry4stChWxSEcSLdUJyJw9kTx0kr13Twb1CmEDEh7V8xhtVwd
yMUwlcjMhh1c523c7Y6VR0sATI+6cl90drxXh0xevE3/uSWat0vFgxOdwV4TAwUhmGGQIlyNbVbI
FIWCyMxJSKcarP/uyUrvUIkOBzhencWtuultazv+rDeTJb9akRnr6LedFCopwPpzPh1bQHbyDoZm
gQc5/aetN5OpXrPQG/dTTVkFIeIOm+MO3E+5fJE4cR5+nHkkOZcpjte1U4mLDJeY3d0uE3Kz61t8
jYXzmiChb5T9Ozne9kD1uj+VJLQjzFtLao0JsEkw5DwfVSmjDOt3nUircY1hO7nxZw6l2EskL4vP
0YRfXUIIs8E+UXWEmdFQQBj4qo0V5HvdjZBsCkWfBjD7y1U0o2SRbTXifyg62IXUUUEcthO9a64M
tVHKN7kcr9ZVPwyKzITda3DDFH/ESfdydlgP6f+EoJUlVQtek0CwFF0wOM/ED8Q26tzih5kmgLtx
AGmrn4WVt8MPGg4r4DpchHlVmKeWao61LZ0nEHm/UHlsI4wqFSXIifhYDV6tcMxiX7ceXoHS929l
W75jnEuudA6o0qVzJ0SCF9VO0sdw9u6EiOqC6wQlNFXX0NAKEorw0E69DOso4SlLHUMxZq86+GzN
IQrfuhY8RRlit+f1EHMlx8bGOm5USN5GjGvKXN/YPVbuaT5U74/Kcca0tNLmGV1OJw0Rga5L//3T
UKJ8S972Xc8EkaedZhk+8ud537EnhaVChGei9DmJvpmkNiUR7pWA+MRKZiv9NIqJ1kZEd7yOPVvo
0TN5d1XmNN10htfasLNBRqr9x4UWSC0oRPiAxwSfenLufJffvNWyZRLnQp1DCZbDcU4IUSWblvF/
zyFcG4crSJjK3pUK3W0VXfKI79U2msWjkKDjOhFPFIlaH/GC7jxlufBNav+A+d4C0sffJEhNGjhR
2ihY0DOxCJZn/af+y6otsi4rhoAYIF022kYblHvxqfW3prj4t62Kdo1WcJgUzy4IQjw4/VFjA8qY
o1prbGLAsHNaum0LKx3P81oLqkSgrjj8pzhS+aDDbRWcbRK37QKY8l0Hb3RtvtQ6MSf/KRvCfjvy
kB0XdV1NQMTKlWqFLgj/cFl/KG/ygdiaHwCT2ZSt61k6BqdhG2dOc+Jd0YuN5NOpsP2oCxZSwcPa
09z2cj/kZahd5hEQ8gIe0cyxLRadc2ehIiKHD3GYxXKpaQvw8lZBgjen5Iad5sMK2e81IOloo3QQ
kdoo/h0S3rAqLmpv/nMhpsaSUzoYEKjmEIs4D/y+kJ85nFiED5AOz7uwYw2FsH+nfmpXD0hhzY1D
XVrIuBLyIWFTefHCRg07b8bLsPNv+aoyMlc80jpmRFJQjLga8uSo6O4YdGPjZP+kODf1pw8iSBn8
QAMeLtNfhVe8C/S262/bhpuQD7gE7hAMhlQ0Fqcj1Rg/sraRJjDG38ly66D15RyPo1nN0YVzwZEo
y6mnlNnDlSl82CHhVjUN1Y1qubzyyJpcTHkoFpmYF5tlRaiaUanDip1hpgiKWpsfmyGhTUzpv2ue
m4z3NC/GnDLpfd0J3izjolkKiJzFLMO3921Ln4rVurdUmFBxxWoL7EaVyZfx+I7t+Il8Zz/K3eaa
ycy8BOK9OG87oA3C0WeaBy7D8aEudy7syvFkZoLtbu9iW68LO44aRxQj7SKWJTwyS9XISR/coMIP
QfQ6GYX1D6HXINVcHdwIiIA+FpnsT2nuVRog5ljVran2fzy2fGMxHlim/nwSAB8zQa7OKdsZGsdd
S0pXP3RcaOmnmAVS2vCMl/jMNJJHuVDg4MMKNGNAl1jjkF7zMBrrP6WNU5bDuphIrk67xz0NmlcN
rD+OQIeJaX3XsI8xqLUHkglsbfit6F0VkknHd6S5/dbBrvGvvgrw+CSCuH3HuwFqXpAIR+MvWdQL
5j6Z1w86g6z05TI2gjZqjt4IvveeBlZoB5sBL/ybn/bVnv+BbrLZK8FODDobCYPNcYmBZGwEB+QM
PbzQIososPD0i6ht9PPSaeVdX00qZGpl9aiu9a8KRmBKwToXQ9Hsp0UtKg5lryDpMdLEJ24kmL94
TdJHONhVKM3i414YxgdPFxC7HwcLNEadSao8BQMIAvZGz5/n4cMt/1DIcRWVWyXa+pygz2ow2maA
OwK/E46xlZUWcAioOCaXqUslJWQR5+ryzOccGTzeBN2+BpU9ttoA9BPBHi2VJ5D4F1vsbFi/GJ95
T/+3Uf8OCTXrClKqFBUdUSdBt403emxz5qNWUppZOrnAUbXxcK+3FqtZjG3fVP+3hryukJ4g8uso
gdHgW2W5m8WmK8IShjBjwnz9FLRGT+1+V4W0mAvUZQyBA5fV4JuVZqxejyL+3S/pq0ggtk3RpIxQ
RDJmUdCq9RV0KyvqiFNDHgC0r27QaZI1VjQsL0eUQ8Rmd/m+rJNSHCiXHanhUc5QpS1XbHs0Zyzv
oEGEgbPm+dCRmwm8Lp2ILwd78DY2yHW7LxuiLTyxkVX++cXrpWin5rr0mzynXWq/fU6sQtd/OUqI
gu0D2ZiAf6322LDsE4a3xdM64MZ0+tOSYjULVlEldTjfJ/6hiYpYnik54itGAaE7k6Cy4i32dHdA
rpfdBtJaENa15Uuy/GqHNgjvO2dKUMfdjxMuuDfCICPhKOcoNHuOjakTesAJmwRKFMSRyWKOOil6
0DOysm8A8UfUW6wr5Iq8k5UVZOX80KKIn6kZO5gXJS2+eC5EcDXMCQt3IfzT2lerNjh/ceWsmRIc
V8Pj0UrKbSJebaO6sjtivvrz/s3YwSyf5eLBluFGiy20uOBLI7mymOMEqZ3EN3uNEQfW/H2AShDT
c15VmPmJO0XXIIj8GOJjW5EYA4oFqTGehSqclUh2OIdQVd78s9Fd0isXRjfTRSsD7HrfVWGQo8Oq
lLf9bLHJ2yfu2+iml3cY0KuXbbaZGg83zkK75/hl9gXEIyeEsKJBTye6PdMxo6vY9xabY4mJZEkX
VvVgvUFZqk+92pYNrL8JDOgjZZ5X8uDLKvHaHLx6wOw1De5HVkDnPdRuoTBeXTHr1SvJQYBJZ9Rh
ynNetPeW8sxfBeGw7IYBddI0eeC9yaXnoemrJN7XUZ6Sw4Ij8cXZVRbu6vwC3e4gmVR1GfZK7e6O
TltcUdUJyKeaaAal08v7dqvS5KOe9QNBQHFz/WxUvidG5VNp0qfL2TYNQWuy6H2CwNaxMefjimBc
m6ZABS7bCzwR8QT2qUZLaq0YEtLkYqC3zLPlaB5h+dHqIZP2v7Ho8UZq83NMoTF7gaA4r7tpJ99u
cqOgnJt4cPzyu+JQE0aJ+zvkOJI5SkLTKRSqaLqXJELP/UOf7dr+GmzTXnWRkyp7HdUZ1X7q5B4+
3IPRFgxRK3okJjfEGXGV0PcO8fW9njs+dZVRpqjEOPqQJl8bBEph//SC8t/wkm71Kk+pUS2DQkVy
ZejF1DE5HN++E9MN6a6JtNUTFXNT2U7BOT6xh4pDtngLA3lARB7ZyKOfHHgkS18rAOISFOk9HK9x
JvnShaemniMPG4cJYuZD652M+/RSPIE2i6pPk45j4C/olNAMG08dHXazaNnnEsAPkMxknROUqLGR
tNftrY8lOA3GAUvxBEOVL4J0CGj81pXqerD9aTh+lLJfMjiRGVD3ePeBGmP5KZGhKl3J4dU/PIhl
TQJjLNrX14qnD2icjwoD+rEY6MKOMWhdUuMhPCNmrGiHcwPN9azhEG8EPzFUzYGHlvhVA/9+SYpH
F9a3WBOZt/qpTXYhA3Si7lnNF4T9Ko1XxlK5j7WCPoyWl0z2OtDrHXVrqAetUaDCAkbRJTYqNzcf
b4PDotQMqQlvRJh6rRf8qvqN5KedjAO54R0vs0LPb3auV2WymSRbGuaLwdb978HAxYGA9rHBVsM0
cp+e+Oh9Z16vSr3Y3Vkl7/qnzyxtw6+ymx83HIxrB7le78zt7k2q+g1MIhLfo5D3WW8OtgxO/IY0
TJxOpVC0KmcJSv2VJ6SRpGHXwvSyQnviAjITgCiEZKGRZO3wWFjP7NRpngk6rm3ZFHINsYXjtGzt
F69l+Dfo5MxvRuPNrWCl2pkA+Q6GPSE7RaZ1yiAAn2GZvO2wxxeCBdvZGIcyAQXJ7NKiRkJbl3s+
t+8nJ8+C5dWrH5HgWpQHs8VU+1GQocnpkHGdn/rJ6gmlKxGDcCTA7d++YZWRhfVjIUDT9UQSbCkp
qGgUzUsK+AbiDDvbpTSGBgkrOHXgVMcQxd49brOvw1Ek7vtzIjcV8DRhsDV3XYqr6SiYRvSmwETV
V6uRVgxgXx2rzjlidcjO6fV6kj1LOaPYWNHS7uWPGkIFcUmu2WAILPy1CSD9atZj/axg5Fu5QImZ
KIizHSwfX6ZLyyUsz71A2erxqQyM7XK+IR51FOT4BtlU5eWz76FWNdoqpACfayHuRpAOrzgpGxq7
4dxLaxZRjqd1aQmGcBW7Io4KIG7BpDTpcUGVa45cEw5lJ3lAMfrP28OpiIQmlpITWBMRWlQTPBRv
uKLZpUBiKKeTNmIsDn0X5Q2pHhpe4keaIvm84a8l1zXVmigfYIEd0mSfVjeCq8VcpMgh+/D+sEuW
VZLbT3TJK29BM2zaONZ+RNuELh6uvvMdd/XcsdPNKM7Ic22GC/sQTs3l4qrnIKHGfLQ3Zt+36WX6
Y370WejRa28G0YoE4hG+hQjPooAxMwyD+krSbrLDDJRr5KGLhDcPSHJJ6DxmG/3msEVMGkf4do5C
aDTt+RfcHQ9sOSa4AdfR5WjSTs7Y64OBY3zmLS6tQUV4SLvzDqkIJokyhmYjttxnXLN/dtWLZtJG
aEl1sYjH/EQKBs6KjfaJUTdtRW6v8t+aMocYdsqS0D1ykm6bvv9tH6WuJ19tDEg3bVmwhmBvL4KP
YBiRT8r0AJcUnB4xGCxSeEafA5q7dVlWAlSSVIOb7ZHiRRwar7AX4QNA1XLQESNHrKvkA68M6aHl
lmOa0R1lGmAcabOzWHUJMQmhYRobt291EBP3X73M2oSpr01o9TBELV1Fcv9EKgclcFbeotj/jLq7
KagNvT+pTMUpCYzxV79KeYNVaB1Oisr6Y9kUVLREp6hdj7L05b2/cjsuEEYG43vTSFXhM+PNHMdM
qZ3SiHgCVkASxOMSuErXwilhh6xoOcJp4iFjQOnDWoaUmeWWEBqaXVwhVwJaxC1rTqrCZmeQ55Px
RWuPE+7LNQy1sswgJRMF4IzelooOjfnr8Z2ZniCZE/jn4/I9xwvG9SOznxnS+jCMJr8VZeQonakc
As9K9K7LBCjEuln2xc6REDXHABdiCi5owWiIviPVBKxfoYc4LUWWKgnZL5yc3XU3eNuqFkhCVvMO
qJ50CYZZS7E7ccIhpAeTJfUVTVSirDn7TUe9PoTwZsUQCyMZnOSr2Kdjrox2mEZtxUuHSiTt4T7l
DT4Opi6O+hRBJjbfdYUqAwUZ5vz3q+a34dfHD4k/MAglKRWXyjgSBzCDxuicYLISxoDhhM9dTvI1
7Q5OnswYCpqejX7/sVcvxX2d/bisXNCKVafKdYjlqQKt2pp1iOHKbHc0FTcwebpwuzdQhztZkt1L
RfpEDY8kbQ/WDrnQtn6Cx2RV/5/Rrx629EL/xPW2OzkSg7qIQM1PGnnsjdpOyZjMsDvyyHyBI+8b
19o9PLkAM1DZtyeSvyDbMfEq7V57ityrFYR+MVpM2uu48TbS+Q/RMXAazyTl/U1bdMk6qkkIaye0
Zz2+GSCKBX+S+C+y7HkJ7E/3bSfn02ELX6jYT84XziyWeArpyMI4jJEH0mDCfReTNDEHpCQ7SqCF
SWb5H6ZK64hV7vute/SruR3eTkvJO1ZcvgLPDu46sJMD6d5QczT7DrHjsr8jv6WcqyZXCXcHQ+fv
2eQfAcTX8GlJRJlhpB5cNegqlbPWeTODiuNTV+xbkL8uFqmkn3ZtR4d+qvA+9rcW0nDcPreMDsrh
9wRwDQi2c5tGywmwWOVi4Rg+IdXGali3hSZyURY2qP1nFPU7PGiaGJPGNbIu79BUxWmcnCCQTQQi
q1cLRWGMnMjohuKxkAvt52O4v793owySV+P8e0bhwI6OYr7A6OMMVbHLpzWH21RSmXvbeWr4Xd/R
dVJ+Ae+cSiTTfmkqJbaDY1/vZaRSuuKvOKr7Z11eBjhlOv17qACOVG5DjHVHlZqsSnIm4C1eWfSh
TZQyVa0Xkmneyyopuwp38d14yRmosQpE3MguhG+OLKynfP2IlvFYYPOigWd7HeCEDpOfHcwxQtGz
ktaNQgAg84dFmQUEJu6ptFMEcTIxUfDKa1OjTHL0NNIdFbEpJ0xoE53DXFlqfxMay5ygj6h+6ewT
SfG3pj7ThqHvlRaOdkjd2u6qe3KpN7IE1aGp85y6VTN9NczFJ1rYd8EleIU4LBPyUgpf0jLtXaR+
TwKpP6Xph7J5uJAtmSgDLgK8sBY/G1ZncXv33Oy/Wt+mooxSREXkYhLvAneHd/5ACETIa0txai7q
TNxsGsSp4qpkYP3x371UU1IQAvTDqWWJok/qA/HcVqhNlqBYoqid+Yn+iq9xGFXBWGSyTyunc+1N
E/ABLaQ/HjTMsLn1ehwLP3hnI43RHuApX9MfFSwtwimL0OF2U9fdmNrYBWjumSk/8bISAsgAYKvI
yd6p9/0ALamZYNzC5Vr8HUNVYf7iIiirPjL4nTb70Y36zeA6K97gj0gOoFHFJSX5t+D3p0l9rKS1
9MVcKF8CDZgN+JOptfVQEViaQ4xxBioTQT7MSkiwjQtaLEeMl+y+kQ7jLSgQ1/0t6F2IX9omD51Z
QfysG/VaXSTm3zYvlGF9WOy9uWjuZKDBTbVqKf9Vn+f//i+oUnoCXwLsE6ekqGwxhrgMVrnQFdww
NjQXU7wC5OMQxW1df158ZsXLm5vgGbdhayHrYHyB/wqQrPZpKb6R1AOQz65V9n5rRmryRCSrU5tk
u52v3ugkua6LqBeLffabYgEaE95YWrHb9JqK8PKr/z7W0M+N12VcjZd8QrNS62/rxR98LTS5hmcG
5iTNaDCGv9To+va1ElkR2ehP1LLVWXxAs4lJHTHJrUElX7Ap+XDfgVLo1iuIgmQKsJqSfasJNqDw
sgAEXsPcSlmyY3qVVv8W1uIMbBdgiSTfUdHIxOpqbXEUL6q25NOPZqod+IyQKToOGRwzLgIoNWSd
hNY9R0TIPX+qE25VVRL5DqfG+3S7OHMRPU6iX5q9h76c6U7E9ofh58M6H6pAdcxthc4RJwLE3FGN
KeMdgjxuKSZPjf0T5O4iqvQhDwG8mqE5X1ZqM3p3+l7+UX2CWcj+zCfBGX7sexoDiV+FykGWIIUj
WCTajAJ7xGZ0IT4ueWr2zz0HcgWxie89ScY8YnnfwJRQ8m4hT7qWfZhyNDCJL0d4/TUUp2MWfza7
f3xVoHSTjhSfIxKrfvbmKJEolL6gBCLqJ5B7U7VFfUzojBRlXAmY0VEhVOLkGKosDO+bbnHb678j
LNhvF4c+Wu62BbxzzWYXZI4gmrk2+uOembua/C5Gas/O0LuAEBICLVwLZFwk4Pq4cymmb/Pcd0QQ
OPuM/BFdL/P45zWnoeiI1L18dFROcP59bTqsy/uxFRfVB1aI47TErPr2Cr+lrIeN9+f7s08ptCgX
EnUY4CFj4G4EHGgjbpwtE2qtkpH3p9Kmg8xr1UvVBUliCBgixGRQVH8HNhMexJR2u2PKoBgbuQnb
gyUTPKC1KEZf2dxmnsFaybX18FLgltIe9EJI7BzGb4vNogqiUGaTImBstfXTTNp5Uv4Ib9Tb0onR
UP8yk3/pnLA0MG0nr3pRXu1x8J4gjwuIkrjQ6fjkYB/hV8BNuMQNnewt1EOb6H+KNliy79ypaFwG
aHNNmxHKIswkPDclDruCV79MRM4U8o8TWsABIKXusAJ0QKsIkm6cNp82A66HFdcya0pqBZ12p7ax
xOb0hiHfuzMzTak+CmKEsow4gRvEzqU04iLe7rOi97PYuMFMF2wiUAP4gHgQsXv32cFnA/LdIyof
EGqtC4BbRKamVHnU5UsWT1QgWOjWSbwuz7dZHu+3fNqWJevqrR2DWYFKNDxn66rmeHrSB5XRVvbi
4q8KMyKRVf9c0chVtrvFyfu08dj1iAQ9WafjVpsBU9zql+dXnDzYBfxH7Ufk0rcUh3/IhfHEU76j
+8KxdIGfSgXn2nJPKZBho4yhiTTlyKZm8Nsh2pLROwMjnPkzGoeBid9xkqI1RRwRU2EZ7cfbk8MK
kYsfy8Wkdi+3tCQuXGnGtSh18q4MVGZv7wPGhPCpzrD6DJmZE50TOA6usNlg3PGgAvb+pR1pa8ty
/fod5pa3Wq8TJPRvRCKVTZQe088tSL2YBZ5Ff9QE7H2koiWcJWeVxmYwGXgwfgG2t+PfXzU1A68B
yCCVpK+4xv5tRAZIPEFJbkM3ClRpOME0N81QSYqJ661xJUG8n/yFtb77eQk2iscQO7rwVqAQJXgw
sQyUU7qr5Hi5ISKryZdnqa3ccnATTX3D3htBIn396VK5tzcjO0xtdxd0OXk/2kDCoJP5ukLGL1mk
aR48PaKU4f1eiD3Vf6mCo5TuVTsa7hxBG/mfJuOFMO2pGvBSSptxMTycVX2L02oVgy0+9XEnhaFF
I46rNXfqOGvaPOiF5ulIfnvJA+opk4c1j4yZsc6B2wI73+Bt6a8JoxTkjFybkIrpVb32jP8DAe8I
Rpx+6KsXGujdu+HQzQIB19APRGlCTzdH92jTZ35uzlfTUCLU/TaU75WmUZ6ip792r9lFeeHaseL3
j5+owGB/XPG6/MVdzyAUmXvzuh0JzpY91JNfjq7EUEniodSylOpOBx0PIVbzGt4upn2XzaF0pggk
ev0T5Vx/tNzWif3aUKl4KK6J1JnLFNOGRU8hWLbiJoBNeqLyfJErgKbhB0q5VQa46QfNmJGw5DEY
aN5BSEq8n3TAhkC0cDcsoFjSIJEJCktuSAPLExwA1ax6PG6NMI8BnjXPDCbM8tHJDsb7yuEkBeWZ
T7a+XVkvKlbmozhMvyB1RBKI3g1TeRq32OQk0c8EyYx5MpNohZwK7tF7+l/oiDsSE6ZxvaDoari8
l/ERYFrqsVNpE0tELS2hlQ32OUdU55RVcQHVdi2baR9zDGCOqiOWfTS2ZOJI5nSHxEa0lMrJHJd2
86tA3ekSvYZQ/KV3VnfzQLAEJhFhK4OJLd4zY306glYSxWl693Xm3Xw40I7wI4DaO0+ecJc8M5oI
k9Fbcsp6nKjbrYRNcnvxrjzrVJ95Q7c154ZMRsXtkWFgCkHbA1YqO0Usii+fN9luxa0last7/ofP
0Rj4+hl2fhz+opHyCZWXdFbW12H2VQnI6vLwZCAIyQQcaC3xgcAPdPoVk6Ultv0/EeDxmXgpIY5y
YMnM8lDJz4iGPl3ZMM5wwPFaF9W+0e2Vk0pYzDur6kJsj9D/Nanvo+sVXIHHPMxPNghSmUrO2Xrx
HAyTy+nGbpbvOyRoYDB0tp31E6DqMr6xIGlLJnbelGyFXpVDKoBeABesT1vFrDClrK+TKgtfvNUk
wSsudzgyjj8C02nZiMVSmlN0bEfgdjiAKL/npQ0iGxN65/wmKiC/lp83Qfc4o2ca4tOmK+clLYMK
ZhAB2g/fWk9aDh7omD0Yrht+h13P/SR7NiR71u2ps50tSIjcrSYj+vklKRPTb0/bpLnQpqU++ESf
+2DmUgjMzFQ84L6pWdv29kZx0qWMR7XJ+P857XiZHQHKhVLUwMpPEQ0ppMn1P6S2C7nCV/wu/O04
1lsZEdm1v9OSwexgdhQ04MFMJLLRykRrj1ciXnhyH+W5MScaLPBkpatViUrgUwyGeYPezcRbyL0V
cUe6/KEeiHhXSymf//GDihYiL/awOP/ID0KV/el4WPpUEDNk3rBeP1Wrwuzwtmk9+1RkY6dnpPMH
WjvEeV1pumwtITTVyedyuzq21Iuo+h7JSo2qp3GvQT0VfYOq9NqcOXTUI3EjvP2SJctNGshAq+ZY
koAJnTAQ+A95rPownPF/EOjqQ7jffN2yfE1BSq2vKmhcjmT4Bw6llZf0IHnJOPXSqZQAk11Ur9DI
+2u+5yXyAe9peeeUD/ICwRvletMKcc2ew9QiGhjJxIfSyReyzM1PDsNQaDYRjlSaQylzlKKNKrPg
ZhChbb2UbUwfJcVD2VYnRTlPgFJ2cDFwNxT5ZL7lhx3CKjXVNYk1zZuh8kbWt3rmI8DCphRiS5kR
jL16IZGPKZWWDizs3YBkP10WZgPDNcdL1BEi+9pzpo1yRDGvPU22W4pXaRkm97yg1/NE6PitODWz
u8r/ViL6La5SQFqBoTs6hK0BYILpcxa+I2M41V7bWCBLAo792fDaAt7vqbrALN9NTBXcphV3OYEJ
pWJ6tmFd94CRRqyyg4AQYjPODkktoVOY9BjRvqEmyodnwN8sVe2C1eoa1RZiu3JiJrg3JvlCJDED
q/xDmv5w0i6QxYl/o3FIkm4jg3tXTSTUmww2P2R2SVAAHXfOpQdSdSZ9AoWRg8t7mhy0kYFJi1EI
jZvFYymZ24nTA4t0+fvt5NCbRa2ApUrLAJNiC+gSHXO8FJGgvhjIn5q6R37CWuJpDvOfZf9g4D/y
0BOHsanGhkjELuoGQEl79ccyJod56I+KNxyRMPEsfDLKf91bk497DCVItdWTQ4FJPTtW22zeLEFn
fL7q1z66u4JFjcqTYOtJ6XNflXNWhF0I3Ra+z8Yc/Dj4NbSLya4wMThNrOp1ptGrFexqfxL3BCMF
WuMHECN9y9aljDexqFsdRmRZ937zRGtOdulqdQPqWfAN7id1FmRCOlERGT7VquUR+e5AO4Y4Z8rv
+vClWfqssG3J9P5UjFFi7hBYAa1J/K+amQ96k6UBz5JboK8S8D25lkXVlKJlbQEVjK73fCmGbUQX
pflFGbOrMQSVh4Jdn3tjJTo4IBApvIYdu2RC+UYdb52tktaCCblyHMMj+2XDHChfiiUWnpq9Kx0T
B0WxSdSWdNly46/IzKUPQI8I1GK90vK4+A9/E7iC9zzO/8ytSA2HmFugGrgF7Rrff0UB+8F3/E7P
hbgWCdsMAAVgxfbJwg8/A+DcmOwUvE2TqdLI7aBwP1iC7WE2WfHpwTMP+igG8Udmx1Dogg3ggcyD
0OMqvxvawbxdYfYOB+2NswObJ7jQ4wOccqzzczpx9Gbw6yK+fo5MtINkGjFpfDopEc4UcAUxlrJN
l7MQtNyr4CCePISa1lmk7XZOe4FbJVYK5D/JdEyU6ICF5sqHwaPoZ8oedtERmbYGOYW0YNxoUCkF
rj45dyI4q+7pXF2ueQMnKsrPKxQGT8L2me4WrPDWOMOBPIRxo8bLiY9Y0IWoXpNTazgOOgeuSbj1
o1g+y6vauzpGsmcNUhw3928xC/jCFwxCvgWJlXj+HJ9Qn3TK40x82LYcK5MM74o7PO38jJtkqkfy
8DdMR81EhH03si8hWZgMCXQsNAt7zRGs/cfDlP5dj4pA+kNKD7DWNjJ9IggW3uWPFSeyJ4l60jou
WhAr6ND/hr6DiCKAHztQsov43xjSPHMg4ULuwDAGMqH0mCa9Z+DCYONk3v1Edd+90384i+FtCBT8
mL9ky+xHh5438VxqZB1w21CFNKX2PXTxF+ef3qqLFTLew0//tlJfvQecqDy+7CVaxRn6psMBLffe
u5oqxDyaVw9Hy/RpYwnJ+0PeFU2MXTFvmUkW9JZw62XPCEQKTIxcNNj9MjWUfqTzkO4kufJeIgJ0
uTyO3WwNbzQ0IkdQUxqZxeDvjgXqclRSO49aDYaJRm0PusyBN4bMD3Y0SJRpFCMZem1eCdDZZmPQ
FoZBo/AGqGLw959NVnGFTnuISng7dHocaiaKS8sWoAjcgkN/7goNBiNE0z1QzFayyn5D0pkQZBHu
Eza8N6m6w1cLMfwhmghc31/3FbAhknhVH2HDdrTdhnlgRn/w0r18ZXPC/kNjMo+idZfqufHr2ujx
MdOGTt87xudOPDyxs0YPqQ3v/hwS8q40dL5TJjBA9yUrnoc3jBtk3YeYrdTxTM/pk04xrMF/AM3z
RlSBkIBWZTsln4PBD5rRjYVV91XxwtnFEE2YQcK93wslU1R2cfDyoh+qUvB/D3Zvm7pnk8hXWY7h
6BACC/1lf8AwKivPcwsZdyZYFeoxP++S/pBrCygpbVcCrSUXBLqvvs0ldXlVQJqUa2lz+Q+jYLIA
7P6+rGHIs9kN5ZIbljD/B4RSWFvT789KSgV3rEI3XGQHe1bA1PDuIdflamQyFGEWzdbdnqDIa9+o
blYgS1bAs2G+c5ludUsbQxpw2c4hM0qq+0MShHGXDhjQFSBDH5yB6SIFG5sp9Vs4IyeUwrwel5pk
FkHKn0rkJf2u4lBkYSd4Nikzu1kA1cR0Jyi9j/aTKL4OQV6gTHOE9AuHJCeGz43DcvIDEdx2VEyq
vddv4cBIGbYgtsZraJcUZRiq2jh9z6kDV7hvfL1R7rQWQiFDJ8OR4VLjhM58IUfK5SAwArVQfvwO
AW4oS32RhMr6ji1oeobwtiNiyS2DuZeESFgk2w039n9Wup7sROQfOUfYkE7mGUg6yPCZlbL9bJce
xGkqnVMGeNTRjt1hOpejJ9ALBIBNj1sfr98aV3sBAk9/AaL9ci3TfJMmjq12Iqeg8Cmr2+FsN48f
cpza9MhSh5rf+DvBmvJ8RhfHIHALVLrUGoaciKfpXwrH1LNz+OQ6lt1b2N7sCJbP39v629BxWct+
HFvU8660Mwuer4SU+jPRjebTqdmp5a/9q4CrhOfHJnc+JYxmByBUqFt0Q1wV3VOIpimdoGiX6zXN
ggw5heegeLXEIY16KYsie6Ti8LgSgSPDZvJM/Gy9Jnv0gBNMo6mJIgt4t2DZ5seZNgESfhTCX3dA
WhKr9/ocQwMhABD97HrDBPMTPPLUk/f2FY5YFHzMM01ObGL4zHsPasbJiKGRQzfWztT4EoE0+U3h
G0U0kdo3xQByQcMfnyhkxAGvgM4uABAhu2TcgtRJJ6J4BUqYaK/7oqrZW70adMz+sf5h1gMrjMpV
hDVjzgHHBKcZgPnPBGFigl4+g4+mAgJXE4KyjMsqZ7MX4W+APbHY1fRNDgZT4uzLau6Gm/8q/hKe
ssuM1s3geIIIqy0moLOEmZnuj5PAYktO3+5kmdW0awIeB0C6/qYdcAk3itMUMSVF4uXQNKoV5TPk
mTFmvrP35sKQezG9UvPp18M+9glwgaBBrgm/TtNTh98X+22BRMYOkzW0004WcCSYRX80lc5qtXxh
mUjvpp/M7jKr/6r8rZCiZZqr/6rRwpRKaYGLvp1op0eHTFYMOUxzT5M6SGYbXDM6DweJr1t3FzDk
DkpXbsJKmgFH9HfpFKmENHoQTE2rl/lAN4wQ1+TygbgyRWXUT4SuITmSWunNdYCpdkJ0PDug0n/u
neE+LnM4A0pbP7LJ4jb43nPk2dq9dMl7jBCUZMF05oAqFVycWlPX5Bf1heDUSngRYDjXpZ526MRw
t2iT0ZmL015Gse/zTOJZ4jnDeiMYoHaQzG+ckoZDMLvQc6P5Qqo88a1YtRH+iT2FhklDWnyb8vq3
xMsByHiKfmck21rB+sOgD8khXzJ11t0pS63oLmk0T6B0e7dRuAMq42ZI6BItpj0SqN4h3cxY+V7W
krRuJEhBRkYjQwrkyrFgirkHZ/iRfzB+zF80Qy5COIMVkEpPDQElyvMCfuydm3Kz8l/6i83chLNl
Ao/ezhfa7TZlExtqA8eVk/Ym3X46R8h9WwNGpWDglTBkjIg/Z7U9x6XX0iSuVJI2mViAQzO4Ni5z
h3wzrzVNo025MdTmfCZcGT6/d/Uhw5ZoZAweMb5EOTwm/VVBfqyHFGGmz4yEtDt+I8M6Ib2JWK86
ENz5cibLZlk6KvBiTSpgLVlAI89DzonBaymTJLpW7R2RpyMELaiSquD1d1hQ23zWAg9Fr2Hf7r5f
gMpkuYJZxjsWcaOx8xTDCnaywqIaaK8u4pV/NkUYnfQY310tOfmHQE0XjIJjF7wqWEsh/ysjtKP3
dytcffyCQzGom7aNcrnj4C+Kt42Soca3iVWS+6krA/Plds7eR5ynfY5IX5XKvcrcsiccrkd3CsXY
53dZBKojHmX2Mpi0h8osIYJaapuKdL/VD8GmVju8FzNwDrYwAtA4dBoEBS5sChmxM4SUSSjPwUGv
kCoNN/TK1fsyoyRL+r+bt8FhlN8Uq0mEhR6+JppJ7UXfZghQhCrKUuNKVEVLQCXM1LtpzHaIn4fr
ag1+Am4fkG4JIRLYDV/i7kiDN0NxjqiZGucts0jSj4lvQomb4KsC8dxqlfBsfT4nJSgu+E9FZ/tB
0EXEyMK/tgqEEChnPzVEiRJ4KEYG5zon1pDY3xVk19Yu11N+s0Qm5SkGF1fOXqJNzuTdGpIhmkit
mJp9pKbgdGn3a0xb/yM8rm+mrKOYvJ7xcELn5MVuFzOLSmsexb4xRvwMxNFeOD6tigBSH3RyqFoQ
LKPzX73CLQeQZiAJSIbaKyHPIzYvUVdgjN7jOlhyaKp+rC2F1oOB6oDYsBKn8VmPDgzj0Ba2LNPg
1VMo07+kxGlLVs9LdWHSHpqiHG39LoCmxhXEA0Q/78cHBC4/ZmJvPOdrPcYzsNcr+lOgwJapmae1
U6B8l1Zke0dA5X8eZMqx1WwJ2mi24GR0UWsa0hlX9EBZzHecnMNiWXyqJGEwjYw0fqxf5PWWfxSM
nvTqw6xZlgh5RvhPWfKuiA+BrPLBlPt1eyMJ+TJ0llBcaGGlFpBy5f+ciymUVmlJU6lt9eoYRuIZ
t1qPDkfyT4EjQVB01C0m2IcVrTUqQpxgfN6oZkL7Lz4Dzj59Mk0ka0A8opkI/zfr9DI4LHbZLFuk
Y1aARgGaopTXf/5Ilkihs37z7tvHksuIZYfUzDqtJnDGs/Q8BlHRAASu2T0GiUIuYK2UpmLV53TD
nY9RGr4ueOPeXeBR+oZ4kX2ERkuTgVfHLsHPfedFicRoUACZ2V9H4oBfSUSLqMKX/1FcHdE2vXLU
tMNTUcWsDQIcfsBzvZJq2qee1nVzII5oi2deOGJpiu0X3wZ9gmE7PB9v+A+q9u8DH8oIObZ7rhCt
8gjbBbE54buctRUA38XxAjB0mAR8H72PTB/N4vEZsF25q39SYkpBRe96wICmPnmKhrDBhelvIJDX
S9nUB5dcQLFowJ87HB8BSe8daeU3fSZHicrvRjs/azL1EtFxUarepW3/du5U8q3x6FGXPgTabi2D
jEbdslNLISVEkN2XsLG02Nrr+hKDDtfdaj+xxN8lbM//Z8zdO8bakpPhMLSQXpxWukq7CnFaBGQz
P/iUpvfXfbvJR2GWVGqI4HrVzs0pvcc1eE+iS0WFcbQywvQmmLGMfQiH3qvByXcFn4a9IkSNNoIa
haJbMyhI1MYq6rNQNaJNOtdldKsN77zHXqXFGwAsGpHBtVarooIsUAc0TaSsaOf9GqaNRA0zIe8L
apCaXoJbjE325xZA7ZtiJ5Xz3cEdHnf847201XXfvFt417UxqZSbcshPKAfXUPXUwfeKkj5NxoKo
mW56xEyH80QSKn7ioLlKK0KaFhof9w0DDSKQWvBeXRssG0hTqLlgWV8PZHFs1UXKJSHeoWgTryjI
xjAQg6ZdBu5inrE1aI/EXyiVuB5IM7mwegyqEei2iEtGS46/AYs0g/8X8VZYG5wQUlx76eRN0G0r
HEILHNnlfMYb2OW8RV8JsYey2meqkt57l4ANepywp/cRFb1UOiksH7Blz9MWu8M6QBROQAw3ogd/
n4nzOBe/I18aR4qmip2siVNffhSYBP+0p/4lbY/yn9ZNdu/NzdmbtO33G/wS/mdYzfl5wMAHjIUu
Y52Exm0a3hPV1Swm31E7BDvGBlliDBDR9LAG6SHVDCoelEu6YvXFyvaaN5k40tdclhFRF5UWbBP/
OUqUycAx6qwQC45xpNwMTDlt/EKziC5ONOokNRDwCNboiPz1GnfI971RSsbXJVlGCUWXKANo6WRK
rMR7vNqGw2w/TWhADDZPyWdNiU1ABwndlQcWSnp+kUsqFiZtAm9brMiUP+KKxt9NJP1IaCoPUYTf
HYwdk2YS13WUXdA1wY9lX5ahmKhx7KyA+rZgOIql9bTPQgA7x5rOhO4LfPfPG41k4Z+aGrN4a221
0Y0AgPovgsIpz342dierPoRvn1n4qRGOxDeo42aR9LGs3i40xkvoHsqXmMOClFLLtHMENDZNkTel
Djfx6yMZRDK41mAesb9fo/79dVrhA07OR2Go7O8G72Lsl5J8rGi6KCWeqZcfcrhSiL6bQYb2Ir7X
SgcCe+9C/G78nb5DEfnn42d/lb2dd8gyP9ILPS3tyEj6ub8DnBE+ipaZdk+OQVFqDcVSrVsy28Af
ioItJRM0Y13PFyjDNjiUrtYLFBf08FcGj01hxAimbF7v+VLFmq9z5aQxafY/f47QB/9D2Z2XqRuY
j34b0m8WAeh4nE7Y2uzjcaS6W0oC9dHniYDPXuAQlRRQJHatoSZKmd/YLDesSmpOT0M6OJAeKmei
LVT85YHlQHa9Iba/xbjib7/Q0JL5gjqTpAuCltTTdArB+lUo4LbT9cqF56HmUHKf4em6lWwjzOuu
mwppBhDtx9q7PmXJ/1pzvvw0d0/2UFp2iI8Qbx9VOd6fQj0mwCmhJz6MuPCdIZFd2GSFaF9h3//n
yRoIVvKdPQ0XnHmPRx6rRNxCf2YlUKuoRkn20z7PUM2EYlgTEKW2coKwEBELOhp+PpsXwu2vzwXH
X14Fl+Vv06KBDiZ1UVKpNBUSeBHwP4Dm6IjKP8KlFlBLjSqaZqQsAWHjmHUUdmKXc0MwuYHGgk+N
OHXPvuED4uxs7H7wPeOFmCLgynKaGF09HNzuqOUKgLepEw7CljUOOrCPn2v84jqNZtiCFmcRzT1K
vqfmaWo9qZBrx9NER6JOKTMobEUgj0hwv9YCStZZhbsRzZFGr4/CcmdD8SPxNvru/A2Fof0BBxoE
UhFU2G+i03JvSychwhnqlpe1vz4R+Y4ZmhLcccoG1Qhx/3WR4hQk1CBT74QIgICqB/r6IusCnLri
ztzi84UZx+lJMbsWvlcMKm3yIkdPmfbcmeObi8KP5XiSJB8Iq1yq6YsX7brQrPaTDV1Eecft2FuE
U9ratzgNRKTD6ywdAwJke/UfmbYZCs3BtAuHEfQhFv+88pwqZD6jzjVCSQkmn5wZipQDk38bRHZm
VEsAKQ0FI4Yq7XaIhE0ScztxIzcwzqllWPPzdMQN+NFsuGtBBaNZvkfqVsCXPoUI2rVm3XuxAFvL
PkuhBt4TUSPiaIz9NJI6eWkXQfxCmsUeh1j9XuXTOxE4tF1xokBvp44cg6ZFdj+k8GdFfSzobKBJ
tSQZZlbFsRei6wNXGlqHE9zow/hMUOqkR9sF5mdxfqqGdatVp//FwfLrRnbKmOGVi+n4P2aN1SnE
4XW5XoVVZc6cEAH/QS/tmRkYpL752J8V0eG5zlFmJA1N7DQNI/FUuuVrw6F6tHjMQn2lPFY7kRmt
KvIT3yqKUZyyMvcb80Bv20WeHC+nBuIDLYgcAPT7gXsmVuGTWWQWJHCbkGfHmBIO0ElGwP++h46t
yQl/l0RAM0vRrsp1K4dBrlPpJt6ePZiHWXv6okHBigF8pEF+QZOS1df4guCnIZn17xtTAVlGxk14
icSLKRO10A5609uQTXq8SCAgSM93AGekHjh4yBJCXLalEznvWdh6dcds7jaPeZR8J8DOEwpYEEQs
DLBzahO8llnFR2v1Dqi0dop5mljuLRsJcmzo2bN0ifdKotA0h6OiPVCMMiNFEhE9QAWOWECRj8ND
Pt1NXlQV2YC3HAj7JQ6v+L9sqpTetc+KgEzOHh9UIIiM1VXv9cSNSyBGl5H4CI/2RQUh1X/4OjaD
q049C5Cbrh5gDuf0Evj/ffR9trGz4ABMe6vJE+U0k+hbsVgC06v1D6yvrOqIl3cic80XwyGYyrxJ
C3RFKPSLiMNV1XAudqVvcvvCzjLvV9fKAoyrlN4bmhPxvoEjywfFotmcnEXU+M8mtdB8r2UFvtPS
b7I6FFWT4i8cMBpoGze0F8hD4MtEeZ1mQ3TlXHNW8+b4lEbJik4DHMR9ILBUICTTOs6T9caCH57r
xOnyvHNZIG2vDk/0zQL/eqxfijJv69qz9XWVr2JCQN0RwW0YZ3SwmfZGpDhRc9JyUe88VF6i8uvk
Ql5xaYJfjLr05A14f+2lQSU40pMpDmB3xrR1DkJvzqhmEgT1WAmaodJqIihShe+sot7Degs9EuRK
XDNxiGR/iKWeVmx5NyWCg/O5jhgNKUw2S2f69B7AWOyWwCKm0pDanudKbyyf0mHgxzttsSsRPTz1
fLdJ86zamcszQFxBLegNYar12KcjOMXMRGzZCOacr68c/afGVYz9Ew6N7IfuCALYS0RxCIVtz9hP
0wJx9aiE4Vi3qPNBxOhqE5vHL4X8CP2XmjJ0d+wHlMC2H+KUvdbYd0J2GnHDoEoi1DUMF0ipg5YG
ubS0WPqKA7S+GcQdQ3ZkvJ7EnBDz/GA/pMN3yvudajRxG7A9RuY8N8VQIwieOREtfmhROYAIcRGb
Xzt2jcp9EKs3gXAGHkaHTdazg7KSe/Wz8K277qmkZXA6XCzweiU3B8R7i2fi+s7hilvaZamF71Hb
L9veOu/pMtRXnqyWwWi8IDkHVpQCwYkBgpFqZPC8jQ+CAlPxHe/1Vn2Q7aYccZvWPqBcdw1rCZSc
iEX2CMA+TZTdFQ2RUzspsyCR1/nQQpOLteRI6MFr8MIgrqJgELSJV7JjZ/BjmZswFtsb5VW3OBl+
HNJTplCAiWt0ocjKzwaCfjoICmGqtSZxWPRioIeNGZ6SyDk9oDKxStwhgIEC+4YzRsc1nrmsTdDa
nRhsjpr5iyb3VsRAZg8CJbxO2qHOUVfeYUWel6BV0g9rIEmMBrjlbhvss/40MJK8xHePtsIi8b4Y
1NVP4KD1bKUYFcWImUDUM+M7QZ8PWdmJPUkTTz5OcNhOjYIv+RhaFM5tehbnlm9yYjK4A2dP5+B9
iUGRZHQuRX7aFwEHbTBfNfdjS2QLISSn4P6aAXUuLTuTdS9HJDlJNx7RueOytWG7RJl0x7+yc5cg
sKUbWJCK6MqUF+htO4kwtqqZu9dbxQCXY6suSVTjhiMOSKU/kUTvoSgue1ooRkZKkcxFYcmZbbZB
pEAK8+g6iGB8Me+0v/08fykdoQS8wXc1HB9OmHbY0LUoQ/ujijbwfoBoxdu5Oe3k9X2hmqIMbYSO
G+GkGJq/GoL5LFD7Tx24/yUt4qShUxi4AXpF52nvQwi0BRrX8XtFdczMDMiYknfHyAcS1grAE8OP
6imnifRVPuDNAi4lbfjqbTdqPGdiTnyuojpBpy518b5gECbj/jEyNEC4kEzDCwvRz5Yq0sgmFXC0
zY2615wg2JznHPOju/ETnXFRKACd2p9x9aZJ7aXQR3I96ht6XgbmJ/yXG/ADveLe9dwWgtmrNx0J
wtBFZY+WFTo+Ys1oJrneu6gOMTR72D7/uq1XjH7qABSvjzLkIo9qzLXfzWaJERnt/BUoAvkMFp4X
PH99UG1959i2Xxhl99X7rZLliH3ZKl4NNXyf+XAqxTnvVusEsR890jfbe1i1MMtpVCEwZJje/V7z
gn7xNloF7svq9A7sPtW5EZCycWM8XtJZt1q9c8weZi91kirZpcjYQcU5yj+8Xrh1yBegkXFxLwxd
SxQ3Z1FUtRQO4+reyaaMaedmzqN4f2ZOol7BoHJ6PiPzhZ4zKfgdpB/a/XM81dqAZQRHhwUq/CQb
9IfggICma91oJbHi0yQr5sMMs7rPXE8VCQtT1HBawJdiiQDPHZx2JBicd0oyaYRvMVXC4dqhkea9
WGVMD0+jmshgux98fZ0WjRXA8CF6zD2Ra4yCLRuT3/Kv1eztKbV2ZAtFIt5eaFuiM8iS0AMKBefi
y123O5qRbzBDyP65wme5p3KzUC4awrPb2lx8rH/+U62wJjHS/3ilAhSv3dleswDzLMqhSptOx58H
LRSpJek8OgL7p+IrJ1P0a4Nu4Nm0A0Px2JiGzglNIoQ/KH4emqlUkP7eg7WECGtQQjfF7EljiU0K
V7JLlGJmEpLQYSU9+s3lOW0DwB+rgtxlG8LkNJ8nHSd4V6NvuBQjOGWFe8dgXE1DJhRIrzHlN89K
0b9Eh4Td9nipBZ5+8oX8hMbsyMlQFBBwId/TU6QqFz66hvi5vp4WrbYpMq7flRl7NF5RMYhKuFjy
zqmnL/DTKadwNpUYeK6Jg95zaR++EcyA5Qa5GkaSAw+WccyDmlXf3I3TZO0s6nweOTozGwiQgy63
rKKeK/6Dr6MC5zNsz9uq31Bpfs1DFYbo0SPtZE8DRgzU/poBM6uubZlZOEMulvBlbRA/fjL7X4EE
RIEXV4Pai5kuRx++fifhORLUmEgYrbVq1MafI38VsXZVqpOZZJ6Z7zLM+qDOU8WoQfbGE5Er7zKg
INdlBz9nan+wjbWuknG3qITJ6SQ4ZCFKO3mHOAqApFSYmVNKIpYH0K28XFSL1sCwzOWE9he8tAWx
1LTcCJ9eQwA5VmOjiJ3Jx1wZ+H8715MElMyXLSRf5tmtBAoGzLLc9ZktTYfyu0izg7mRFpjc0KL1
oTOnuq5umeALigxxoJK7FHD2SNyrSX+CPsD/bOXfRWxegvEAsqs1eDnlPwRysikvERW9BLiK6aZt
JGoKtFFC4FUQ3R4UiCXaRCE3+1H2dEveOL8PwT89SNmbAUPVJGnU5guR20K6y9lyWav10PzCzI3D
UBS6+lSsg3bv5pmC0J077vAz5/oWZ+4zErzoSE5/tIQ0VWEfeVhFstTIsKHb6TnpKdXc5++eVxuf
b5qNvpAiBU08sui6PfKcY2qhBE1TGJmiCrZKA2ywR3aE+tJj79eKQtx6uJaik8gcAYLBqWw1JgE4
m62boSE6X8tsLe3ivRAo+nDi5XJz8gn/d5zj5PhNSLkEPxWOmXanG9rR2QSDdylCvX4IaM0waE51
VcmTJyCuimq3q7ZPEqOKOBrtqXHVOqCGNmnDZp4yWK+JQ6YuHujlje+59oFi6W4i4zqD9XEUG75F
qO9iSVp3RGYjt3A9TNkOKeSXZbYvOqspmoUfJrlGva/DtXMjcFv1FsGM63RJzVSKiLa+oXO1Xkzh
ZcqrQ/JdOiDXkXnHWMUpyEDLQ/g1MPeF+TGxkC71X8el24HwdBN1NJZjRmNdTcgvIwTUlERSVMNG
hPFGzja5weT6H5xZcYArVc43CLkG6vj1wWuvYHLOFhjuqudkEjWBbAuoXuCCewWobZLgC90EMCMp
g7IM6jcT/MTB3+nwuXD2ZOuehOCrQv+bpjU3b+QGV37adBI4/xzRoJq9gaNhhloD4xuIZqmHC9qH
c7dOl1EHyiWE5q9fprslUZmvUhdccHoXnqb4gEQY2qtGYV3Xd5+gRp+dA2FE1asPf4nsj/PJztVb
il7s8NFYT70Rk7qMYtThghGORduqPxhRRStVm8Ai5mu+JR0CLN/tkPng+fMmS1JjVdPu7TYJq52V
eRR/BR6yugAKahcviwNeglpe3qZxahuxaDS/Efz+xb1mqXYfTPmDdKLwSo+eNjuOrQCnw54fTtuk
Hox9VO90C8sahx+2HliNNaFU+6eITgiQNoySZd1heKNSqCNk8ARAXLt/xJw5VR+ym1H4OBAsaf9t
+gVFY0oCm4ZXAPGjGea6FR1DaD9BKd5xIsrhHy9Qo41W5Z2rXV+6XUzFw+j5+ABt15ZEtfbcpLLs
uBkXulbZkGLPUj2kA0AC9gWXDWaCuWYxm+6Nlqa9cZExzm/AAZkTx/S49yxfZmyzGGzusf8MC1AX
gFOoVljaS1VexgjmiE6wB3CXVoQxIdM3GwNwagkWak2TaueRybRt6uR5+yq6EoJ6stk5KoiUxcn+
K1RT7bZPOp4N1A+zMPwlpPs2ULXm0IwqDJuHrLFfZpbPemmLARimPkHun+pH+0Vutv6bzRxWYfz0
deDdu0VtlqcJR7SrOEStwv6KVBDtkkChtkY/KZYPS/OVXmrgg4DorPmnRQ2i188vBKB8zKxYTv8P
yejCfn8gvhpmgkMsIdiGQAdrFrba7R9e2axn+iqoTV0jn6zGOvqZ1H7d6v8gWxJeLAWvsGB9Yq6H
odD9bXlqdDxkz+KqtcQD9ombAI3CCXOsj9q7kFifEA+qxx49ovytp0FJifS+B3itaXeEdXNG2v5y
R/dKQubDeOF1qOSuSVxYUk/25AH+5FgRykLy2ggUQ73W72PbnM7qodu43z1O2X8xrRmgAwTU6gK5
0iGyunlF1QOyXK9LpwTgXV6crAD/tk0eS1Ec1mjafjAN+lskdxblvTdWze+urhAURXcL2kOblN3s
vbqJtZ5dEhmgZwHl9DLLFa9wtGxUaPvNYm6l23Y2p93hzqUSm6/Jjx5gvOegd9XVZ2KjKRY0eVbB
iRDssB+G2FusBqATFqzoEoezU1vBAgJlQ5Xpf4YM8IWcnhA42sO65u4J3jZtNZifMKbrNNXwvppd
7459GJ0v/ovaMf7bUYP1Hh03yKMckPymMhfKMG9/M3d0QGowxsy1UNeIXXSIdGEh+qY55q7Ht3Z0
JG6K8kKSFZb4aJYumpwJUYMgvE1u+5r16KCJ+sC62BeDZgvyeAOfYt5slGifExyauJVCq+enpPBb
gh11evCiZztEjR/PT8fucnqPvIFsEptanR0blQrHbqYuATLpKVWtmg0zRZ1RoFxW/IGtGV6laZAY
eyvRK/bJYeOd2zqxc6Aa+14UnalkieqotYALnlr6RFUC9XAPjVriJOcfYLHt5pe7WzfD4gezuZe/
29uagw3NO+BP+Y7xgbbdkXIt2958tBJFwyj4ufahfgTyeWb5RViDhzUx0MHDh6qDkBW10nVViqa2
yb8N/D/ufFvVZclssvvhn9Ydmg3XYwPwbWsizsadFkVcHqNjqFenP0QaUeXBKMwauHOUHUcjsyiS
W+q4Kj1JGA/1VZcI8eKhQhZBstcOZrkE2JVrnUeVGFD2Gs0+sGrnNgf4AMucHDTeYk/cZJWasSTD
t0yD8XUUVRVczMNbhsWHHOIfKvHY6kNXVy7IrybsJQNVwjWKHN5vA6Gm4NjhZw8y3311M/uVOvjd
T0xZhZzL/9o/lPNtYx3aO4nj0eTxWZNlZcuN3W8zvkqfCiLkhX//DjnBApm6LN9aIvUpK11nKYkz
K7B5tLqW1KCkxoBBO8yJpijTvVcjVtavyA9Dfkq6mEgiPpLXKqJk6QPP30k2i6dyd9/IMWC947tm
hdMAnDj9XlcqtPtXxm44WeJVeLlonCH/XVXXph3Qo/SkiiLxNxuanZJHTdy6M7uJYJx+MdUut/KJ
oENzGFT1MFnbrn/mITPYsKFpgJLMqlEKNotObOK3jVGJ7ipjecw9oL/m3O0GXrRIBvj5NSRse7AT
OGIz038cGq5Lgsl4wfudW4l3f0N2eZwMCWxBKbsmXgBilf0MiZ5xnTjReOTriyN4gmpcR0qtsE/L
jhGWnMh1xsMXOWo5ig+eNaKwlTXHIhSVtkkh/KknWj6qEHpmIKpWWTE+8HKgqzYEJ17XwBx2dQ7h
C8hQJHXgGAqagzJ5oIZ7BNOsfvkzR1TfnZHnowTI+TOsmZtFCU05GjhS/Z6ke/jiQgthYdbhuEui
v63+GuJbWgKIAqcO2SnBMBILC+BTybAX1iVZnlqw2KJQq2q0lHN/J2rFHo1OgqKN5i08owtxEQQR
n1gnJnOVEsqa2RA4prsTeyxL3hDOq8yznaR8I2Njc+oqdvBFhph2Ggtrfyr3hyts4rOeN7TdLvJt
13cDL6PlmI/Kp3cQ+OdVgxE8LL5EYt21VhDpyHR3RHxPxB3FMHZzSKHfzICgtix7YhC1mcbhVmyc
rakvAvprjQrWUGEeEPEvBQzb8q661ZiBOYzRD4a62nGbFkvTXBo4DiMW0LersPlSaCiVcHd2kzdz
zyf9sMx3eIcoAk8zWrXH9TQOpXvvsGGjKVgfk64LFrrH+KLq+1BHHWHh6EymtTM2BCVPCsmtiaoc
SUbzZkS/GwZwk5iD5pOqMYhiwA6S88NxfZh7OF/tGfgaiwPYHPCzC+FSsAw4R6+QIl+Ly8gCEOsP
p+JduQTieuqHfK2pxDl3v6MVs/W/PY9VxKOueqO+mj9ff4taKq0hdr4bZMIDRlVYZDHt575T6SdD
buoJnefMuzfe29R5t9DJcOAgVdDfhb4oAwINnmKOBUracxn+vQNnrVHInDJhNYqW0qYfvkL01GHC
UHgTKNPtMiyXhuaOwMm0kOaQFkRIfK/lmsNKQ7rg6u+Apppg5Jm5NyxmyIVMmCFVgaWhtFpjNuvm
31GmIdC3H6vrRnn5cLK1Y/TnhBdjuAwL+9UqOnvDYLjSvJXZf0qVPVr6EL5BNEWvxVrheqAUtnqU
AqtqRlCYecnyiaZE5Ky5cSGRDqjZP2TYHYuEOqseGyk4Re/lujjbQHvDh7S0REllkQEmdz+JYOip
sgtzvX3I8tq5MRKI136JnZeF2ugL58iYgDV2tZA9XfagC2db380mr1hWr+k9xwsFQ+hZHUPVLio4
D99uMg57pFr9EtScnHu3cFFAhrepBhf6vF/j36HJtvIq21AQo+JiP6SAUXpliz39Mv/vV1p8GNJk
L+VzbzWXioq3x2WBubIIzgt7GNpOzz1CQSzyJt3nTtMlmJiqOVUZNCmGmo3ZXCnGtpTSBk3W7jqj
0NH1sEpZ/VMBGxi+RRYivr85M6zcJCSOCzlCtqm7t0fAvBVmMibYY7QWrOajG5MuUKFCLZgVLuo8
IBgRscNJRVYGnW72gxcNqE1WHO0WzzaJQdX2Hx/P/Rj5b0N1O4immMDxdK++OOgOn8EaDtwMAmXP
3oD9viOZgo4rZzkE6vA90FRXKJ8p5TJqwH4Sxj9NXeBwE2x2446pVni6IT7ZbC8Q51JSGtaTzhx+
y4vXmSzQPhTl9jhUsbBRKhkqJD9PHn6E3uwuMo4Ovub3SIzRx6xgbBlKUEwilsyJvotXZ80JmbhB
PcOVDClyrbXzv2H/TbcDS1WofDtFc/GSvkUy76fhajj+XJHl9/wJncQ2uh4fBPVTJALaxiTlll8A
Ydm5l3ostKGfKPciiDQvrZAPw9GjgV4H2HLzJy9dwR5aMk89prc7999ohk3LwBDkuEGGV0RwtbZB
/rkyekRVGU82AHDyzo7ZkwUpcKhu2IH4O9DWKTZxaY9O1YqAeEcXolVt+hzWcE59BTSwIboNcomi
vO6mOzA46HQPJcMbXILRdSicvwxALsFwervE8NrE825Ll4PN+7TNPyv4xGwawfnwcHif+D2jEeN/
J/6c5Fdj1JgLDc1CfeZMc6QQxwhYf+CSRxfERDwQod8qXhyUWwUWjsAlPQE6tHPwg4gy5SIsogRq
0EcfFG0BBdGUDmtxiqbfft+eMOqivEah+QVhjN0y5x0d/EQbiJvoM7X/AijNtfNgx4R3BcQ3eUn7
EOIO/NrzBWsDCXcb5fjTgMuKPVUU/s6PLH3cF6NgHW33JrEO5B3EOhEFnuoajLp8kofOoEZ8twFT
4V1YzSlQumsGqzD/Cdf9zRnhkQaDOfNNbQGgcZCgtYEqHmbg4qWca7Vb8UwK+xPV4AJVHGLpTwuL
Emt1VeV+Vwt2IKvdmcAl4J4RP3t2wCQG3t40MqmhHQwMPloP5ulfzKpWS5kgaRVbtsnK30fnda9H
fchXgm2qDVyHeq0T8Vn9YDnR/cYZDNvW8r+XWuQjGxpNV7ZGIRExBZ5Fx7VHp4fqDWzZuH8WXH8y
CsIrGHYQpbRE/pYFaBAMFvUFIyFhybPX4XYgv2ygf537GiB9zxP8xN2kX88fZlYgpWiaI4Xm0p0h
HvQh8sJ/VWAJDploNl3f2jWfVJBuaKZ1brRkB14zradGo6+F1ddPisb1D5pb3KHUwa1pSpakiT+K
6enX4vHENlKTqp96JkuV/ya99zpsTFoH3rE+FNINMyRiSQ2Bujt0RcSCKXcbDDwrkBSD7bL/P19S
hhXxQEGQeC2w7E3HoTVWDPxqHANoMfIICdCse6p4otCS6r9y86t8umUEBYnOy0G39r1aE3asqb2a
ePnn7uvKe5u+zXABiZQ4yW1xR2Rt1wy9KlwNjrard3Lb+aAeSNa/3a1/krjfWz0/oif/1ENMkApa
tJOJA60PlBl9QaqKWl2GDWozcKW4WDKCts0ZdSFH7E8zKH9ruZ0wWq9/h34d+ow3/aBIBCzWvkWx
LgfugS99eoiugd8f5V+gSmjiPr9zsBE5pcMwRiNjtVJD64hsDxa/az5TjY0SVutRUkfSpP3AodgB
MTW84K7kLLwoFKajgQmvz/hlaZ3nByzDarAYarcln7y0LOkbCJaMEYR0haE0uYUe230BC7I0I1To
kF5NBnCZmWjPxLJMAkNQI9Bz5JKMWX2roEcHUHOC73Rt4FY3/aBNtkU+8P9iwA2pV7b/OcfSL1HT
sEj0jGIzZSdwie2AqkDzQkm+H474VgcMagJs/0cJrbqjJbX4Xdm1FT/f8M+RQt8UVBbilZPiu8+b
/UNe6JFwvveMOT1qFFpz8ha6LkhPVt0FGnV17PxLPxIL7VrbFlDqTj+DffsOISHuiuJZXQcJ98cZ
WjCKn02SlCdYQlC8TTiWytXzvqO9VuoGyCAtm0SSmj3/AcwoCc/68UyQpQJo2YPIcAkU899MJvqb
CZUHhPq6EQn8yRAMycYCd7ApZ+KtHib+lOiM/9c+L15l+hIkKkX8sLoCVOaeNUpdKD4jXBvelJdl
6Lix3RtnswicR+z6MdNJcCYGN08PXMhkCllnS+5A8pP520XGJKCsrdeI2R5Vipfho+ZUakEd4HlR
rermss0AOPlyNM2u3SFNFILNTlytWWNPbQ1SPqUW1dEgy+Y5tS5yWn77Dj6X8vF9v6w+D2hdIwcc
NGoo1QoustAZFa7AUll3Cc8PbVzBWHnjMJHMCnclHYidTkoBVppKrga8URP//JIiIdCjeahN0OhV
eKwod7rqHFq6M5f3m1IM1D7QBehi79s3ue3EdYx5kUi3wkFOaQJGWysEE/bklTCU5WuasSegLDvk
QHVbbDSuOQhgzLYlfY9+MG/UUQwqTMd/6+ohSjAOlWouDYcAB1VhRvEOWaxMnXgd7ZhwomorJrnJ
SCOLONrzNBqj47gfwILx0nJ0Pf7rBWsrxHs+ccCiifldtPpG4zYhNDZjYFHBrdxPrGwVx4Q9lvN1
QEFkWOwb3PkcrrNiTsPmTIM+h8AIdoEKi+9hca9oCxlslwCAH9CLqCLhna86OzA47XlU4OpOur8+
B2XJXCZxxxCBSTe9zEAXebXlRsUUqnVh5FyIW5YjfD7iGmMD5elj3vyVRe8e5ucJjGNDVBasCaXu
ePAX0YTP+IJ2FRAR7mc0M68gzjGrDrpA0foGw7GJuls2nXA3ZUScD513edT/AsN6HB2rkC+ciVqo
WCAD3YyT82vYrZzeRTaH9+8FGb40GBHFT3QmMDqbnnRfEfLvRbjOIOxIrEDQf5KQtAI+EgGD14Ct
ZvAG5NFM/0cFeIo6XF91qPJQ7zH+LuGfYC6R9i3Aj0LJij+jf9OwxaHx1cmOk0A7lir36LanL3jc
/Y1v8F1lP7eZP2OB6sMP338mVzvQcAXHJ0Od64idxy1etD5+9DG/GDrJQ0SEtaJJHp1VNXVyaD5S
9bNDmQrBSSnrn4wC4Vk16uS32lkeF8tjeOO31mr+QWvbzBEVG5vm3ODuHQhAKcRQ/ZiYgMHRtViQ
9f9RlrK8EjZeVHnKvRTtEcMfEuZHzeRU3/i/zjP4OTIVBDCrTBTDomcJgif28SyoXX0uqXPstwMu
QAXRk8iE0iYdsqoT6qTR2KoD8wbizFm1l6IF5+8s7GjyZy5SAZAUEJkwBukVx1dX3PT3yPq21If4
EAYSmz9iRdb/TOsaRrJxmbSa3gF+eC/1u+Kbt89C4kspdS6d4Vnv8j3GcV4VxAysXOaqain4e8Kw
gRr01xW8BewzuQdWkAvflfMK2NJK0LUg+x4qhgykWRJ5hoFWQXKJdi0JmcVcyYx5jlk1vyG/2Nvq
RjFP3R8cPX3OuiL9JeNobMH0Jks5dg3X5VBkaL3gxc7QAWfMMoeY7Tf9f0gSLARx8XuIl0am/RyI
LfOxaAoiSwYrHHQ4wuZNxytm9/XvTZ9cDtRgrts44qEGeKzYGy62LHxBYa8w1Q+7Gy8aPQqREy9f
TA89p4X9m4zcYa1CSUjjekgaq+amxMjW/+gISJOXRJmPk7WMzRbvANl299KJ2klktm7Zm0ikPqpo
PHx5m20vuFTIVJYbuD6SODc1yAoBo+/mX256XgNRSgATG9sNKCKkxA/95q0ykB7fSZMqV9UVc10Z
wiATQOffej7eYhQceGOrivzwbEjve0ipSAe2OEItctGQ6sHsdg7mElp+GBzwrXnDgc8vzAMEkwbb
Z0MfggLEZepknGs86fOKclMb+CNi/OYeKYKD4sj9BunNmUr3ug0PAVdBWuf7eo0C8y4SWULb2MPv
KO46hSq2l0Ndot+4HLHwhWynogdVo+9tmELMBEZPSgpeyDPzrJ3a7SZirNm75Q7K7mcuS9vEaMej
cQkNDGwQnFGcTcj5y7wL2sS7IqTqAnZmKBQMXcvjyf1fBft1fp5kh/AVtGQ4dVRA/bA4OaRYUVRo
pH17HmnB9N4JRzckr0gVomnVQZAStKr5t4ANTSpDTbtzFU2kIYVb4kGJ1a79ssMOafpm+MsGs7L4
JBVaEVOjbOjnzyk9y1I7CpDOhz/M85m/h0P4L0+uLXg+2qtvmR51xeH2Rm0asA2kXlcsvcMgR8rq
aln6Zo+BCqnQefcFrnqtiJSB7tlFF0WXkD7zQw7IOd3ttGhuyo7bQ44L9WlghwCkhyH/vXtJ+cak
QltfEHYi0KfPoObKg23Ah7XCZiMMzMeB0RzOOCadvaxZzS7gjLub/2seaGAw4z9sfhPNpdV5/tJ2
nTEs7ikHDjwMMuuIz9Z5C0g8xbHwW+MZsn1W4UW8lsbZr0e/13HezJrrCOysMCLTBI3TH824aYIY
UsdYWZ1qI+RP42fWfbit5oBaBpiumD6PiR63Bb4a6mvaioOvmcMdbOMyQM6P7tjr+puAtA6+aR3K
wubs/O06QERFMdISRwrSL/eDuHyAhSoyHAK7M6P7JvtfnxkTmIWJdRudktyybz270cawT5KTe9Cz
KLLMMfPj2DkNGsOmAz5HIWHJ/fUXIlqTfxeeJX0d9vjyQ7aYtYKzE4JR8ELsr2IwY3vH5A9bN3Sk
DYXDhQwDgUBtfYQQMnsX4hJs5JXcR0Pnr7Q7igSC+82k2bMJiX6IbkBIPZwpxH99rzu7k0QyneRR
I1Qa0f+RhZzO0ZGdAVOaHhhCxxKulyy6/46RnMYHTlrVMWBEShUAYwCCaxzVqQqkS5tBXQfazc7n
jYVaE5sXI6zdPWNIKNS2KWnBX9klEbY++wWR5WuvHz5pDzqyOnqWKdnBlsIOx9giRHKQ4wAqfe8t
CZbbiecslaL9D5EjrKHuAc5aMIRTFfvRzDluHIvDCDsRvYiq+UPXF2/50I3mZlLA4H6stRCGcUEM
e+v6ZMtOv2om/qkZpEOZ7cNkPHrRny/ygfmeJ1tiDVLXIUA4slpJntB+vwsabAdYgTXvZ9qCfake
/XCXdSD1OqS/kEyYoMAtnjSbs5VnjteUxGSTVGEETHb5kxe7Zubmhi7aodWnm3HTef+iksrwrBQT
T7xIv9NHPQy6jGCi9+Vn6gfeAb78JITLEc8iTWehN3/KZzyGyAtlbvsOqcad54d+etQOIMSNcn5R
B1r+N07JcUOxVqnrM56VtM4zD+pJW23vcKPU5+EZyE5UtFJa9eoQ/AFZ+1B8sm1/m/3Ya1/1FeXy
BT4Mn/oYQPFSL32PdeQZxTORjV/AaxVeRFWKGhda2HM1yZb65Ui0r6sSRB14Wr7mNnbUJp+iGeoI
X80t6rDju91LfQSDrdzI5cBjBuaAKJgkR/cwNGYn0VE4TI+ld4P1tFHpLITAbcLyOzw5OOAJNbWM
TgI4sLCkMLNw35WxHaCEyH/5nfZLGL5cHJrkW2ChUXmugedIJz2ChnRCI0LqxuojzYgYHPz1rTTb
D/fpjop6cip3Lr4uCYg52bQvbvNRCzX1al29OXgpvsJ39qwZzoNFI8WchcrZYofVfREKvVzbucHb
sLHjX5fzMlvOjQoSvW9VSygIA0+sV5cYTUUkbWbfubb3UzS5MrWXKcGKLZNTn8oeu2Jb4lRE38RI
G1rOlipjRDEPQqhR4lnrPXAax1XPfX/Ky2t1zINpCIRcyuxPqhBowfvuqeWSEn0TnN30bfwypY9f
qX5hIF0uwaiFYpoyXjsLua7B0AhCbJ4+cLtmwmL1zErhqC2COm0N/WlXrIHtcJNsH3RPju9tTndP
TBR4KpRpnVMJ4DLmEwxNkvOsf1GUprI2gYYiVZ0I6RA4/ak3Leidxj8GcBf/GRSE5ouzxo1MaHEu
xh5se2sRUf9yxx036+HUIYAJ6I4bO3L4x2LUU2LAeDUWiJyyV3brrFPUZ43AUp1lWQNtquLVsr4P
gV0gIfhfKAgBTyTXL7ABAMA/BDpzXUsq8eHY2twfJZGMdjb3yqtvyrOPZ3eL9ygR4x0bhH2WAveN
Kll2NSbHDWYpKV6xAMNYxs6GO7ztE8KCK6UgII3yPkNhOox3t7ThyZJMoRDuAW8tAnJ6pvGy5TTq
GN3A7I2LLqIr20MVOr0S2NNDOzplZWY0rQRYQKVFzUkiQ+ZpCjoFeZecn7XsUA1kNnQ7Dv66fqJu
WqK+29v64/CIvow+2oMW0mB8T4yJxRd3OLpS/O57cXhIKbB+XuotvohdQsvN3urrtarnkEEQRWwH
IC8wmbyAyR10oE9egeYKsawduwhUBOyX4qVwLG7uFw1u0uozlxo/LbcJdEYdbaYIy0Bbn/TQ0ptH
mG/cA8ckfzS5fJtQ7VkEmUCINC+GeKObqLYzXr1QwIxxNZtBlbfofV+WlX+ly6m/bZuic2hhpr6O
b2Ol6mN6OfuUnMrEwGNDyA3VlvPAnK8EsTCNKj0UNYmEORiwYld9KqePKTYjmvtxTzXVmiozu3hg
aeUkteTRVXhrrtmYtftAddZ5qJ5Jt/GRZ2VkGMMRfuf5f5zG+K4lDvQq6JMmvoYbASGzh8GnA7rk
1Djm/RZdGlF2Yk4z29sENE8EIF2VphUcBn1XL5+pPl2jH6uIY0lwHN+gMamJBfSWPs/1uGFIDsp2
s88fhn+dAuemVerurQh4EUspDo6D3cT3bErur4+keLWFPj6D0x3PC4J48lL6qQtzaD63bF3z4/iM
o+OtG2cAMnTkC2nn6PNahHJ1SKXs30SPLbOg7IsZB2M1FDrl4c2ZAkdJhlOgRi0Us9ozGUTy+PS1
7ThLMdsFORJVKW2xhCL44jAx8J0/PX9TrymU5gU6cZg9T5X7mwp027JIS9oyV4A5g1RPAZoyJQWs
fAIqngZU0sL/m4t1MJU76Mx3X32kAgUHEK0kHbN2kAhAJ+Y+S3IhQO94aP6GzBLIBBK8WRHyy9FJ
fl4hI0RlsrsIDOUFPibc3e1dP8iKgGkA+ELQpWDiKGnOmaXQn/4u15Yz0dRY6KZgc8Olm1JHVeLH
wrXzqK0XZOHWA9U+DPZoFQKclEa3EupJsxeTMB45klgcj0Lg9Vov1Npdr6V+ZMUO/3BEGtu475Yj
l+Bs9deGZSPYSUFJrpb6ckr13feyPnq8XuvqTUt2OjdSFrcmsgX5WlRMo3MbGqsH+VWqzoZ83Kub
kMdahKRD3ivy/sNbFnEB5EBnCTDI8MqIn4OixD0OiMSN3tF2RaKZ8PnIGjD7SJz0cUXc2Vv1jeXm
UEupFJhP4zd3jBhw2+fpFWt+eNuMMTgRunMjagZt8T5jVwWtwMy8mFAd2ZsBh/TGuvSEXinOKG1/
ycmFE5iQ6GqGgzjiYLnIko1N3XtrD0q4sG8QsfqYUvZScD9kGFnm2RikIUTwbcvr6BEkO0YLX6DJ
4niQXBnqA2YtiLmrxCkNXWIGQUa+s/YYRTBoSCayU3jTYSvUHc1c9E5/olN3JH+xOwQ+nOiZ22t4
V6PkY4Cj6xfJLfeji3qnmMx2ye7/fidjIFxAGS4bAcdFO3V1iPzULHN0mjjwMedcENCuoy/i9tOu
Uxyfw8B5hXerKhzMiI6mfJ2y0COBXhWXG+FpXrDXZE7FhvMsWccxjJf/RERFOtDVq6/W8BWn8y0d
9St2XqQs/eM4GEiqnGqbJZBDeAU4KjvZ63RlJYRs9EfrIcV5dR99vnk8QOsieDLps/rLiIHO2uNp
jErVDenRD9V11WcqO9M2Gr2LJysoT+mzOFvq9zpUmwfMuuajks02ouacmK68ZBAbMlGDg7GTyLCL
fRyTAZQ868UxHwMUPj7l0W2zVcPvavU4F0lgvoqhOHKWEBEyaxJtaiCnr7zPS8lNMSzSJikPvejX
IeekF5JIe8QLdYzpjjVDcjeaK1OzAeA2ebKj0HLpDuc14XSwdG/l3l2w7+PQxv7wEr8Z09MvaVaM
mGNr/1dF8wk2iO9jRuX6WSF2OtnUcxd0cnk6YJiyP7Fy0lDiyPTer3y+0oGsRSxoNv53aOQEOf67
MXAF3BbNoCJtG3M6/IrDueNFteVQ66pUNPdJR4Lh1TH13bMzt+Q7i137zIWFCsH7XN9G2R0iN46/
u6jmEYtQIzkegmOHa+bDip8sIm8KWWPM+hMQf7caHgSQUZewNO6WlH4oU+G9MNuCxATG6d6r67y4
FKY59L28BfoTpSVe+wj0/hGQzI+rn7xFT+vSWkHwRUHa6LiOft463ytFBDDCLVes43V1RyUQYQ5v
7gxGnHw7crfMTA7gCGmNQALJutA+beEADqj43VlUdeWNogV9hlvQ04bM3x0a52ZqEhtnQEuULAYO
GAysMgc6J7nUnsyILn2zBlE20YmMB6B7lSD7ow6vTl6VTlbWLskK/p8XJmFEcwJKtYsPPIlh1D8p
uwP0ojPNYS4g73ST78WjLUP+Fjg0EbpFqCozFQF+6frwF2825A5UNQIeOCK/WwCEBJZTV0zgTwsh
UF/I5BtBssRO3NvEi6mKcMMDpdboGozXANEyhXZo/82FJkC57zNVSQD9msQhtuQEPC7ywaP+s8Ce
UAGy4fsnhuqUGmwGjjAdPIW0BEChAU1B8iNOnnqEZO7fbj0rf+45h9pvB4WyfoKaCLueTAJoeuWt
YLmd4hoGLhZu1lIHJ/eLbDpdYSucepHhKuI6tUbDmLz0U6/lLOJjbO3wZLee3NdvNNDQQ7GIS/sr
3hguClpXAPFGhPj8txjAV+XPObYjfBKYJ0zoUdcttqj31fDADpQoDb5G6bNV2OimoDuX+qtKYqLb
3hdwW177B2hzXTnO4ktLeI6RMDkycsshYald6P0WbPj49EQpdDxn4gRg++lSSTQhtvxYlrYDA8jw
Xmy8+prmL8lO0ZybjsZPZn6eNA2QeeYXylk11CNzdvl6V18vx6SN6fYyjoRB8QPE6DIzA/h3/fvw
tI8Lj87kxhXp56frgfqiPQ4yjBdPhmWtEYCPEg5gj2t/MSBAhLRjpsuqt2wsVqOob43jOMJ0YiwW
u+fgSoWXenAsk78gjKGLKyHx6CkSbvdyQypDgC+ioERWUIrJ2+Cg2SinwkXjsZ2jLADg4vmLlo/V
oFZ8eJiHoCqjFg0dUS5SVj96XBq7ZMkB42QBIiP3W+B2k+8YlQRmRvRzmF13FzSER2gXDxPyUbcZ
EB8WJaeeF8K+4EE8UusBm8788BSP917A/hMDg9V6bspybB75x30MTNQGZlkhTf5roKl36EVJVJFj
Nhbc1dKFDKz00dhtLUxTgAoagF6HSNsunuhIbAhoMk+3OcnbmQVtZT7x3RIbemDRnlPAePeDI0Qj
Xjreb2SQ0tKdi1K9lKBTfDsR6uWL9mvkg+nHPFrl3RNe51wIpuUgFIcb7+yol7+30B1zwQvsRfp3
yKwJ/h4x7v3utguosMlhdLc6KECDGqELFmqtlvU0lQT+h9yELt7YMkTRupChZqnDGDDC1Vgp4cUo
LXNC2q0BLVBjIW5p6hTY7BjLk0h5L66ISk1iTd0IJbqIWIiTuzKqyX9/Ntcll9k2ov4L39bG76J8
cMDELjaYjysGfaOaLsFSElx6tTDMsc2a+IFyggZra1VQ49JkWffyrb5PyhEJ3D3q5viAPufCeTOP
CmGV+AyorFe9bb3sPtvcTF3oI1OHz+Z1z7qcKyIp/W5+pl6ZyyIW8BoqPu5WRYufD33dJaf8R0DZ
Ry1wROx0Ji1naRLNWTKJohadmgUMeWt5xDY4ocTkE4hva1Mp5njKIFlFuc4QI1t/GiYjNyvPwsbp
tUi0oCo3UCwKxlAxn9nEHwrF+qkcgGpMhMCNKbgrpU6koYQlTGNotU4csDzQ7mCePvNAfe6x+9FL
kzjdonP5CWAogXuG2DZdVfSCCI7g1SqHzjyPClWyKVncocVEY2f/T0muiJtyqd1HPcRADOpOPJY9
ljIp9jMXTPvtt+VJTQ1yaKMXSydpznUiCJ9q2nlbqH4SdrOsqB1m0Z1AYFUNrp/sNFzNVqTIP8eq
ToAm+xYg/H+5VPxhoLwIRgaIHjYE7zC8QTpH15W6p2jziOwtx/T1cvhaSq50Ag/oZaLOrWA4jbDO
tve1UghMYr1vyBFMdRJFmw3BhGygYoMCtQqhzcoEnsRXZTjI0jcHb2fVqlci3vl4IhwM10ZEKeA4
jicMTSsKMzYK5yhVVw2oe9BOt2tZv5qIdAYmcltLokp37QkT/V2jhBzcEbaBFShdZ7RdvhWK3p1X
VOc4p4LkVvmjccpQQQGI49X7Lz2GuV2y8S6vyafOwxdSy2SroO3srdcuPX6bxB9Dfc5pmbauNvbF
viW1yPrVUMsbl6pkSK15Ipg75UlXjcvxJbC3qU4rUJJRDhbUvgJJUDCJHenFMBTxNkAWulGx0V/b
urG3BD2s7GOEFySSgubRiA1sHHcmh1fMdwzZ+uNQZWbJ++0gVy4PpatZuZvSEjrmd18GYvvQojgd
2dVoLKuo2zrpQbeHuqg6OdEdGhw/ZSqS+7FLDZnzcYphh1USF7vwMqzSMQntu4GCeXUgSIGlujIU
Mt9HD0yzQTrNzAjySEp4u2PINH4iaZC/C0LVn1hsgyPPk+mcFaOT3ooSTVOlrZYDcBWsuwiUWfVm
OJsxilfJP3Ro6/UyiSl6jXPBM7/w9oB/yaNMNWZQNR6pzqFUPkeJ+GQr2Oz+B+xZgEghzbZNm1en
55sGttR5YS08NVgrDH9ymmEQ5hzu4hiIYwa97O7DV0skIA2tkR4LxzucQaIe/Qqjc9JQ0VAEZn7t
UHSs8tQRlIj52raqVmM0TRsiKHfwVHejia4k190pEhLdrI/XHwUb7HXjenVbscj+i8zf/dbYNilc
TGOl92Dwc24enrbMsHEl6CWINmwjvWtxMFt7Ky1l1R41OFA48yUm49gSwe95jtUh0GS2c/9RoQbS
4TnCCNJrwAa3jABigLejZTWqRFkVF78pLnY2UUc1zfI7fV02Wnu8dylFVMJswFatwqB9ecMEIjKd
acIPxNa01UpBoB4GnXOGW5n3q5j3zlqnIJJDWQgxVHJls1Wn9QgTU9NKtLXfeANYnGhSAorqbuII
a0FEQ3mNwO085BgVUMPTGKiHlEtkJRFNRa+EpwnopA0o9a27WOy2xzclWiUjjCBMssgzdFCXKtmI
LqR0GW2z1l83NOiv397oumcZZSIcIVU+YdB7HckA/i6lmjPGeSbeCaBefC4YCvaSdiGvnobqLMjQ
64U5pnEvkaOwVMYMY74skImClSaPiXb3YP0bYpNaB9hmRAC7U1IbzQvH7mKSjh0q2FRgJiWrzeXo
5BdBpb5iCQDVxUpKLE3pCrat469ZObp+RqAq3tmKcASofU8oMBZ0y/gWbluKAdyTu41WVQCupdpt
TIZ9/K39hp3HH49FBb5O6Vlu7PmNeiYu0c+8hLKUiqP3vye0oYN3d+2rfBUkygT8JKX8+gf+AsT4
/CC9gsJycuPBgxF/3r5XiyXIvMhcc0adwzHiajwItyzWPVs4a/AIKf4BXvmfbXrwo/9fZoNPj0YL
p0FAg2MvNfRw/sRCO2/Y1QKCuisZNcHtdtJcqlrc1ySqZMUIBghFrJefnFTj4o1goHajT8uJYVhD
GdA5GkANw/k/UJUletO2wbpZsayqi/I2146NlfH04ZVz6UGSDXtbnnCR4uDouBoU1XSFiTVWW0yd
b8LCrIJWvqI647Zh4orVLwb+nnGYPI17bHFEBwcB3LMoBL4QJFZFPhUUSdsxbdV43mk9LnxO+H3F
aqquX3Vn1CkizfLBzvRkGuQW4mTuHqRr6vrgCVbvYn7i1c98KhviDxPCWHRbQ/4t+3TiGvpTKucl
H/7v3mDSllNRxieyKafgxL2T8Z7IiGcnV3iVctdZssT+XzIks0te2fZHKaUBPqi5dx+M3qhdB1XJ
QGZ4cZWTcf5YSlBo/Ge5PODCoWetzARm7KA1CT9ykPLmrqqjFfVx3wsRWt6LmrfGjIRxtKfzCBc7
wMYrer1YUp2KQIbSUKcg22A7Xp9c872bSIJ1aUsNhPMI6rylLP+UVy+LOJZC2ilCfqACuP/H1Uv9
7lpVSe9msYLNpRZL213Ol9Na1udTOKFEIrqxr2MmrAaVxouP9uW2GRo59etfzjDJmr7DZkhXmpuz
kG3P3z+QRj4026rUOR4dx9GFXixwTm0y+ajiyqgngDFKZ+oD1qvPgSDp6b/Isx7Boxk3a0Qthr1+
kXfV31pa2oQ6SlI0A8C2umS+liOV1Nh4F+Rv5Q86/NCHRipxIjxdH5ncb5tahwRgETfQcXnvlzyS
o4O3+VL28Iba5PZubVnS4jE5JcaV/HlG59GrG3l8pV+045KQpCgZR9DGMxM1f489OzhWkoD36ax/
clhTZPvEl3eKHMtK29szBP/cNCYHs45aucy5T6ZA59bKmKsmh2aWrGicDQhwFG6TTm/Zn99Vc0w0
ENJkVFQ2MGLMb/ZoseWf8yJIp+wFb+dvitenG0i86FSpybbj3IFajj9LMKPB6SYFRemAiFGSrdH9
W+BRyduJvmzxlv7NRAkHpp72ZxMQBaycFVC4JdhQxcxAUnnsvmPL52PJWob1+s55sxPaMOez2Yar
VWUUT9LaDpxQfncRifHW8gQszaFx4iDIgdhuRCZfv7xCCQwSj85Of5nHuZuqFfP86HwaZ6bhyv9i
tkT4BZoF+foV9cgy/wW9pKo0kp5WxcU4tzE8JqMMRmScMGFYgT80svIKTRl2oVa6764wAY7pLrbC
rMNEuRyVS0lbPjsOaLAigDmVUXblMgqyU5lhBlOX848X9b352aoQZgCEg0pXTwzrKZ7+gUOamG1O
Apc4Y55//Q7UDceq+rrIoVBdDaFDLlyOivZjXDMU3qFulBUU/B49IIqWGH5eKJ6e38rXPvGbb2Ro
W5lWM5+BEgCZTbt2oSQNENGY5fqCNRfLUC1E8ZfHnWxAfBU7a00C6QtEvuILQNwLzXll0NSbsD9i
+FJT3fUv4bsTGa04qXal+TcCrotvUQubrLqc0eUedbN/+xGcGyHG8oh+Kt/gaxd+fslJ0YRBqr+x
2/fw1T9/7/IhAw1xeS5uZip1OVOyN1gHtvzBfgqFuy9vpwa5J976KFtLQ7XEFEt6T3j2dhuFCw9t
ZygiagP9QQEsFP/1FX2OJNcwzjVrpbO6KeBT1uWF2dRVyckOD1Sxtgv1biBVqqkv6pB+8VOSc2uq
0khA4Pmf+WPIGeslu7CRSrZPqkX4EF0ph44MTcpwfKnclSjiIkywYy2K3BXABhZRF6/letK8kO0G
bPbLO9Qk3Q7AYe7iul33g+1nQZrP0BxyxRLHBAxe51TBNYNno3WMjmFhWUkNya+7pg7TICl3ludk
a+oR0nEymqu7kNrOwDkD9asA/rS/0rysw9ZK+2duOB6HQbYOc+uxo8VfwzmawhPe3AEiBAE9WY6g
HCoDuP0WKtdfBGkvWsBT5OU7Dwrd8VvkxbnHS4SBCEBuOe/Kakqxyy63x52xrWWfyJRMvmLS3J+L
Ttzb+pzGTcBsgbzn+l5A/9uQm4RA9SYRbEKIUu/TVrCfalxcdJ8yYn2o/EXlGU7YGEd7wU2E/o67
2VFDWltjVwUYMz4eKPWIhuulJxXx3ahcDb2JCAXgY7s3vq3Kz2lCbBAhF6OxZtMWLZmAJpIbxMlW
JBrYOI4v6pEKj/HXHW9DU6nsZa3eA9ej3r9LE3c+NrqLPqefKcIbKhRhQSqUtauhtvIXVqpXoP/b
PLXWYe6xZDVelWbzOLzuf3k80JDzpeETZMO9MqiZMNyrLiFdzF9F7FNeTU8ExWDPtIOGi+yRcZ6o
00ba0HkpGi3QcgUqz0Qkpjq5skVuA1YsUvoLwTKqJQBQGTymJ3TKPTKEHoitWJdABSFty4i2clC/
GOHXWF2bJzGGC4Ui2K2gT51YSVJQ6ztWiE9XJWoYNynTWzmkffkWzFLyTok55cM+POjwSGAh0iJf
3JNQv9EyPe79G5FwQHKntZVJrY/zuoThITJOua3t1dZeUI265dKeZ5/CX32GReSZY3mvOBA8i8tI
2Ca4Bdim1qAU1PqHGCjYRe/5EFDYQz6xGoUDKHoPyo1tBEVTfd/7Zosp2G27utiflmKMuIhuA+WD
LTFeytwl/+rru23VFBCLhgW9Oyt/rbS97fw93K5YPAP1f6ibA22PxQXW6pJxoIzWhKpX5BwBuLPm
PLNmqIo9SETOe4w3mRCqFTvIERy3S2jM4ifvVTMx0q51A8y1wkQ36gqEu/114eG6co6OGzM4fXlk
zNsIc2DXZRuoLyt0jYCuI0ZBP8qmOQL0BK3GbzoeAno0UGaf5aHenAQyg6sqndG303Vxgg3HgJps
ke2RoO+ZNBj5mBDl2X1tAzzOg3T2bEttGLf6a0mg9VH8kwAcnIF19XXN+mEtguDHr0FIHWbMuKUb
SophsewpBU0TXrrjqwCn/eIdbsr3DxN/jH5xe22vewgum2cv3jmYipQwycvtenCyrB8dUlxVE44/
pNB03EcLuspiL1xDuorLV/IIz10hEpZSHHmpz8OQIHe6B8JraZlyJxVjcy76UApU5VqPH5R8+e7G
DUm1qeWVhCPmYT8NsPJl6d6MaAlOcH3b+a/B05WlTX+gaquKvd33oxgQjz7yxAB3HG1GI4K4vJ06
LfNT1IQYSOhtUSlKSlTRBmvP4WPISJDKdIuksdvR/RDlRa/ruALs6EaY5OTo5vE3j9f63NqPiCyG
xf0AvIe6Warp2xFSidai+/vLYEwdbyGYxK92Y9AG1ewsjZkgVyJ1yulYC10kpTG9aYRjSwtWR5Gt
kXOGlRMySnpvz6JfECJ1cw+7irn670vU/3EcXR51EeQ0Cnb/mrgWnXBfdBlSmhIIQlzYTHflmw3o
dMOdlF1WL9qLrCurlxVar6/SmkuoAISRTl+2zZNoxViVBf/kiB3wSzGsIRVQacitMJaf4ziZeVdD
v4RX1g2pRgkB7GDglhjxJPZwuoBjcRxTjmCSQZYlx04kgauFQ78xRIKr88K0O8UNDO7NTd1CMoFc
E+IFNvY9zTvQmkqlV7g8UpkGeflDaO7BJSnQj36o/i2R21zFvrh2hAKoFRVtL5hKZpypNCW7ZEQl
BhMasVnITmjJvKQjaXfnbTLOsDRplMeDJgfChl3ZNzGwcgViw0VWiljYP6YpV1C8pxEyV4k0w5AI
GHFmzcxKq0G7JNWoWory/0tRJ1mLSpUxkOcXUfXJ03PE2LsEZ/N9pVcGCbKB3hLNJQdJ3frpOirb
HS0PdYx1chasS1ZO886jXGHdW500Y1UJxIIljRqH4jZfPhzQhcLf1aLYjfHwET1FdrhhFXbm5tUu
HxjOL1YvlemtYEmtSbFVOVSsn5pxkYKUGCjTm6ILUj0yajOziR3FJMqUI99HWK955BN72McA1zLV
wP1ccF3+Ftf14G6niPo1BZJCz0zOWAoRHaOzBrSMKUP3qMDQ3BG51BoODXpNJROmesE0Q6y8qnS5
Ua0ibIGFBdFr4YmbJZ7IHGbj4TUpisNDFvzwfPAdoCzv873Ni8jVwtMvCpC+Z6yLls9FdC75qR4u
3nNW9kYSt0+2PTxHBWcwBlxgO7uwQqpTHsl/85GX6AZezGL68AEWvMq1OGYlC4LwsV3SamRRcCt4
YL7pv4poYkDF7Cy9J0/whVzn/jWJj4mdrCwu1U8gQakVEG6yBcTEsYXzb+4SdkLaSTTkvXno0ym9
4cRcUFHegI7qHVe78y0KFJH9lVSSPf6cI6btvGoIOVXbGRCrKTfr/YixoBvzOdKCmjjWC5cuk3kR
NU2BoDoWJIh4ltpsyM1tfK4scDaOEd4N+E322JQyiw9/HUNJWK9Z29txKHyLGz/CKXRfmzk9KwYp
2aclc5TpXHIDIFohNLr22ccgFDI5j360kmbZo2gkzRVchw3V6q12u5RKZvK874opncCMV+DFA+BO
nA7oqoc7nfX1wEwp8GkbGYy5gthOHKvc2QX0FzKO8NX4bdgYZK9Aj1XKQ/tba+dJpkhSMaQ9v449
6AQiOqMzIB6imoSRjAqQvsBEJCp7kI3a36mvovS/WSuCvuvVJvHIRBeXSxHPyNlqi+Hlfk1UurB3
nyDouCW1mygJJb+mf9CPEilm0uuZUsFDZf6EePkHYgCRloqBTFA33gzaKe/Dk2eyQ5AsmTnUwXfL
lWUijdj5lQcgPdai1Nz8RX+uUgoco6SBHdEJS85JQ8Ov0rVfiCHrTc4GAajudUbEcrPODfHeznRB
YhrjI3lTwfvt5wh7YKKriig4bpo16PkMpUjBys5y75fQIjeZL9s+h0nF3B8EoL5VwKMU1ppw2ZU3
OgmLYcpYeTmQdsG1Lhl/81ODjOioe38hUCZ0/DwSIcSu+Ni066sPXqCuWbm36z4PP9hg2zrE/zB7
Ot2h13c0TRkxH2WZx8VCRxXSiY2I3y/PuYtYpNBaZ5wu/JePxuxOUF7Ybz30JXdeTU+Nel2sSLXy
2URMOIuvqBaRArZoTXApl7Z7XJamDAxZAh7xi0Dp2a96MvUndW+T9DE4dXLurSik/EXLrheSfgEi
K5u7yRdvyslMHxCN6sAt3tll2zhTX9zfvsqNSkQIuxL0vQQG6qNSHiegNsm5HCnhCXuGUoGX17xg
/GQQM3h10TSeEhdOkDPq7YXXKHCPxmPowQIq0sseiJ/Sd5f3Z2ZjJnBBKQcZy7iYMiypJ8qRs1MM
UA9HIX/s7RRWIxJ711uGxAIQdPRH2KKnqFSNVFfqi//zn4AOJT1jWAsv923rqpjSD/TjjNFo3/Sb
43u+G3Iqogy8rjUq1VndE7QiONWjgklhCgD6QoNhl//Hsi1MmoUU1qnAlRhTgY1p8Xe+p+XEVTBk
RjY354WUw1eSmLK6tCxrUdonBV+ti+vJswuCmu8jiwU6xHkLr2hpBA6zmUSuOUMHZGK6SogUWEzk
O81WLw4MVwT+jE3eI5ytgfR3RIJnwGrz05Nj2HG7o7JFCdeHvH9Q5y6EGzWSGvP+9slTxIXnoQ+2
1xofHOe5usBupB9EWvG3HDWpRx2rjyD4RsyXoUWIAJLIxGkAbR8b5lXybBVzB4HLIVGEWn/Toebv
oBOc3rLk6Xa7VcgIsyhRVnbBdzhJnuUWi5azDqjN6CqChpg90j78CvCIml7/aeEeJwPLrpNQuhe7
ToZSyJt9dTYIRtPwDzUXHzXMjesa7HxY6pWYxYQdx2CI0Fet7akKUlV5R48ir0FZIrLpwP55MLBB
I/45NfmgxCZTjAJ4PEgP5MbKqX+sVy4bkgrVua2+PY64ia2V+ehX1ueVS6NVC4NSawoJjXy6PJ+d
9y6NfxYi5AVAyG6uw/+VEQTD/uSBhtjqIWlzA+aZTmujt+YQ7kPTqd1lY/KAc2arHSAO7ISg7n/H
JPCNSSBuwZXzk9pAdyanJkS+HOBYFle+jvwHEcG0K6nYAtqBh1S8VRkkPqLh8GnvFm0qJKtQ63HZ
bd87/A6rHUmqneJH/B0PLYOnXGyYS0YWf9r+OL8CnZi5vhyDrr3vuH1DYodQtSomYhn5XAtcKvrA
tnx9IwdKlvDeXSvuPN6JzdqqCI0FnO0Kw50wYuzHuc4UZEaE0FSxmHzB9zNDKNwQqB6V0jdvDg03
jfbU0ExZgyCry5WiQmblNdXIRNKavRLvPFTL3XTP1tVXXtKRCB3jZpAlHwZWG5IX1qDR53m9rssZ
E5a+5Ltphs7QtUjj691dYiHHVJ6cZsjwcXpNji+9f9WmXrNyC+/2XgrQmxRd/yzMnsvpe7LyCWvf
+yW0uz+3SLpdKTYD4Gol5viz8K6wscYnvo58NNgjjD6sFqkHoLBnfDAXjDnAfJ9gDdNYxta9mrUe
DKZ7v5St9JiMj4coPcRX62+8inpujCQqn2AoHDScUneAOfWoY+H92KTdjGCVHnBV9D6iJSGNZzrX
Bs4TpdobRds5v+l/JK4yC42wadHOWRH3fmTjFSgpMvdLGYlaXUxYAK9KWttglGLqW0g58YTB8wIm
POlAPb1JyWj+HE59oxptsskNOOrkC2eLgzVCU/awrKul3c4eW6djDd1duowdAQ16jsGzl+VmuAVh
5XZjjm4Tewh3EQvFHfxyOj7dtr/09ybj/kzTmqXr7PJxztafb5v5c9EPqBm/P4MAM0oQE3AZw9kf
PM5OLU3YYrOXD/nrAsk2/FVUZ9EQrws+ARLVz5Cs6IlZMIOvN1xNsXgOn6i6LFtl3k9Qs2wkBfyj
MEI4wj4jLcEfM8Ep9AgkynV5w5Zfok/K+rg6LXUt/Xa+0AUuQT0tI3KMNvETNfe8Rev0dXoZTmKT
1AWZFzsTtHOzw1zPzR3RqyFXPjTyUGMNjOz/xmfCmq37TGXd0OXxd0rhQd26gm0C8jQg3B+16lMd
SKoqO7eX2tXoNy1ktjczqtzNQAoNbWgzEsxV471lEzq4wS4kQcgXOTciCpW8zB+WPTfZiYuGUeS9
FlNV3UWjHEMukRJL8jjO2xmKLgiRYqHRzCigs3K2TgnbzInNX4hhXIiVWgkZVTjL+D8D+kO6wvOK
jhZ1i1AIkE5mSsaau7US/YukTNdmVhaegfolbqjLYZRIV6rmxYF5q6cXSbwK2YaY8J7wx4q6ctX1
oibhHUa0BmcSF5xofUoelwIU9//NwElD2m9MjpuRltKCRkWLOKgtriWyTBSw9DATPYmmx8e1zUgN
gMFEvcG2Lu/J7ZiBctpwzGPGbrnwbPcC6Yus0uodNcEqQnT0cBlQGj+fBQwBGZwNkTYjrXGj19Ho
uARGJPHQwTX6xVadHReT8WNpP5Hm00upM9VuF26iM+Zn6VxkXNTbHcF4ZJtmojAR3P0N/OP9c9Kx
lNXFNs5LkYX3r/jEw7UFNz/Idtf76XPWKpuiw8PGJQFngJWD1eG7zyJPOoAVTgP5mGGUWzPwxpNi
yHvV5zeQMl4UCg+BbzLPsCxKg+8ia4EMJgz3NfMe5RrugfC03jpicNjKoSZhxFhU47VF8HuzU7as
BFkuGeFnnlogOvmOGHfbiyti9Ijim0Sk069yTvyoFqAB9/hVC5yaB/Cwn/Pzz8F6W7uE0b29vEnp
7/68QFIh9H7KdfHfEJ3U6qLJZ0khta7qMpE28uhfghdmuvJbgq/6Nl4eC4Azc7BXm+Oaa5+wTZHG
GJ+zrM29KHVSVBx4v4WBP5O1brsmD6zg/omzFUvJiAkw+46WDSdr8kYV5CQrJn0p6PghY8LzFeF9
lpH2hHvu2wyZQ7B2tAQiTibRt4d61Mrj4Xj1KUiNfH59BqN1iOgH6lPnnds5tF4Bv3M0e7qVp4Er
uZUCR4d5QB+SYN2z0MdTUkPhSTaZrISJaxeHQmGmPwZ2NjzN17cSK+t7aQ/L+/a3ftNniGmnC/q5
Gi0IgWZf27m1KVRX8KCHpBJOfweibZrP1dmuAbl3zhBQ2PNTaGXwxuwCh4P9Ma19joxkWvZL0l3h
ccWwJUF+8VuJHnY9j7DAaO8omvlfYIng6rmmnQEGfbSSxgiBz7ZazN0JQc5L3c0OY1f4C7A3yQ1X
BN8Y9HMKmli1WyxYPia7Sz+uF3GtryDHVkqCH1KuQjn6YAKKhrKGweIy7fN4nv2ibjbyX8tZ87Tb
Yk18+bfacDjKpmggG/++TGVVgNiyXNs47uSnoKcxPvy/PqxhtYw+WBc9nziIu/vgEgb1QV1AapMV
NBUPcw7avzfJ4qXolnNGzAoFjw/efhaiHAJyJgar2Yp6UjFplgZpSRwj9RowjJdA2689/qIeDWfM
UX9k7K+3es8cu+4V7upjymf3b7958+2Yw8nahcwbhVuSmrOIXHAHw62KL7q28wpicB3PQH/eqU6w
gwJ8hGKUfSImfQ3eTVJrwRwfnqvpUOszAhmnLUYWrsmM5+7saTPvPgKWQjNnfihkWtUFwYR7cZ1s
CEu+0AIK6ICtV4nIC1P0gUnc4fKwbLltxw9f0J2PoLnBJQvTQ0a1RtjxivR9Klsqnql8o3rY04wM
BJPiyd/+FheDlLtOpb7icOm+rxwwbTK51RrL2P7BslyRLpeqQZzFxfpBHDFXUaRn7BLTvKl0tGnz
w12RsTaMx2W/J0oSWLS2Oe0IdC/NmtfXELtGYse9N/rjmuGczT+KZitEoeKsEo6x6c4+866/PwrQ
hXU2xesfMezFFnu4RJ6WpPhfr9nd8hIS3kMUnbFo3SDd1hcgyXaFHuC5LgN6QNLLbqD1J8bjotvj
vkLlAa7GyrMOpwmowqiiW/XFTwXe9Bsm/D+DjdWRBeS6PTEzum9Y7Us9ZG8qWraFn/POBFKeoDSR
rodyO4kD2tK1fMYJ67PGXt1XDW/STPXkZd1uNaYob6pQh/ePID2aVtslwqKbNC3GapXb0u3iBFoJ
4sANPtBSv4w88E8je+LAh4FieC1sV7wHBBpUL/fxxuDKIcsK/LfXyKGE81oM+vqF9G1kU+xUTXHE
5oXOUiYxiVu9zedqgRND8aTzwfdABSBk0+0cSA3VT8eYv7bNeCPvhYNtk8TyriGoawikmJGNBWty
RM5kCPSuT1eDCLvJuILChMDVK59PMmTHovnAlRN19Rc1m49NPGX5iMVyKwkP8aK0jUCWFsK4l4eD
yPdKtlR3IPvX9gSZ9YEmoE9FLZM8i8dW5yj2UpJpWk3WIgv/KFl2OSG7VKG6KTpNyELI3cbUoiOt
IuH0P3mYXm0ipKYNjEZWNKz54PlfCFU13/suPwPsWaROAG8J8mDstl2dmggfRT//c4Wny7ZWXv13
Z8mYnmhTlKfhv8V7v2h9NE4WGrbONglrt9b5frHhv5liX+e81zG7Sb0N/78igJprpepL9NamZUqH
espKiN1KeEjcXJoaaoXS08tqvr8KP64XIyt1DEOcttlgsoKvMDrF2/4f3TuZNaTwb6vrBMNLPsGx
KO3mL0IA7E1BEruTXblc6TZf6aEljyFbVAVOUwEBA8RpUUUtKGY9cEnpdEh0FOCxc17Se9Xreo2F
AxP5euuaRhiRRDh13hitPS1FvfhpvU1BSgx9P5powfHgumNVqK5L1VTtPkV81hzHKnsOqAZosKaH
J1twiGKuSjWVmvDwd59ompUOSJ3hMFFOebftW/iubqKvH2dkKUKhRsvoM3dcLmaKbb3P/s/vPtNW
rIYWwqZ0dcmmFUH+wwzUHUN752rFS00vcvawC8SVo12Xhiy0fG8mTpZ+Vu3G4Nc7BMWA9BtCmpSe
ZvaeD8uIOch1jHMHbb1q+Sdz935l0nwA6dhXAQ81u8XvuL26MkoZFbI6G7B3RDNafQqt6KV2P6lm
VaRreq7I28ZxQPUMkw/aiaZR2iGFUSJCXauQOIQX09vUUr8i0it82phdJ47/ZLVoACN3v1btfqxU
BeSq6wF7IWegdbjxC0vXCViN5Bmu8yzKvVEGeyh9Kv+aI+rPIlOIESAoj7+tSzoFIjaQNve9ADNu
ubC3V3VV7SuRCXgujpm7sv4aINMK3kmU0DCoOvF/B7uA1UjPXHkcw7QYJfsDLS77xcsgDEEJHT5g
ja8GggnTkUQhN5natgCr1ajjWqF0wNIxG74Go6iOBMqosxjBoRUmhzz0cXMgVOfsoV/DGyUrcON6
qWD41aoJAnM0tPYeekxQgaPVxfF3zxRosyR2dkdbN0QSFRTuWwXXCEOyYY2sPVtczAWrRBC7MLgV
kLpFHxRqkL4bXF01dYeYyLQxNrlF1IK0mB8Njgaoi+Xa0jZHRC7tYlOKHcGqa4vwPVWUP0buXlgP
w5Wk74b1Zmn+ktH17TGTmPNt7px619TI2Fs2tl9UDxYKK0lJu+uNHy8a6/jmK1Yy3a6F2+OZI1um
4eauhFzwrMGiXgaKzzVCfonvsj0yR/Y7Q4LZkd7O7BrF00EVSLkbOYxCesYyofhHEQyb8PoMnuG2
WiY+Ka/p/NwIPzKOIrZ4ga09UCjbirNC46WK0x8yT8pzRiCbnBKSEAs5QQDNrQ4phtboRLH97uTz
HtPvJUEkLHDTnSo6DHM2NlB+4HWxMnl0VOkXg/eVSXj87rN7iUqTZqqqh1RI+MhmgPz1MCbUrsC6
fkmchNVL7Ld5KR563qfP09nOMb0mvjmKb2JmEaPsQWiBCDvXICOheUrUohOH+Mq53V+4GdvwxVGR
kCMaXiIdAGZSXlTBdxr13EwnLMcd28cSH9Pg1QzPwaC2LIuOsgPcnFtgc40A+4EVc5pcXg4JZBFn
L+wN11lVgWcC8O3socTRBi52zrIBBRN1mArw0J/o8gyLKTwPjahI3EIKuFajx8ZQmLfOZP1ZclOy
eWjWkcX1Fpex4Zpg3h1iagn3JpPYy8l9NjyZkOPWb7BWrp6wLsGixFkrhCOEtPDRcvhfOtLL+Me7
CtuOy3SXcVV4AJC0PipwDWe6l85v8OuoNnzXUdntznxfz9rF1YUea+HyKddDMIejI9AZhPErMHrd
RRD3mkyDtVjHNRlyYn2HDN+Qp6X8Mxv3G9o1I+fy7q3VCTyE1KBV9tmoGTTWDv2jm88xcEQSKrkZ
vVUDTtRyOMQunCLoh4z7qTlquLu0vvFznYiPV6kA4q5ulPBGGDixmJHCY+LY5XfUQ1vgIRc0jl0H
Ul2U8Qwlz0m9HtcKNxVnG4JwGII30yKhRZrLcKcJV5zGR8YFoNCCPlY/eyLraULLspxK4qAL9WtT
jjhbsv6pLLms32miqjqiBKUc4iKGbMrTjDQkOqX2igiEtqfdI79FTy3gDdeoGkCcbJYf49eguZZC
cPPBRMhM/npbr48BCjnI2HghqJaSD2It/Ncc1HTN1BLry/9wsmg2RJL1GFkYnZHyBvvEiUFLPF5K
/jouUVwWw4CGrOeAETXFSCH4qsiWS9JRSmGBcmoKhwlkPgNv5IUorbJTaPNru8XmJvrvgZKt4hDH
PFl/GOCT17+lzlZyhC2Ahc5ts0WcKBbSM+qd9boYo0hi3vvGx8PB2C0NyOihFwzkPYFHlT1eWGUD
IcfX7Hrs+oy8np2GSNh+gu+9HMpfhdc1U087NtXoevpJdaQGYqy81VhDHtK1yoOU4nabbZNhzMj/
xggCxH47BDHzq8dxpBTSkiWOn9RwPVax2Gcz9OoOxxdWefbywARzj1NOp/ufKgFzDj/uwnJppxG9
5Diele2JmzywrTGPwu1t2eLgqkJhaPhoqJCjFleKr5gPxyim+75GKwDGF3AO0ueR46FMijjkRsyU
XEviYjUVZTd6eU4IH2b3367DOlzDpAyHfrX/CIsD6eEdq3JH9NepS8HDPXOhViBR242EHUCGZold
ubRqCQCd0YsDm0B1ohmzvkRHcJ24qGuNaNpH66llyQVA0Rdjd14yZd71y9KO+kRLg5OVr6QMrZ2i
L8aLfLBPlK/JEw12uX571FAOg2kwQgl4cm1CjgA/SdB7+jhlqNjLTdUu1Ty1BwfgRYdpLD2H/4Du
DqrApdj3Jq8UyctPoH5nLLiilqx6IdZ/n+sn1Qtf5NoPzPiWTz8FnKgOXLTzmVgXEDblBqWNnxxr
4THzDu97lnDJ03uM9oePthy1oCjrbY73/wDl+aysviKR619zpSkuv/AVBNWmgx4IXmV8Ei9mm9NE
kKWHhqGzTvz32htUmqT0p/VOmRqJuoS4wm+LR1Jzmpo84ZCz5S27QSju/MkR3bbbSFONIoSbmuLr
t4TpLETTfVOoS7JfJipenarN84wt2WLU6zEiPGvqY+stcw5OwdOrTQ72d+DLKUbOQaR/xWr8Pbr7
TJUHV0+LUisV+0be2Vt42opd0idSZOx6LCvkffuShlxM8JscBCxaPBEfDgvgY6mW1Wi8AWszm0U5
6lo2jxhO5QcgX3Zfv6EpI4Y3rO6bQdK+Ki4uUr93vPgtWi5lpqfBMZvaslwQ0J9o0Kp8Yp8xhS50
F1hC5KRQvB6MVwQSqs5ilCdQwgAiAGPlD0LsTWSScriTS+dO44AyA4bj7PfyVQZps1XLmitltC/9
xLtoKxKLVHuN51THaJ86fjekt2GvQc8iWj5k+AH+SEKEruCtPxua03+VvtAc5IuPW+WF1T3J6A/8
F5Sz36PPh8OB48QnBIGyEZqsTXMXuPsCetwPy7YO++MNeXmLGutnZXQ3NA52y6togL7/do94bnVt
lU+FiV5ViwbBefmBrstTzcryfmUvzCE0puTbi8I7KR913pxjLMpg8p1Xt5UOzZuC+dsZqaK7z3Od
/v+IO+zeCEGb9k6oHUUCwMfAMmjlWHz54YgrAN1TN+eHlIQY4Eiz/Lh8azarR2XbtQjqWTBQ/XLn
pLVcUNHNBIIOFb1Z3WnV2Y0iZaCelW3PB4+y+6wGqTopb/OWPwR8jKYjhPlXnKrIL2fZR9oXkQgM
/hlobkcEAUFvjXQJSnOdYGf/LYaiFeCrWecG3eU/e0AgUvtDltzfSRkSwzAUiaLtF6y5jZ97NAfl
xFm7rZW7oEKqdrdPWIBtE0Lq2pBKtYcVfOAXbKl0yMxZ6GJcElJ+TgtoAU04qk98/uQQlp3joxBF
rkugAl71nDFmpcBnwWAB9ks0a9PbaijlRhNf5NG5hvpo6NNKm7PkFHvh+2XjokVe+/G0L/HBsp3C
94yWAxE+vKFkR7zOXMd9xlbD3S0tigovcFfsJV6ynK54jy95dw/nzE4kGteYgmXRo7JHCzhXO0Ec
vQGGBGEQ7UJpERyrRKzcPwqyA6MEu3yoWNzyaWgm6doeo4o3OZwOLWh38QXGQQobwT5d/b8qaCJa
rfudivG76D5fdxr3dpEdYSIrOAjDrD0T0uZF1zoNi/HDFwKfxRV2gntatHNtMeB0828Zd98JaAoE
Dmn8VL2L4p+Fk4AQgd0lDK8G0AIhJyQP7TMHEMmK7ws4vjcVIo05kwCTtNAuUs8AmEj1Fhx0s+QP
rs9MW93PyVNdUpezyIhi9tAHqZsxQ5fwGr4ui38Vwk8h9AzQBAiedAOmn7MmazzIA+69ActcoQXi
1HxJo7m3RiMAG+vpwsO3IyusBukz/Nn8hM5MvCeyg9BRCw7pbb+vQluBvbHAj2b5fcqazrF5JcUm
52JXYBMynLDLrhzg+PIvoUg+eiMGrU7mjnzYG1sYOUBwWqiWrkizlvnPlkvQxTsDh6WElC3dCwu+
St7lyyYfS586tFFIBzRyJNyc95uesU8hmTu2hHQNbtojr1zPMJU/bcvJGemuoekjEs+uxxfOtxbr
bZ9CEQu1ayRHbcto+Ej72WNwqnRqvg3AfCvdXyKJrZjudCUh5kF6XJPE2IMkfXnlaE4KStwQcztK
lTXWBn0BCUAcaL0/IpBAfwvuJJuA/RsyCvF/Cx+KxRuhlRFEPzvihVJhyd9kQauVnJqiVbKo2fVo
8QB5HW+zxqaZ579Zh5N6FqWmZp9291YO1L4OaBuSkATlCjU80Cs0K3dFQKEnhyre2zamCjNAhu5l
ylb9oh+4aEbVDg0pJgHzl6nW/wh/Jfla7VOuGgEzJFwOciq92YiisARdctU35bO4G/oJHu5ICmZ7
cv+O5zFSXbrWLBON1UePNO5rnQsKiaODYESo6ed4RBBhOaq/0pk7cf6R5rKFqk/HETYgtS2PCvMt
vp4DTcD9cnZH5yy2jyYeCpoP6aGUrW35eLUuv1J8qFlHArlm8WAUpYaFYd1Ne3oktwQNd3o8bXYH
95ngo6abfxwGCCAjSNVWkBS6WVjSUU2fS6+sXyL5ciM+ctDnmm9nXL6nDFSkMXinmp5qYKveQrp4
hA5uCKLQNOlUZ9pOncfd+7RC+/GKNP//IV9ClTvmP83Cqx1TqX49FqYqt8U8Xq3NuQgdzki9baLp
k3yhvPkKIljdhg9c4Ki+6S8Q5XmCHqxTNPZki2uOR7yhd6uxqm4G0O5U0o6gv0DNMK6VRCJp9p3S
TzaVzthO0B/aqPHOt/UNPbt3mhOEV8W3mM5H4L/EX+2pF1LHSChqZ/bkK9teE9wHqsJ+jpcVEWJ3
wehY/LDNSqN+4n8HiA8YVLzgdHzUoYUVOsBYDfonxrY/rtqDgagvHR3WjAq2z4k/3ZQ0nzznbfd8
O/TzRZa/6lDpBgka7XfKcXoeA+X4Tri4NeHdYw2kGDpmpifuv95Ssi0Ohki+PFtIrC7FKkcQk72p
3ZvP+bspiA3CZ2cFCZI3scFPGM+7+UmN362WUi3BlRi/xeJHX5GWMMbzvcmA4ifni5By2Dlu+E9V
onZmwG6LmfMlYOLc8sM7riyaO6gavTzlCnjvSZ/4BxW1GgBrd7ToN/8BHvyNCqSGE0lNkm4r5l1z
Q0AOkYt4kJ5CtI5qBq6dVsoPzEgwKg6fhJPQVnOhqaQLSOjpM55+SUTZk3kN+GW2ZJ6wYfeXxPdw
rLm1gTatSKVvr9mucPrCADCazz4ZMCTalJAVy4QhLTihisin0uvHiMjgnQacxx6ByYEawtVzywl8
3EbpbCc4LhnP7LpWcR2zuV8e1cFdB8NGSLrVjg6TWa1dtEUWD/xiPhgFYXkVQkDm8BT73gun1eFM
FnLp8e/gZQ8RHEZnlB1iL9rCWJs+tHBx+7TgNdxPfvJgaCNc2pNS1D0lDjlh9O9vrAkbDK6azhqD
LAwi9eSHi7jFmRdV5t4V3x4FoZyNMmLW+ruoRMsA77z6AtGa1j/pKXGvh1szupgDzY7848Suetzb
fUI0rPrh43ld/jbouYMlUISySrsZ5eeJ44AbuA9B6DfY8f5dh7/ScnupjtT+sTy1U9QJ2TcZ5Vkx
85in+MiYWZ03RAPwX1FW3RhvJ5B4M1sN15aG4hHW4m4AlJs5Hmo+JKZVkE7l527A2h8fmtL2bJUN
shxTnbNtEr8H0arISHRQf8tfzgX7KuvFOyqyhhgo/HiEOu9aUtZ2zLxX4MCF4ZB7se/743UbPr3O
zeQelAuGNlCc84WE3Y5hRkH7TLnHy6Gzeg266Z1I/28RVOAa1jRggbnyqeqb6PIWcXn6zdpZdYJI
gN+K1hctrJvwh4UjiARaT0Hd+o/kNVtlxdwzihUFZ+gA9wpDuZjQb+WlqQQItX7ekWXWVaGQnSnp
Ios8OnsZOsuZbLmLGrFQhXJj2XOphVRPg7v1sNDbJgY/UAXKt0xJH6TmIhczPyj24mqz8W8tFzgl
fRREjErFefA01hJn+cLnNfCbeO/O2l3/KEsWXbdvkmies+HiC5Q7XY3aih3KBD8sinCZhgJX8bdx
++nnt7chKGy3C6f0Sya8x2iA9G5zY4+di7wP+ig1BuYZWYk8LbEBatagnGJYbB6B60SYDrudMwKX
YMxhEucc5kFTPpwmd3huGYhJL4+vvo8d1+07LGcgk24JgYGJ85Soa32vY2moiqNhJhIgP0dbbisg
rSD+qKC/WsBZUNBM2QsDthDqrULKaPuHLM8ZHQG60/ar5/PT6Y413SrqaZiPri0UKUtNpJbjutNE
VMZ3IC4AmQo4405mTu5bVqNu8TCXFFbPOTr+tBYpTdF1AG3K2uKGY+tOyWhIQf7yq+4x5QSJ82it
Y1bn7Yea8OnZXaAtnJNBhmUZNhARAFsxY/HYk7bKH5KoyCxpJIZH3DdWdHKJniPdglHbsRo4t6UN
HE4VD6LhBaEbHPPAluNHe6XpVCkv0lt0Trez0DBbeZtZxQrqG3NayQU2dfiUUjSAjQyK98PIBKFH
FkRZ40z9Dk+9aedXGvkBazxOq2tNddpLJ5qzSIm4B7K5lxzxNROQedsHPvIlC5ryAj/w4d0M+LbU
HQ/ht+LTfY6WcfUvzjQJMavcJMW4T6CKaHjCmA1Ilnvn5obayS3hILbbT1YGtib6NRyDczhdulnW
4Q6NBOA5cXKYbM+AQjgokYpYnRhZfmNHjQJo1ktekT3K5jEB/VRG1G7o1WjSRx5zifraJnqf7fl3
uwrr73rNR9Tfixpx24H8UW9SdRsXx/0oIFPFzIAxrvtUmXo8ZAjXVhCEYFBgK028Kh+RXxtcf3Is
2/SmudjF5HTcwpZibodYZUmaKNsUQfuohQJjWD3kKGe3oavPtKSEPSs9ei8CNkyU42jjij23ScK6
GkOMhmW02ynms3nbJC22rzh7BvjXrh72ZFANH9W7m5LwSle+xnwqRrRK1PlyIJiQYvMom2UzJoLa
eTntT293fzwKinFeWWwj4jooQWJNFBWCWJX0+UmES5VZCZU1Sya4WnM9g2E2kxZKCpI8RJiw0kgx
Du+kJiqct4gPYAET1qaeZ6SEyxoEwo9oP/kFe15nZmJmw4q2HcDYCT73ctOjqEZv8Wbaxgh8cyrb
7P6gPv6slNGDyCSOo9PuTolTofZl/E9T5dg87oLv6x0cYzYBhoNt9w1zXZKxUJ0NIE6MCizTQAVF
CHd1iThkhBSW605AwIJxWbkpld2LGrb3jM+ewD1lPpPyPKr6IuX805FoOk3+x6ME63cpC08F99ed
cnYqWur6VpRDCU19etmiDw08TqCIEz/rJQoBh3wOeWZtXcOxLo+2iUZdmohN9fQ2v5a0MNcFUdgJ
Swb6aD7TZPXRGbyYNf6QmCRXRmHgryLcknesPief1T8QRSmAEWyIrIIRJm1IrfXaV6CLoEUp1UjY
+chcw/3F0K761fbeUj4vlAN0ei1MyRscoEb0yXU1GECSb/HG6sySvorgqg2Wtc5wvFZ6y0VtGNAZ
d06RC5r7Gr91a9QDGZJiq5xrWgB+ADoJn2xxuAgTKCC48bSzn7ah0fhNgI37rIVoMVtTRBH+KQgY
kZIPJZS3N36oTOQ5Y/CZ3nGx7NH1O2iP2bkdIUNEvHnO599zeTJjmeiv70pA+xtWzs+voWEVKf+5
hX1681UmUbnL4L7wQqpsxKVSQWtP9T69wKNperQQ2+y/tB4MVHKZnyaMYpkEfR3YlEJdV6SKzMt2
Nbs1rDf1AjhyqSafBlxaWFMEUzm9irgXL5aQ6ZGvLH/JMLl/6Abxz/MTOxk0ceqdO57qFMF6Espj
4xsvoNgt+KgyZG28UQxY8MFCrSK9uCh1Kuoz5aUrrWsVgUTW5A8KFAhnBQ0Iw7i5h7D0ljKc6Sa3
tIsUts6/BGNbnSQ46hl/FcILzWCkv8yfPrRsmpfd4CGw+6Xx7Wvn23ct5lUpbTL/RTAblXfvV6Bn
/MB1vTcgDdcxUI2hB2cu8xrxBotyjRGl/FmytS9BtotXT+Lq0ij6YYY2z8lvIk5ff67baMJ82Loh
12B4isqp06AcRhRYwoX7Hk3c+Va1Pfu7vNctay/eGoh2eEa14xTGisj1ANkpk4gQTGYruhmV0TwM
aLMvtim6SpUQYjcI6gclg1cP7JFQ1FCmYYHcC0s6278BWis0vWMJak1Bkc9C8Direb/tZfK7IlzL
jw0KNALYs3a3SnlXdyspV42d4+LZFUadCfkUtYnxtF+p0B07AbqvvQUkIwK7Yly+4JOQtHN6Sg6/
XvL3C33K7Zs5n3qDt9n4GdY+WuEqjZReqgvCr5kbvsgiuzA4UrrwsLryBTbEb+z4XpbcjtTIMA16
x3yEwtuhjfNMujeTphUJgoU00eP9VWIOS+uZOgDlcbRPQfPQ5a9X2fsx7Q564vbKrESbzljI45O2
4BX5NcxwVwIAWBpjMELA/cdr9aNJDPbKTuXsIHMSchrRakwWzBKO+GH4uSDQNyZRdQhXDwq8Svx0
tQBHFrKjuSBhrQWS8V1E/gqGsU71xg1PnmCTAenjGOSAaide8AzDg3RZNm+osAqMif0P0z0QLaeR
Xn6CI8bqAaUuCnaz5TvdOxIMCExbp3pMThDDsThFpLZ8zOVX+egHLr1p9HoiEsZvU223z8h9MIVl
td8jrHJ0L3fYRg2H1LOrj+NwQtZSeB44DlQ6W3p/fKuOab46Q81DxEMmz+qhibuK3thc62oM1y22
Fq831tVX1widUaqSfvNFvBL8lgD6pwvj2266606VswTNFSgVUkk1ksWcvw7KdYTWIC6q4fLudSqd
1zTDqIj5diA/M2TQtnXoTOVFYOgEgc4NNkeT7+AIHLlv9sC5cpiX5ABoiOkcS5CiMh55Kc8IKLRQ
HyE9kjcOEbmdsOIV70WVYXhZbpaS/xvru5DCwSX3CuHoAYPJtxvF4iHP/2o6UhIZxS1E7m7kkY9c
0Y1UuSlYsKjomXq7BoIzLIbG9PQ5Stsgq4xFzEElvVDbX7EjaYoiKXYXD9/G/vLqIe7Cfvn12o8/
+9rBXLcXd+qNVmR9GEFpOH2QLTvCEHckNf6EXm2N+telrcvOqX9EJp21ZwVS2CHCZWhLAYljczak
TK1siGvRH8fkNllJ6U5IqTsCy/ur5MF0DtgqF4aeZJyCdb8o+j7eee1l9mDBXIBatoTW/EzeBer6
n9dv+i0RRnGm25yz6xCP4e/Qrp/yuNp2Tbg6knRzJmutwwIChhLrQKU4nrDRQl5dpylCHnOtqIJr
RcyNuEozm/oiWU8ahlDN8hWRFPaysJIjCqnSDxHyhagb4yPrY8+KDoL+eNc9ky64JMODhMD8Fj7u
+EJwfQTPg2kJ9n9o24JRXY9fhmWFeaq7W9VryEcL7mW8dyln4QMpP47TyjT5+ozyWDdYCCAKi26x
OcSURH1cLVBFl+vb7RPAg+bZdPap6g6LyRxdAkcZ2mVukDipVlxzwZp3CFekPpYKwtxS7AOBiSLi
Ocbl2SxdP7O+1XgOGP9viw9IgbhVELEcADdQRGY7fTapL5i3O/kNyUxODXVRb0yUldHBfy7RSI1i
1bicg91aH0bR3gKJ9BAGBbQ//yYbWFMv9AC78WQfDbiKkl/lwy/avl3CxuoF7FIzDIsP2ff1lmgm
IBdZXXlF9T4d2exPocgkd1e+hRgBfs0/Ho0VQmY9vEiBgBANiDoVThnp7VmW+arMGPQxA9E/uAUs
IovIoDcMHt4KpEQhH95iGXzC2LaW7Iq0qxZN7sIbOmc3SrZ5fQ+doIxj9G25jvYSRj/6Q6z4IyOM
/cM6u5iGfN4c4QcbDSCrVsFK3MqZ7NAkdFN61ol8nwRGdOooBPO+n9Ehtjba/zIsrUBU/zSudr+8
k3eL5P8FL/3kDcjplyRpcGY2LCYkaGPvPJpr5emd/4hVmJS6dgCBAncadAALAhJ6eYcOLcGLLbVB
uIoAufmofyY8My2fFjcdcaDYl3jtKYR/zs1d4zKyQJWo02EMnXb8v61RMt3hm3CVmXy8fbUL7+GE
drxKjnnpc0wdbAofcdThJ5IWdfZlQwblrGvqwcop0ZTBjE9VKTDiRiS1JgLM/VTT6aMQgwiQTrsD
RJFHvgckgG0T+CTVHnAYCDucQ2HfC0Uw2xSxzLu9GkXSzs6Ok0056Zv8luDRbC68nPjWSECB5ncZ
onUrKEpYWRlIT0vocu0sG9HjJ8adEw+fV9UPM0aojE/F8+7OGgRVFnaDrTQK1O9EDGia/F386V/A
imznuoeKKSFrz71NGLI3/G5Oid+NAM4SO46A5ptqFZHEANRl9oN6P7iS0sE8sUPA15ED8WqKrdXP
KbDeuPIBwqkE1Td+rTOsOvoiPrpM8yHsKjPGD2XqAL5qFE/5SpUNNoOr8I72TJknutkb33H/t25f
K9NddNiZ3Aq9c4mEJSlZCLaERSD0mBi1iC0lrF9MDSQyRqAxjUq4CnJtVwPh4PcLrEyMSDV5MW3J
VPe0YfkDzttt6EEm0/pQVSXauS0Zcz3YE7LZ+yfyHTM6NiKm1tC8UEkMKTXktP+ecqefEJSNTWKY
4D5H/EX7NurexYF6RNaNG071qmBTpcEJ33R+lULZ6i4uHyUMASXcJ9PbTx4uhz8IHk6azt/KCw+s
SqBK3Kg49TBN25WXzOv8mr2C1jBMvb8vHH+G8gCLw3GrRDlVOQtUoJJ625TTzHQqqCZ2ta9EYlR1
HWxwptjcZQ6qVhnnBEwGAu+k7LGxccUGvxf5XLiVzZ+9YrohmNSLchsOYVgW0yaV3JT4ZocwhrGk
r5MClK8HuZSCnFt5mK9CBfhdWv1p74gNuqpxGEqnGXhPLzH1EnPaeRmEAKz2fDaRwOTdS3T7drCm
xfROkQQHZkCYCYSfwF/IUBrCrlGFuh3fwwl5bpYqpVHrBAm3Mp582998uM2Ei1Om958Ly2bS0Ij4
I84vp+IczEp86c84aeipM41h6qa9AbA6Q0tzMdwnycNlJItjJ0t74UGLpm1v97rwzWuTAz6nccwD
eswwqyCgGJIzYW3fmiA/8mBnBTPbOfoTqU5tu6pGkLk+wuhPcVCN0vCSI6phnFUqT2Lr9sOT+ofT
3DUPt2Gs2CYBIcIZ5JsS96tvHK07g6jHDLJjq1lKsezoS0iITBAwdjXI4cFXdE1k8vHgHWIeLJDk
gEFMDCY5m+loAE9TNGkBxOzRb+TQAsZDP+M7kPT0s7nYVUhBENrHD5i5lXnnXlb3xvqwTme/uQVq
u0a8w9UgqRxMXyC/oLE5bFeZR7z2TCsg17gqpH36DVZ7iZ+1I9Dt6X12RCMV08adoQMtTleVV6vt
3loA2PPDXRAHpte83zfxVkp3+z0T5bWlsIZWi/O4YVS24RWZYXLFokM0j4FxaT0kH0V3ZY/HRTZl
3s+A02h+7n29hN4z9QVxStUZOxtRJuDRSsRI6LYQAU/8ZvGg1gKHHYnWUuWt6XobAI7ukDZg3izB
NWqzt6UvZJdRpFx2zEH8/7yKl1W5BNX80f71MCcsaR52xL36AoVmbHSGmm6kCwZvj1oHg1e+kd3h
bq8Bv4kHo/y/O9cS/b8IxCpEOoOm6GE/rcWWyFnl4am5hVF6JYRPyMi4oahuq4PiLSywro7nFiST
hdqcixvtpQeAhgIiX5Fm1kTMlOJAMMRgXKYaIaFtEc4tn1rnkSlNACxFto7L5BLPfFkRdjgLe6s+
hcB7Yz50Rpoz9R8krH/G2h8VG+qtqNmHiCo8TSbR1hq/+g0W7UPuUueOCiVVhSE2D69UxluTZujk
+ut5sNDFcQkqsNe/qCWnEApHBD/3/bttWOvJ0mPW1v7PgAV2QUxzILB6MiW70vE8OS4C8Ax+zfbv
ItClfKtwP9SH1lhDsqGacPS36qbGTb11sS9waGzhbMmly17ETAO2m+O0ZPJI3/daJvKnngmASq6a
0biJe+Yo7Y60hqz0ow+ISt8Yr+BWB/gpCDcSVeoOHqROECrZsvISIzSwaCfdKXmIgiF4VMrbxGex
Gak2hS73ponDeThTh8sG8u2BSo9a9BSMxC5N1hYv2bNFI0rdGcBKUNvzbPaxz5wvtXiMTlCyDGxf
n6b9zvVn0n2naJPfhCvJNXXFcJl4M54e/rJuaPlkt1zQ8Hbd8uzKfcv7h4BqRcd5SZ/YiYcaXJR9
sIWt3P3+vmQ914DKGaS11yFFL+XUzCLNBlLohnypq1+eX4tWzbWG8+0ulDby2STHy3+WypAnSpS0
daNxsql217NZfGzWnoUIzs/nYXZaPPerxlhLzH9qz35+iqWIcIN99/1svkUtHk2b6oyNPbKN43sk
RYCmcpKKMmCUIvmc0mpNE705P1E1HsRb/EWkN3e/SJS9kjEOSTUyEu91ekeOD3PEV5Kvrqcda9y5
efbo01tMvF2Do73147pQgX76zx9hcckxyfUAV5dGjcvPLBToVK/lzqw1zldoOJwDpqFAA7i+TI41
tJwQLg53G0/cKx+qFjH5XTfOtyFGrGENCbdIJSANvnOdJ+4gjt+iuQM6LbT+mD6OpCUnCuTwDOWL
RcUtbqMYZhSLy8a+D+CbvZF8+g4XfF3/MOaH6cY6qWuzuVlSLI+p2LnTEazeOs9myfRhpQHAj9tx
gz2ibfDV4JnUXyF70mEBu5VFGjZcPUsbcechxmEm6seyO/ZEKWzhfNG8FkAR+cn9CWoj9/4LkvwF
J828IlCxIWL4znMFb5hdNV9NArGU2NfYjtp2RToROMzWfZrrcWB/+cAqXUXc/pjkDb3c2QcxOnKy
RaIpuoGkaR4iF7JOE70AL/6ABvHJgHe3MyxMp8kVoo4S2GMYd1lzzWN6noJFA6LIAVwrCw0daPRF
c4tg2s95TYl27Qx6fWwOaqIqhmde3DGc5283C9Qhkk+tFLVoBfxAmnQpoDEsehSkC6zg+PLLBxqw
n7VWqqcYUnmMVidtvVZ/OE60RMia5/nmD7rMjblfrSXOrACAlDE1hBsQu7swJi6JF9xoklFocwip
Pr76wwV93VsxY4kUZ6XpMxVDdOd2N4AeHeAXY5cxyqMDkQeHVSDY26Hp2GlBrlnnJ7IZf1iSessq
Hh3Kj2yzxX5YqP3clyQ+Q457tdISAOnT4sn1RNybxYp9LeyQmyTcQEfNaCeX5rSB1fOvTbfV7EZK
P7nJEkMaB+hcjjf62tRVHb60AvQfgEoNCJB6YOD93M/sv8lqL4bpxoUMrjsqVojkXM2gePBLQj04
b5HhduOT1MuABHaiVOx0RT3iqn1LO4JfI4Mr2kPuCVQ+Jctf+p/nkHU5hUdRUGRPKziTcLgAWvd8
wG6eoCIw9YsEbFV/EHRx8dzJZFMy3yn+4YJVKQQp8wwXh2dtBUofNUnrip3a61x/juN3xWoC0plF
uGKPzcDtkz1LG1BNEuP7s/bGOANWDQe5q/hYodTosglYbWxuEr1UtFeYVebCqnW+41UUGX0hsici
WwIop+X54UA3JiAs6S0W6NAEgXpENZzDvH90aMn8h4cWR9tVPD0Qe55wXadJIqAM1H24Ayx5ipFM
mkyD/lCfUzHZstCYSbLiyUgLzwJ7LN+dPbzRTlPMWCHKODZSVTfaRvA9Y+NKzDkhGTkMTAQhesc+
ih7c2aH8b1Qu3mu2KighvolzR+ypLLIBIjV4Y9+k06rf3HeC2Jzv1EI3H2SuOrH5Rgk3LTRbBrpi
fPWwV1jTOA+FAAy5PlcT937xwMhQ/ZhInx+19asUE+ywZmq46S1aIMYaB5VmoyZPbPnOs3SokRcD
ibs3OuypHdvTj6HqZ276ydnVfhLrXiiAkky703iAXVQ9OpljImDxovwn42QkqzA44rrJz2u2B2T9
jZyDWX2eozSHirUmYW9bjQXMz6+3/F5BeFEc7USG6/nmA7d1ciN+c5IYnlqBEf6A0A127bsXODng
JXxD5BakaO59X8SoU+CypEImcDXdxJzfHsPsUsszDoeRJT8H2trIjoZ19jPMLXOydWQTV4B88yEP
/ab+ZEpl+9mlXnp2lDVcQrLu3xMw4JnP7p/1KLsVmqi8/NeS2yxDyo6jXhDqK7IfcMHgALUh0tio
XGzAar9f7OOA9o7hNluCpgRnsLkMMT9WYFNanuki3eQRUMT6/a6tjBlWorxtg/IFiJtu/1Vg/gl7
bdGRUSv8g7axeZ6BzUxiDOR269oTApwtM3SHX9m+pMKKmJUskhABBj87SjL1IY1KX+/xQJDMSm2z
Nv137w01EAZMZA/5vN9EOmBpwerz4x96o74vdIzvI9xAQ3JxPyNPSZ0CDyk6PhL6A4XhkuEOSCR2
T0CjiXcIYfWpXPbFf1aUqRoV4yKr2xyWP+eNFNUeYORpgm6SJsN5YdpK8W5eQgqulmIxqsdkCFQK
BWx7UQMXY4SyLOTM2pCOFluz0YZzSxaSCGghwDDSO/jFiIW9/qXBQVxySewu1+4XP/NvLWJuTWah
OUhAa/hrVhjI081FDYOao7xfubCeFXV8eonDC6we6r0TsIpdZma/OoRDrn6IskfgxkaRCtI2l4OG
ya1V6+kROWE/s1V+qAqO/wUnC/eN0Vb5CtJk6QTCJIIB9am3cCYSecGMnBr2FxAEtBb3zKrRJW64
rECwfp9m9aBD03IFF4GJvygzw2+OflEgEcS7Z6PIZ0jLTBmaMEgdvM5rRtwFUX9k2GWbTIUfexpj
KC6gf8A0+VxyrmdxXsguw9Crmc9YHwh2LD+ZvBUWWdqRkIxY6VFzQMuU9kqjI5hZ5VU6lEKRu+mH
IOSXw5XAVQ7dPrLUCUEV133mU2bgeeMxBckjg+5ydA7a4/WfabAXnTNl+EtWVUFuIbl3CTVRm+9b
7o8iu7ivXoBBXqDNl7a77WLt5oYPLE+d16zChW4F9pzRQx81IJfOuZea8wvCuVB+k4TopoppG0+Q
1RbGwcarM0rjbK9rnIa6+QMCp5Ttzibvh9KaqEo8dNV/YHHZX7x+7p1q5RHSqTcS3UfsD+9B+i/A
vD/Pc4SpmF8nIo98g+zJrrhaLSg4sBKqFN6K8A8+hXiksGR4rsJSXooIbW5To4CVGu8urizph6/o
/e1V0r5HlvPhfOoU0ybfoTzi1jYopcTjgnNcgJjsY+C+7vIC4oCTsnATs2fWdzF9tdDzVmoIVqCD
XgIdezqBK5s0jKcTEwph+kJPIjPGNhHIAtAbhwhVCxkBR1AU5KiBXTJRzOKn69II5v87uPyJsJKI
g860b0huh8MUW0Wsam7YTIJm116NjwElcpYI5xQgMyBPrLAc9mZHCPlF5qFeVeJHonx6eF++1IZ0
i98iQD896TvFGdL4YbOHX9b7xYPRAG/ylsj5OwOaaPEy3AY2cdA7bK2a297HfDpiRGyFNyFC8CBY
s72yRWpv9caKt4/2cQewLxNEUWbMfHKLzngmEKWQKOPrUuACgFQSCStOxiIsi59OALrMqth7os+m
6CZgYegwoPT5sAcTE8VbvL6HNorGhTbydR4r9gFkuEwQEX4X4dhjQXjeg0R9DMNWcP+B/sPj2cIv
9V+CgP3a0lhpPisXZ5WhIyNsZo+6BU5VcEIUi6fV9XDUxMlk0TqVSTGeYPDxfWSwDFpKgk9axhfx
XlhqCGd4Ws1RS3xfpqodWqqybG/eULtXcUOZv5ajNG//ml4vZxGuHU/yEc1rEUEn6G1LyjDrGK3D
HpU/mNMb6S4y9dEgmQ36qsBUh0lSkU4YyjcG5k/EHH7AX6eYpSUg0UmYxCV4k5kJw0hKB10E0YUc
mVu0JSMsOFY0ft0tS+JActRqcmJpZ+6odFNDmrN1hYkNqqWxK2xiulE0ibj6/w2ZNWmnUxq/EGnH
pWUy/rW2bSUy8P4BDZSJyT6e+BR3/0dUobu8oL7MhTJoCaFTtMa7SajE3N64Ick/z+3xucG2daVt
HV74xiUJEIYAS7B/HFqEQ51clcB4gDbiAapurbEAyFphmBchJznPhoHV7KLgfEEzENKwzJ9Vnz2P
DYgNGAApNfsd7zI/mfxWTl+bqLd08izIdj2ellS7EOi8pAe5L/yhU9ydMXgDeRwLStp9KacZgrU8
84n+7leV4sYh3gKpuvnE2IVPUc78SxfCvweeME7I6216gElpqXLB4NwOxKYWG2SyM5EjO3b9QtgY
c2oqeZCeoPhKUro+A+hF2GpVxU259Pqyguu2dPwT67e+8HdPvfMpQW/WP5I8rd4IzMSydQDNKf1T
XGt55Gb0s6MM9yteOcqB//ANsTKx0rTWmwf11NrXHoJjKgo8+VtKYxFXIKF/i0Q7zpmeWmqwEgBW
sdEdC1gupSrNtPv1SFW65AG81dTy0jkeYl68jl0sytIp3W8+VYYtyUmxaO9+DhEC2glpCmQdOKIT
oSINwUmSw+fxOk89hnzegUI8PVEIm0FTZBNIffin9dPs/eNv+ZQlsIeXlH0IFyqY9PmbBRLe1IPb
Ijplv3sIgCtpMIbbWQAS7RDdBquLx817wymoLvWY3CGTgIoFo/kC8zvPOHAuAMjzPip8vwqBbBsL
yJt8pIJ7ykkH2B0YTE50zSqxb/A9XIBQMCzlAvr8knTjqVMZ9UcavXwmG55lD/Hf1GdI/DNKV1RJ
7b8SsYT0FckeQsjjP1a4KUvKCvZZI4/hniC204gZ+4+96enLD8kjUjkWBBuA2nj+crlmJ2dVi5/p
QslmS824kaaMw2qQ7efrJ2SGtbuQHc9iV4+Us25e9fUL8hX6vvMWxL9VJF0qfAKOWMG3+5zTlOUr
tYUBnYsS2XgMb3wZb7T45Y6fstbmLLgcpvkfkUhXQuXA2A0B8C8tC92XF/tX0B49PcJHswfh7QAh
h2Ao+lBhZtXeLL3Cs3rBlxvPevY5hjsqrPHQl9BLyvEWqFD63bdZzPrZYgh2W4yhHEzjdI+2lm3T
7smM6S9e8hSR/4ltfjThXgckzqOjz2r7I5Tw6k2PfAuDjRpVqrZY5dmCI0bzzFO3uk/wna9Rl+ds
FLB/uuOrmk/EK8+nBD1Tt7o9vbrA3a7qwJPHkZTrO34EZdsPbFZd9KPjQyTo0u2eZkJUggdEr5cx
dP4l1QsN1aeF78znkngMjWOFn7Xf1bBsAOW3pOMkt9jAzK1GKibExLJZT6dD0YVVsxtbH8acOw+Z
h+ASXtbRbjXsVX3h1R6HEIymsxpE6Z+Pvs6vH/JJ7zqCFBmdylKEbomfL4Mh4sHGHkLCK589mUTh
gXI/ycgtyQgE2e00JLceqiZte/yjkENzZP+lKkpP5eUkXQvxSj8+dTJwdxVZFJk1OpwefX2vxWR6
KWjR3S4QEU+XTZg8LSYmx1JguturwcunIddX4hCRoihQsNKQ2wyAe//1rqBkfQ9gwkCYzrbByES0
z6q8Y8lC+xEqt1f0AoxJuSDtFBHVqPBZo14NHLDA+mnVWZlH4ErF9+fOdVzAhiPtOmAdPdmHXQy0
sK1vJ8Go9gGep251BLAGvDv8jNe8WHO+3AqpZijhlPbbrzyp1MJdICGqsZnsKh+EK0Oxsd4Nxvix
m5jpzIwqMQ6eHk/6uSd2ezS7n21QGUfMccoBIgAa7aVk64fr7o6GduJoUnltqQ2aF8ochPW3VN8C
BVhCdUCLLfFSr1BvrxQjNc9tXZl1FMca5b/0dxnP3ZWMHNTtLS3UBdGa7dD1MPdgcD8qQorx+hvk
iBkzKKaGQssSvZtHMzR11nCQ9+UMbxT3Te3L7QhoA1xUbNOBOyp9iW6PNcoQB+QoYNbURSOdcHS9
QihSHD/O1kCBKQ+dp1c5eiiq0xH7DW8OQnIMoHQjeFvyYrtUh+yKLeXlysspw3Y7F2W42FWfro4T
w4QgrTTDiAaodXVqzrFauEurq0j6MYjOXVay6KIXvPvaLS/FQoHFuS2IJt4RR/fvOxYZEzrYWEcH
IDb2QOEUwNUGdHUvftWGMsi2MlyFWpmwc1QToNlr6V1Nz8FuLKmVs6Sup7t6lEjHeiI56I4oHOlz
wkX/lLBy02nIk9+I0r4fnEdAxdlfvS6Pg+K878XMRTqcuifhdnYsDjex01r+zytWsD+Qfp+/0eeg
AY90wb5lMRwV4J/hGv9yJ2mwT50Km0M9HcYkZlpnu8lVi6W6NmGvv8JaEZp6mkL+YVsav2lwpnC5
2/Wezqe0D8ngwpn4CpKowsR0xJtavn4D2me67i1RB4AXcFtC7IX/gXLqz03k+ShMBUvCG0YF3Y+e
JhthOwmBTNaEXCc3LE+2BoHvLIHU6d1yJTywxCvpLI5J09DnyTqS7Jn2Z4tgqWMtC1mvpHwpThzw
MZoJpO+zXZl/NrQMw2FXBoC3EHCchpPavVEmcTbwM3UuixPpt/gv5Ra4VohEi52BewBOab5Uiz1H
9/SmI1OXwKGzL89iot8h3gyte3IJd71v8ugwmXTwwfPU2niHnBIYypqxRjyVlyk6YEH8wcjS78Vn
WfM2EfILNlM2XOpA57rSsN6S+GpDXsnRsV6BjVv1xbfVh8GbAr+SVyv6RWxn8lvIGlxrLW2Eo/ln
8V1/HqGNw7QtxxkGR76/G8vBNui0tlALXZwp71XKvuBMwY7/fDWM9pJ+xEtcqI3AP7WUJ9DiF+fP
r43PowgPSCPswtvLiVeI54d4EGGfrQWsESkjiKLZOM1/fA5qBwEKvSyVR/tpThtPonT11J8995Ws
HaWaK1oQQg25c7h3l86tR7s7g8f6PYaJEvu6uvTNsR7gZ11rR0tu9G3wmaJ0WVX1Jj5x7ZlV4dsg
dX5jUfVQEJY9+xwZaj0UbKVsNKmu50KsgYPpTI0Fod2qJX5Uaunr5muoMDW4irG0gvRAn6r6+8B8
bYY3qQx2pidpW84wjeBLIGd4vOyZfi38/bEvej9Oa9y+QbwGgwJN5zTkQaWR8AZ0VUw6AVZDV9wq
dfVRoTq3cVb4LYxXZ4utlfVYPzNpd3wqGaykdMkwg/c6ueFTjmCwhIM5RZiSaSvFlJx5+SWLAqZx
Erh8J2MRhF62xxN/X6DV7MXRg11dnXbWQXVCSwAaYif8iHzKsiwofI2KMk06ZaVhn47CyXTfa3ZR
DPA9XVKdk/YUSA/3iVxoi0sBZjWsuAnQMfXjVpKxDo1Gce+1O17mQ+oQ7tyB2a2Gk6uE/6D3rBUC
FlaJPThzEhqdJWTN0OMqAvx0Of+jsh812BoW0OjHO12hcsXKcuCGk2ZTTT2ADbzw9CXJXdjmhrXK
RM/gI6MSUg9cq6xPVa9Roap7fHLN9iG+zVTvpoGadNfyzVDLgh88ZfM7Wc9IIcse8YCpKDpgKV5z
R7MWsPSIm8pXy5p+pvFWUKBzmg2q2eVkdyqNy7M+R39Z56Z2RpgpQHUA2kzq65vV9/cgwz5ropjw
cLddG5P4WMOJ0eG5OJUvQUgc2r2ukWY3+yqAh67K4nrnIofOwZERIXwM9iHxVH3fPN0eD9rVc5Gj
beenCkbR8HQDHuenMrJmXgzlV7jPUWUXj6zK4ULS8T7XmeWXUmE2IR4Nx3Gsaf8x4RsF1D+h1N99
gESJeIaFmx9W5hftAL3zMf2osZyU5bb0CmxB1mGG3TxMosYWCTJuq9Kr55mqEQIwdWd0T6R33RnW
FNxrNnGNc4STE8z1UMrcBeRXUQTa85YUmCoTRliPOIMMq5Ers4yw9JGYdQswoOCSdh6Hjl1Vxb3z
RjA2oYvLXFT82K+Xu7W15yWWXCX9acTkY5FKR++HVhvN48VisBjKdqq5Co7ZtAuKLCr/+4mcQkkV
YnARVOscsHpRZSjydEs5UomRoOvL1a4KbMsUHbDrfx6k89CnsdiVXn1S/lmpu1HoqBUpYU9bjClx
SNMQHy61xg2s7Z+EAR1mTjzV4ZmCGs2gPt2QFQ5sX370Ni1lf73Wmy6zKJyI00SDLGyAliheNRBL
mvpJaBGNennfFbjkPdXKkMbRBV75hMAaHgqK6FVVKG+Ozemmvtoe6lIJUAJsEy7+oCy/XqVQO1bp
4qcSFSqAU5WBDPFEU2P1XDPtHnK8i4QBZN3LpkpHnvZJedgleuggsVYYgm30SMraiCm1Gkh8GT7F
cZ6VuvVpbho7AGmChoLTzMjd3PHFT0QiEKL87Cocq2uc0f6b4ovtyTq/0MSGcl1qoJyggbg4xAzw
0VD8AE2wHdUSfUCwGjIj7I31reJW5F0M3dllOJeKN3Cz0n57v791lLjH7q5R1W4i1GflTwwA/n8j
UXmp/KQ/CN16tEWw+O80jpl+wAQVFfoO6c7GF5WYHXfe0jdkzk1cLqk6yoqspzMxEQn2bMRuUPoe
8taou2rdqwPpTX/RkBTxFJ30ugHoj9B3wN73m3uHa1I4Os876DLwDjDpiNTkl2TVZ9wbjtsYyIAA
5ee6uE8e2/R1to/epCM1+v9zvxJWBbXgDkSHu3YoBg0eiE/iSykGSuCExDhhm0LjDlswdI7yFB8D
mvPa0SV42sVozf7OUraapZtcQeFm8NBzYHcRymU6fNmVZIn3hHXP7nf8GA1gX/mCK4WldUmEYzh9
eVPCVXjXQOI5Pmuh315ueQI2v8PoPLjGgIPd8fq5QBGih1AsV1BVPikqwFvr4F2ylLJx3BHbGg/+
zU8ZKiyvs3CRw34BOc/YcC0uTiPKN+xRMobn7kuehGYvTZqxvyHLXTceG8K77NPmF5KEL8lq2Rzs
Q3c78vRpDbvYsrGcNOQtWnB76UXlKtrqOVqU6VfEDO/6fOWcysPx4/goC+Ip7G/Pnpn2BprYOJjH
JFxsmAuhxlD94IfbrZLPTeyYupIBPi/pwRgcPaPC4lj2vlFw5gimkgZGYAum1BGD4mTPdzioIOSs
msKYq4Zrcb0t39xVJg45Pkasvkawxi9djDftDi10gOLunWsTfYDc/TyvGDrbPCQDMjppSXvcRyhL
QvwuWe6RMXAyRGWMYCYNcehC68Kcxhii7u2VzOB0aPNRY+TjJJOBK+oxdpeSklj4McMOjiIoFC6t
smjWaFhx24qfKMVDf5ZTcHga5vuEy2TYgB0ABLL85x/P0rjpFRXnLc+YZFszmEoS81ufJvFZdQDk
xk8DXfEPaecD8RfXK/mIy68WTZt3uAt1I7sPczBMLv5oz08arbgUQuwh1WJahHsxN9zI1z3dURXE
u1e4tQwtozMqWXx+y2+gcpSPmxl7mOPxxFfqyA0J43KsgKcVtYwHplVcqTZGcZGMi0PM2+B3lAuu
80AmaqbZGrvAg+3x0bTqWgQshMpIBcqTpkG3yb0RzFTKihd1f5J7tkW2LpiFt+tTXgC0wlZbhkFR
t94JFsrsMo8yPdZgz1bMAGPOLWF3PVl7gq+MxosMN8kjgbopzT+zoTPYmXFGs4/BwqUvFr9TKjNH
5cdNX32K1ppd9xLKobBLX99h1QI1r2LEGIDUGEjkahxFhNgXMloDyNbQFlPEbglyNFkIqva6qRK7
Lks1sOkdIXoGVTpl+S+b+0BC/gNMpRtijt13V2Z3CcIPmu8RCNEWy/U1eiHUc6NTNB+9eAjYgv3k
f/1Eu9pLwC1z+O9VncnBR9P/JwtZIwGU5zYoPKoRnjPmg2CiWA7WVzSdx2GRMTZK/xIVrNLpWy93
RNn1df8L/84KLHLSZK1XRSHwTTfXgAmSgzyzN2GtCQHZYsIgTKZJMxNAZv9MeSoAlIhHo4dqwKp7
sya+p9ggk9WfnlW81pPd3WjSnzaRit1xxqrQj1bUG+ZfQmo2AaLn1CjKMyXQWJj7NXVmdMWZZBk1
88x+z/uexoxe/2QoWhBl9yHndQJVEyPl1nnrevgQ/3/CFR36DxMWVH1CuvtJhPgaFMD9u9lFD4Cm
tOIXlADPF0kD46M8zhbNHJPE5snQmWgAwRMYk4qFx/nvmgvqyWJZRrip0Zs6yMcgS6m165NJrzip
jHNNnTpP5vfOAdYchI9pBZUMBFbUcxYEfH/5jpfTuhLRH3GcB0Be0x6KXK5FC+nPI3iEMPMSivKr
4J8r7WOE4fOpj8SIzxMx26V6Sz0HbbG/H/FCpNdjVzPGhJSgosdJLhq15C6ttJtG+oFeSofVuizN
lKOrKxB7Vl+JVXX3BWdbjgoRYOWpJ+x+xOq/HvS7HHJxXYf4HWuHNSLbiA/KxHUyzZ5AXAF0OEyd
TfxFAdvfjKJSRzYmQTxHBJ8r5dQX8XEtL9jCMOqbqUrXbcWmhxOIGX+hcyF2/WKjxJ3AXyCVbxxz
LQNqQbFyTwTtwHZWgw/l1L1cGzt6CqxUy/Hpaub1MNO7kbYTgRMmimQrU4ooywpYJe6yakxuCMmH
+cKUV8JeG9RZaSI8RaVvx/w+BtrIa4VrIaA2nBf7U5RTcr+NK8nLAezkLP5N7WodOCvoXkoUmg5/
jjAwmRKSc7rCjedQC84RfuztJj1PYi34H+v72mOj7VBo3Luvddp52lUt9wbfuRxbsDl75yqwK34w
t2uiWN+h5e3byVDNFjqsUzWvXFGvjKTClDt43jX/uN896WVf/gvA8RVFxUYQS4pDo089P/fpXOXv
8fc5HkHho9sYN3VGU37//lkfOhgp9b32NSQgT8iQn2W8eh7z0NjRt0Haui3PChU1VsHYuntaf5j6
LezfkDK3TcvKtXSUOyV4H/juSNOTri4xzWsEzH2WsPA1ASnv2p3HHJMnNMUcw+KYCkTeuQJ5f2tp
ZVYQNYBA6S66Ia4t7Apb7GcKAog0bZMtNRyef68Ug9M4S9PorrqMFkNYYdkDk1mpG+kKH3ENvQDM
hwmI/8Riu0wSUA3OtyOOBWV8Irh9WlPOOGu757lFNMkv7cukZba/zmLd9aWn2dHKSJa/nt4qEeCz
+QqupdFGgp9WykkOd4bSYG+2obbE+YXo3u8iFFvLkAoyJHfJ2dbEXRI25xQ05W8FxMnTu+WxRAMS
d22lXKFddNYMjExxTfvPVPFfVWV1NKfT98Jlb8Sd3Rx2iQzEvY+Og4lWtOaxB4Rs/RHRNR7Crjzv
PtzH1i3W0sdbPJNGZ0ze0ne1kH9VcEya8gcXcMnloc29EKEXMUk9r/kKewKecHvM+knNuE3U5JsF
wryRLTAvYNDibO5f6x3vnXq/eGZ08nzdPH/SR/8rKr0d7gS7yEaBv+zYu20XmpuPRyoDJYilWpJm
TIkxA6VTgEbHKaomE02CGooxUZ0yJkkwQHdEzXTTkn1WN+Biby2/KVBdl+1RlbmgI3BK55YjZ06N
CpJGd2+hj6CI40MZ1385kardF7B6NHp6tPl1QgWoSNdDe51qTzTRhfZv+JqpohH9gdVRbB8nixmZ
Qdu7nBgg2Fd067QEAIU/IqJzwXoupyWN2PamEoz3ak7bBE6SWqZG1QymS8UJUIJQRZlNfeDsJmFr
kRbvrksXju8MLRwt/MyL2Dq1gQHXPIDh6HeHTsXGKGhgkw3yxmCWj5p1xPXv6YPsWaBBAW0X8Qln
gHfbkXSGxNnErIV+RmYKYQOK0ddUo657mOHamQiMY1NKzAm25FKRslhnEgN32WCd5W3YHvWzMWjx
JqSpk6MLz9rNVj3c6ekUEahI/+q5gYgNAyrUR9lyH2rKwsopyTFrKqzR3If/iBTD386xFl8x7DfT
sDH5Anvh2NKioArgfC8JDVyHYL3CLyjr0YhP/Mo7bGKTHJXu2FOyeDzO+jV4nm5NIb8peO1SJBJb
J0HQY/eCpq9xyqNWuzyyHLTJc8lo10lbgyz77AnnsahrIwsyBuOWZD6ZvoXPaxpTUkGyXrv2Mu72
VLddtQCYIjFCwmcAJdaNeh4s2KHhJHkO4d1ZV3M37NN1LmgTRRof1ixOTTU8DNYTlPElNQpJbgiM
55AdGQGl8/KqqpBh6PjlokcbJA+DX/NCPeHt+tglyX+b8kPzfr3QcBHkrlMGWhc80jIMgAAKBOQO
EKPkrGKn8N0nGzSNrbkMEGlaOBWdysKsfc5dX7SrdQJqkq1+78iR2VZOKoIW3/9V3fpeXPBVmXYB
HVbqk7XeAyPgKBzEEijH8aIRpCXHhY2UCVTM0Qvnu31Y9I0ZcCV9DYwvQvWIrJHAVIucVo23zmdW
vvgOPOo8FhSZ81NE/vHqatioJLByU2bR5IXlMKwr0wF8JAdEBo5Erjp1qeGahg6PcPEcKuN9LSy+
W19iM5VTWLe0Z1qY2HhvNOCbg5uACxLT24XB2zqnHO2L6k5PfyrsPRalzq+ZdBKEwnY8VeoPcSpc
lkR4a5J5d38kwmHLlVEousDroWH8ebiWxhyBeWtgwzecRGW9F/5ecwoBlv3I7zOri1ktndzY0zom
SzatCbEux+D2ALdPeaC21+wK3m8s/vjp2GrN/2iNlOBYkMUrPBwDiiZAKHpFSzZ/Xre2KiZxtLg3
H5zBZ4XOuBhcpv1LJW8IxSgh8GLIld75KbC15dEeJ+IH4MOWTrgY5NgaXQpCwroHdJo34+0NvCos
2Y2U/D+zYp41iGiCSonU5428ZOJBETsq5YP82+pscZgBwuK8Hl5+A4uOxp1R6q4MXLlxVW4GIxX3
WuODEMzvNeuUTDmDTewy2TiM9l+x7EsiePE4S+VTZAAVVBr3l7MNVaFtUViPjMdJ7d5aaQFQf4gb
i0eXk8EoKyOD/Cn0hSYbiWGrzZjUgSX0RbQFkCTcTKy9SijAuGheU2sY1w8ieCs/V6Q+YxG2qbcp
geQXzggDEVwnKCcHToxlX/0PJ1Is0lHM0Dbfiu+pkQ8eFzE/FI0f+kvbek+H9oZHGbYoLLCEVxNg
IXFxfb85t43gdEMpBW297B1hybZVVQfHRUOQ4SPM4SfmDSylTBM8ujjcVwcSBf+IPxy0HaP9Gp/Y
2VGkMc1/9pINUl+npbwBN5NW5jk0FxHXUsg0rhxprQOvm5bQYeZWZ/nVOXwep6oO2ROyjwBF/duE
Zc00lKOiIDsVxRGPVs1R+R+cYnbmR4XmqT9caz/uwP2P7NDL6Uw0MP5Unjt6DsdYhGS11guLMVfv
t9spbLG48SBuoNVKK4cZmWNJLJg6mWChn6OqS16uN7Y0G7whJOOrDNEXpH6bLjIVo31w1PRgBh1v
nzIIpde0XXXNPszO4BFhFydMggd6XSaGpfyGNiF4Ov4K//vi8jfYv4kkpzuzjjclGWr1vZWgxVpP
jXnxWk2W38+dYjuX2wjW7y3XaV3I2ORpHj+qq8ot+kMJ2mCrUhdg0vcM9rDGiXjyuDBIUhK2Q2rR
aOHiQ+jdU0S6KpFHM47H7LopIm9JHzm+Jczu99zHoN9KJ3UAU++XRNG85goRz7j6q/YtAxrfpEgv
1FtutXu/MRmHSzdgrbFmweh4meqH374Hl676T9/XV932E0RmAm+wLNXmMWsel3+TwL/u6CRfJLQ5
J0PdmFnkCWPXmKadC1PcISCN8KYa9DfY0uCcl2OUAJkkUzmGKlHRFm/HipUS0ZXP/iD1tRv6v7EQ
iE50VOnLJIWFnE69nmLRIztqEloZaw0KTHnrn6s87HuZAbaIp2A/1D49/IiGRSrjcTQsZZ96skOD
50mwvcBdU90S85DvSBA+iHRnGB/iAeuPV+EWXhuJA3XogMOK6oy/miYfu1TKy24Kk5XEY90lrjSc
loFB4ANGhKaxeHvR+2pH5JpmzxtKiUjxaYnJRWP9nTedzQt2sFlHosTtuw0YfrCdjsHTuhOfxaXJ
UERWVMIXnDCqfA8MQgv6u4lGGNO3feTrR0gR0FP+QttSK9GXdCyqZVfEATtMoC6MLv+NNCIel6Ck
VhXZIirLvnH1Jt8nIZuB3NCHatzaOTeJ00U7xKi9mcUOYSnXswZrijjxIJtJmCuTrDdfXnDPoaA7
U8dreWBpEtrC2WoKtIcyjv79bjcDUOSGkb6zmZmSF+IBrabmzZwWJAO4KZYe0+Y01MHqICC6CmOG
+LV21fgZYz2pEA2nMFbR0jfdiFAWVo8g5pagUi+9JGV82GU8Spj2qh3Ce0MDmNyJaEARMLLrFl6d
/vKI/vUu6udsIWGSr8U3LGpCOWLem42ty1jkkYxWTocaUAEAqPAt0hX0aQwtUxldjjSVcNSjMe5w
7HX3yw2ts0BdminvbTbMFjFwJtsGQAfK47d2WVY13sEaU2z+jJU5cOdaczs3Wvqd4qIsE1Qlds1i
49AAPILfF/0ua8YLcTctN3V4/R6emrVOYDpuzxFsNEji7+crScIbpQQSQAPaCf1N9yjAVZCIkWHh
wMYlFiJi+NaP8v9KjB+I6078mlFNxhQk6JOZJ69zbdQvFf4TRUSVvUvcr+gfRvNsDFtJuvFjEjm6
rsp9Epu7Tpct7Yth3l+X3I3fRseqjXcoWfXmkiwgqDB+3wQQpZ5cxPH2l1ozfzkLEYA7SRJCiNEQ
QufEXMONOcpA/bBkwrBu/tq2GWUOJnCV+FK5NjgFeO7yNL59rsc2nc6tWPjhzl2WbcX7We2qZy3T
JZAg8JjnXN3ko1EtI4zhH3uPctnXbwV6mkzLbRj3GIKgM8B7HtIyv4X0FMR1xek9Y6Y7rV2gPK1M
kb5oWdFqL2rlUqMNSEsLVsCebqGdLL7CzCAgsS9s+tsGJAHnT51oDd8HDpeYG07siOUqVJ3GbwTU
ihh5W2TqQ3/XQSW6x+DRx+iNPewn1ekiNXW/63/OIHaTCSpdvUjNCOcBbuZBDNiK3sbSmPrsEXoR
maj4sDRMwiAGYEuQrziPVHp5OmBXgRB+M9tM2mTrhBCD6tzon2jkNOoajbCZq+AQBH51SFO3vQNh
qlnSsxLCUdZiaLm/NOW/q8VcDqxP2jsMc+WluEbCVrkDPjzFycxFNjrYx0ZNYiEDHVpjDDOOS1Hh
6uZQQm5JTUHeyiFh1hn01wNyss1OJo2cDhxwz6es44Kt5erjVGrMlRC9HkNTA+dizteAwe4IU8tg
TKCrAGV/Pdo7qh+yjb+wfgfYV8y6grsa61lkgXJ0QOOnVadsveucVNFrcmwZpOU8zbpHrZZDCJO9
jt00GAd85idq4UKdazwsXv5rhV3tyhgsAW3YlKyASCFCfLx/FTrAZBOOyxp6H7Gkgo25ft0ht2cE
rk7S1hvhaZzIEvUm6aT0mWd6ItOGzLxLl0+HtLUaHV7X3l0HvcMSt+Yak092eO+VD4yWkZcNj8Db
dCtilfeD/h0c2k612KVx6kwrVvmUG9za4+sqjTW7MuKa8/V1OlTptAynxJQB73yW/y2qxq2Wuq3l
U3X5HKpOV09l8B7kx8MX1m/I+NOYh8lWYKn/8PFk85P5PykIbcUumnqiilIOr/FSOoVXPlmNTrqz
4IWQCfQM7BFOf875Rw1Ex13ZDO31YzA0NtOPNQqiIaalgejdZhEBPx05CyrKtGwD9xpirrWuodv0
PAevG7pvpjbgG1+roSeS3XTtnKS2W48QKEpu0SkmkijDCOZyp6gQdMNgxvSWhcrl2GI3wiEd5a2Y
NshWXPF2EjOsCOST4CQ8tqPM930EcuFOm5HjawedS5mLADbVG1BagU73aVGOw101BtjXrwwH35xX
xbfob1XlV3iv4L88Cl0qhBZt6PByuW8+ck+fuhVEKw+2eD0249ne514JmRO0LksRtWU1oXdroUGI
jvk+Oth9hRvUsDcum+21foVIUmkOQ8noboXKssq9CGwrNcqfutDGdOgwRA88waIwaT/zsxyIs3J2
UdSl6rw+4EmxOhK/fPHAuI2/x7SCfuJS1rci05DhDETTlnxGqWJzMsIiBfH3fv8bYAdeEhP87twm
fYnTywpposgZlXD635rSeBgJQHrfIZ+I694i7kEjAJwnL4EnidwMXhZ4s/2lzbtpfFKqYg/fLp9W
jC9E08N/F9TRpdf1WJLYj4UsnbQCUCS/+CI563S/Ou5jIkpUTwCTPgc/TF5kPcpmXhIOoEmogDZA
oPZMbRBZ2i2lsH+VIDuLzFx3f2iK7kMi8gL4g1+4rsHMRN9FsgtmG5TBMgjUXf4sW31WwloN2adJ
W+uOaPSN1gqJt9gzFrO8szdH+mgoTa+WHbht/2Jt5Bw+69r5GzyWOlj7cNcZSbhrheqvKrKHIQmr
D6q2vsCp6wpphAhT2oLT43WTawe7wXcrjtlo9hT4Psns2ZJzMB8f9yqEN5d0BCrDSE+Can4BPK6U
zkGAzfOAns0gL6gGqrig4GxiGrNo4FHYpKWsV1JdaYiEQFrQtkvXRkJ7OvpM36d50ROWcCfmIyRJ
pVPj7HVshsa5SHD+KH2H5UhTsUvGUqVRl4qbehaRaE+CZYh3xJsBLER3vZ4lgSrPacsWJXXv0mN8
oeKK93ZhUH7pqjpPB9p5fxh0cNMHxOtVpOJpqzOqd+0UBT1pqG2cxy5NXQW1AcDEDPQCw23vQoUz
RAE4ZLiTqkje69C4bMHuDc2vfnL4adDwyEsCK8BKZ19GVAQQwJoeqdWGQjCLWw/0pkpULf9nZ1Ta
n/bjI+mn/huAC9s5kLf2Yra3GhgPLHhK1MsEvA5YoAb94huyRFEcnu3X2c5JNNpjvkKVw7s0AyKn
bVSJtyF6sxJ3WOknCQDv9FKV5UydChhe6Xme8o2uf2SKwzzAThy6u+PRgUpJsfKoL5XHS1I51qGM
FyXfUnhgtEywVomnrtNfF5WvwN/j41NTZoOGWd9Pft6ZXarNSReeT2PbdMLIb7ZqGY4Zw+jgBySX
mTOjxkmrvr2AKVKPXrPqeYKvepA3lLlHUQYr1Ua5x8f5FKhtBku7E9JeQAl36/UsMqRjtfw97bgq
wyPGxwbXTDYTVcldt6KZQ69jbdYxQ0Jk3LJXRZZvbfZjU88Xq9h6D8orlaHDWlpXcFIhq721SBTV
P6VcZw6kZeDUVyHdUhzwUNG1/AtDh8aECiNyrdee9uaFbqvdmCK7wi1qVNMRdNx+d39h21D0/Cpl
7NSoW+WFHuweBBITBp2ip4dLHz1qVUt/aKj9YywE3c3gL7GrzhtcGMvZBkT6cfn6zko5pQxmf6Wm
6nQuT6Fnxtx0CiecIKs/CGU5W/IlMK7p4/d+qfnTUJQpzSeDS4BqXh0W3erZWm4xLNOVpDQNabi+
64IujDI+B9CzPh8HsiY2nqKspu4apWStgcJ7uaOlPrjEQbvJ3TPGW79jb6PSxnovR+so6wz154IW
LD1wxkSsYskNTxy1rlkTZ5bEMNOQfjfZ7hXPkYnRPrLveUXpG/vhwhtWwiEftqLgBQPYBcRbtsqu
1UaDiqApR0Qv58ks7WqhXzwK0999zBg1crZvdJUhyU5QL9MQzeyCosCvYqZh0oLH3DErBbt116fR
bzAsfSodeaK8hwLjILp9EUBqgJJO0mwj2/NwuivCM6tdsa50ovxC3VZSs/zVVUftoq8xm02oWmjC
pQTDerzTB5rZPx3ERw/Kn+0li2OrgOwMKkyBsrE3TQTKlBGxsgKZ1aggQAJspWFM/Vn8az5ltFQp
kW2sXxiPvvr/cURwoN8rudb18isIO4oFaWqm8Fwwtv+CAXU05hsEPQjD/e+80/UPGx+kzipgstpn
w4YHJZO6HFR4Q8PrsVWYI7Waq5jg+n1jw4n6332xA/26/WE3J71/npyIndx614mptCpa3p7YnvqM
uVlSi1meV+tVYOhjqzc8aDWkRrF518I2aIQxOJVGbz0fdS3knBnn990jXaz2HCjbHqyXJA8lkkH+
1yX2A0GIp5pb6i0JWoZnXfk+5MtYyS7wjZx7H/36qVB7NK6IDEh19nsSxr3/+zPE9DnKyqquvUPW
SB2Pg9FGvL2/UdM7Q2Wgc3BOj+PKAAgB/BwSr/HHmcSnoOisSmkGM5CG7JN4IGhqEnLvOGrVv9dq
ktMhcqJhqRxM1aaD97gx/BuMkgw63NNqBFGm4Uh0vzlHrVQPgceJku/Ec/wq80IpEp/YpRK/dgl9
rFscKD2h1jDunOXhA9jW06UlOOECZgO3QJkJGnMlpgIo7vouRqzNA5T/jNIFNLKsqe0596iyjW0o
p7VSPYhqZr2rxvZX4uR9nuCDHatFUxyAsbCIOXY5eq43nGgz4++DePfDVXN5n6Uv3pYXY6cNadmM
CSKUUJ8bBdzgNCJ5WDSgYu/B/FRvIifcZsCM+9CpCfJhqN7l5z9TdOCAAtC2zCpDcBlLdXoYbwce
rUk3/leH9wjtyuEVk/oVYD4rnl5VRynCnqARwrDFGDv47Jgon5WznjGYSsctt0490wg6B1nGlJ8y
KqrVHFtFwUGXvZXTN8tDmmR5BVswUFwY/DI9mzfBSNfN7MM0hBi4NJKayMDZiR+StZJuZ9jnIqTB
1YEUr8eIGbhPUqwtOTy2rnndKgEsk7I4744EhcHYgFkwtJRlZiZC1LR6k/+mJPlg16KbwH2WKo22
Q/H76IUPvdBOl0LT2vYam8mWNV/gNTYxZa57mykdYyWue0j694u7HI+ToDfLvfPK3FdMkAuQ14+Y
J6sGXZE90ha2wXtx2P4LqyUSrsuBEVmHhNZkjXnA3usDEXnoh++RzbjnSUogyJ19ku3tOcJp1pd4
Ff0xC43Q/vIGTtTVi5vT87PuO1B4gqFHhV5gSDj45SsRQVgYBDee8OHdiXUvTsHvfm6SsB/VMTo6
kM43KuXYUkDfdugNZClO3JYLGrtqQAK3llNgWAGk6Wq630HiaA2ZcM2UwKfgMu337/73HMfKaSm2
PdkdiCKayXt3nY77o47/cj3dqpZNkNi6KIufGp80+4MakFcybfao3R41LURw9B+ne2d1KcW/t9Gr
QxdPMKZkn+H3CfAhfwf5lgFuy2P/Abn1B6va06b08tMuMEp83QHCzF0cGVDXpxbd9uSOWraI/pp8
ZzpW5nmDlieBslW2OZ++TqJMcLogFiA0b02Ohzr6AT1vdajxDcnmQmFTSiyazAiRorjb6dCRXgKz
XwsQVJVwWG4YN8yMnx8VLGdBewIPy4aN15PztJ1URsYNCmLR3NPskWHovjoWvIKj5iA4yRcNyVqi
9BnaKwHoKuhQEly2HtV7r/SSI/SpW1JI7Jjc7UOUqEoNPChhdPxwBM10+veH3uM9DEb0v6PE7MMT
cyNEymlSoX/JlCoJp9HQFUq9shWgErn6Ckl95hngwGPVfGEdh2/NstBI7vyZSVk2MZSehcSVaL5C
48TFa17gvoWDwrBSQ33zh5ZNeY60bcD+f9ERl9MrO9s1cGu571h4Dzo7IAFrB4J5MS124uHuktCF
pKskVyfAWPEQoR501j5j/8FnfieMbjrc0909NEspLWuoCUHLayU0xqCUyvEuljFttuiDDl/gMdE3
BmAodPuResiswyEEziSlhMJIyEUHuAeW0WE1v89rPvnbLJPLSDBDl5totbZI1UK8XrJ2hExIhtJc
l6r3eFgGORGeZV/zGZVcoZ1QC2vqea5SAMe+5+hFm69t2f85XCqqh+tiVzXPdvCAZa9Epl7xx5by
mj6OBirP7OAkwkaUssvjFm9KOWKnl92S/beWhWBdUXQXbKlveon4JYOgoxvoFyFPq+jOlqCBaxdp
uBm+51vzJ+x9j1QBxOthbarC09PDhoZ+q+VY/I+lY40pwFYq7XYnkIz2Nmse1eLiQ/SGWEqXOhZH
DvgxLQ1k5S61vK9Ee6sb/pSn2D+xu6/+kRl2LcZAJ9FgN8RBXZIOv5aZzuAPH5DHKlQ5Pj3kpkk+
WOtW0RMLOo3g2b4OU7K9ksEvZGXkp2jvvAj7oWKs47izk5imSK5cVJaJkKyuGpPWdOeXW860/83v
SVoT9WQNDzUBqOL/4UZ/u8gmkygVyHJqlvBQe4Z+bDu8tJ4ZyLJIIGG6WAu/71/y+kqfMN7qS/Ir
VCMY8pGXtUBEuHQ2y1/+ltgzEeTIM7zamiQLI8nXE1j6W/32kU3nD56SlwTPHYeCv3KCWzFq8XyI
svDPOMF/9R5GV0ba+/Gs/Z/f7pgLTQkuDOc7AOQKvFmynqBgIfdzMYA+Y7oCnDxQyEZM3HtqBJTk
AHUz5mRae79XCz+/WPQVWGiaWDjs3gwOtYq+nkSZ7ESo3gESkK9d9ScSzG+wDIi7ZYTC3MMoj0E1
G6IvX0alrkKQNiGXsW8Zkc4mojMJTIXGF/2TpIqVwrqL3ur/LTJUe4mKHE8+PPt3r+fkA7toivO+
2DfNmAQ/Jj/3ToaCxccwJoUfTPxKFrGIkxCrPHH70J6O4gLNL+N/LwHrqq8kgmNXNi40MN2KquC9
e2oJQr6zPqXhWaySnLsr4HkRn0iNsFoGpnBrrO8vbitj1EXYICJHeroO/GOcDuYt2VkNqApywXY6
4KCNWVm5mFM39WOttSyOrjKcA0YHj9FrY3LvK+fkdfwrkQhKwJAzzUV+rr/yhqVgv3Eh0LVk6Fbx
d/3OlxDuPYf9Wl7ftUli+SVgKwhuj1ZxYB/PSyF7nRhUpEHqW+vbxL3lFJV7lBDOoQAaOzHqb+7F
Sq2lAGexlErqAb8bZpNnCV8+NaqvtsiTm1MEVP3ckEu4CjtXu9D65IJHAykY7vuUWijnANk3/R+Q
FIAPmN7I+FrMWi8W1JCEQxfWZQaZsW0H4HrsXraWah2Sp1k+QGZCYD2cPLzRwIKA7XGDNLo5CXyr
reBCXW7D2p+LhNyhWYhnDxGyxti8lTmHKfHXTDlVauSFdovVmDLUwxRtggvKAnjMKcKxseOCE9Nx
2CtxO4p5yrT3OIgocBb5WvG9jP9wGcMeCWY0X97WHH6PEPOjb0MVP5uOMjWsDIxnzhMcW8qsjhl7
g0creod4SVOhs4d62IQtWT/ipGAixi4fczB1A3/643cno1m4yyBxYSfSpyuoGQNqClX+XhtUcCfA
t+2qQh4pOtN7gke6SV3b/0TtRJAbFQAmzhrG1GlPEMLBqWkHqNbZkOhAGLN6+EYmmMHlLxyClff7
+kBlqnrjBpMlghAgNFUoJEljpFdfMvgd/DV0X6q4zkdixt0ojyyRBq6aUsfyt3vNwFbv2mtu1G8d
iN00qxWxKZFmvJ3RBfn4fDRAQT+v1nxfQ1xw7FODwOaDbQapeHogTWEP61+UKLu8bFe5FOV8JCyh
gGQnByvDKxj7W1+axKcFyWeXgsYOOinGWVCumK9y1Bbow5uTAfS/0nuX/lw+t6EzxP5twpQ9FHdC
9H/EC+a+7blUgOMrC9ReHmJzRPcTv4ZBLjFdFOn80WCkgwtWhuyAY03BKNTyqff43N3S/tAK8OZT
YGCxuYUJ0ULm6iNRw227viSuluhby2SNYN0aHKe7SxQIVCNtXNg+6WTsty1W/VEv7q+jpoack2pg
U0AZxeRjD05XDOhr7iJGl/TEhva63DVGdUNRAT5tdQlqJoMyqnyHGcx6H1wedYmuIHLHzEsY0eEe
0Bp+RyQD44lABBZlJWUu2Vsk3H19FyoCIqNAXGlIADHXXabn+yo1KXaGJwfk9+fq9qXkmpDSrtay
UCRK49xpr1/jnXnubWCn7OKnGbWmtye3f/w46Ta+zdV/IeC9lXD6j8P7tpuS7HKvAw5pMrlnWaqk
pSn5AKTMRHnSNzeoNsxZV5m8cWQif9Y+P/mUxS/OH9VjPKyLY4mZwKZ6rt1vHUdkM2fgRM1oUfEr
HQ9b3gdrGaChjpUABd0XDVq8L6j4DnR8YrTSXwm+RcqITOSllwYkRpGpJcabOxjEwrPaoRdASDRB
nMeAekjGUPO8fiU47/no0AaWEb7Kmu55ZsqoMMiygLtUOcFJfD5lIHROQx5u2L6ztBkPIUDkqUBS
MrLv05A07ztEJH7DPpDaOWRhbtXBkybFP16IK8RJRkRueCcosA4xxvWU72aXGtimwMyLZDcOUjIz
3JBDDJg4K4/nkSMSNqylSBQEXlJguPHTP0nyKzKKU1kJ+JLq4mrVI95zMFxm9IlQSu/GB2UHc2Hz
0xur3vKVyeLOQlVM/iwILvVhBppi3zXfYCjbSH8IkFi3aeOoLHWwkdy1aKHq89+2uU4wzHRMrrIh
SRrhR1eoABphGL3plzpA1MTi33MkLm8D8YOuGygt0Q8ydfQjpZf4ox0vy7mfVpuoOXsK//tDjfp3
hIBqbLG663TQpTKGwLtTnRUDmarPQjqSuCenX6kvoHJGu/oHTbqFkFei/I+LpVHqwZAdT3sDs3po
DKjayj7sS/psgNRzs9Ndfoo3J5rnuj5mZUdVACoHZONaqbTlv+v+Bc4rosv8pap06xvS2VLgZ63n
EDgGCeWfS7EYgt7a+38yhfol6JCLrvra32L43i63/rdoSVh9wAB79nPKNcIihTOptZdfHzK5vy3G
V056RNeoh8twirjsZQpVBhzpOOZQcNszfwQMBsDC7XwgXrandeXtmTSYMR/NeOsCu6swlGtKAZJa
g3meP4fcZHQ4y4h1T1ddw0UhsVK6rpLsUI/j0DCdlfLQzYev+0K1Upoq9KTaoLOqfHAna5MhHscJ
qSU2td6iVSUZ2wu0jGHDrpMD0bZ18T2GD80jm39jKVNZjZXeLVKQtCw9jwRpLk8q/sU9OXYZ1sts
Q3XHWpGv0Wi7ofmS6zONYJAmTAuNHYeOkpBsjgyXr3DyB5gKTKMJWWM0L7E6BXMeL3fkzWtfixn2
YMrI9Mu9kAR4KGqoFBftFumTmRun72L2P+zma+KjLwNvaAN1XKoqWcM+Apv7aatbuuY5CEZbS3G9
VxSOeiY7w+VpqzcuMVLGQJ3R8PYPycGuNjFypXAspRsMmaPJOfRRQ/T5cY9JxbOk7L+oZyLwZYzA
EOpypDWYphtCiP/DNPylCf0ySmq7zkintM0Cgr9za9+JdKN4MGmC+NIwRu7hqTuUzfL2y7NF8bcj
WOvFathML7slwHF15extgwJrMNGu8EAH63hvDAa/Wb47h+m13qdnoxXStU41UPHe6cWn+6EDEsgi
+feEeZHnoBGiVe3/ghbiqET7iEekYDjQkKd+FsKcrVx47ITXu8tYxw6/a4HIMO8qmBK3kF/Oo9cz
h6BZ0PHFyItGGc17VXvUDxRHXVp5xJ87a9NQlr687T2/sOVXZfvsIoUCzaF1T43DkMFDI4LkuWkX
EbHOJjrIgL+7YV/XnPXJBixQIblYFh4SNZ2BV7EJieIckOc9mDbbhgrxgGn/tqRYqQlt5Q+Q6/YH
DTI98phAaAjYAv26B4MhoL0a7ssoQW8jBqUXSE477nthrtn0O5dGhyo2pU6TvBwC23xUbnID86Dt
dvpj7bVPAVz/f8E5NTmZ3S6ktoO7fD5lNxdV0b4bdz2Ob7vBK8Aw5UW7IOMgWWE95uzss27iEWPg
+kAVWKat5dgaJgNVT3wgrcLct4dBlDuRk7uP0E+lXKacuB8zOvEQuQuhJ3eDTkY46PFbcnFYwMxZ
jaZfJyVPpmZYsMMKcX3ArONaJJPAVS5U8qHi0HKhNksoXoLcMDzJjvwUhfI9vW8s6tN03zZ74roP
jDkNle1E4HZrYro7HJ+aHlb/zdj1W6HbhP2LHSivZ1Bt72QagFdmqzJ8kjZ4uf/T2NP6MAGrONC+
9IRS0VBHBbvAhAwkV6oWpuBLWPPzZNUM+G6ClS7njdzqNdvJHBTas1r2Ng0rpOAbsYpShPfTY6xJ
F/9kfK2IOyeaMlWphy6M3e7m6EF5ktBtcK0MkoH2AmY4iX5Vy8ZRQrcGz0Qd2Z/PZFhPyig8Y/s7
kO+j+CypdLsRAsJhkwMO1bLRhSUlLrFTJp8egho+x8HFoM4dLIdUUbpRqKwJK43EoH+QZlaTgDii
4tiiBVHJAr2wnExc3/r7CK93Q/2L34pjUOJxnWMiQJjwhmQC4ONL4WXQwb3pi7Cckiv8fL731SPs
J++nHmDkyRp+5cP0FBwlGPQm7tOPEG177P/QwhikD03zwJ5LTtiqfn24SkZgSONJ7c5rwoSZtMMn
fCR4JgQV2R0u1+4WTGytht0UddoUBObQWdNJ925o7132VvRl1iDtsUh5SqKrz94v5RzlWGGl4IxJ
8ZOKAl/pYPgEUjmrsYQhpRSNIp7b2BezDQr+FDoVCnYcdl8i1zbJZJ7cQMOLPU7DU3ZcMPy/G0El
aHsCnDpGpL3g7quPLXtpY56tM0r2em+jaxkkHxmumN/NREqy2aqAxxLi4hz8+Fjc5yYosTpwDq3u
3kzQtiNXMGpfgsTuKzSZ8hZPUIwWROh0a2Xww98AP+o5xd0lArgvcqEAocb+6Pw5rb8SUp/Rh8pz
RMS4sLuKU7hPwcpJUJ07gebvu1NUhTHIZWc0IIyE80ThtBmlc6sqE9EdRz3+207nltN3U0PyIte9
ggQUeuafVSv6gNu7DFN8cKxa8b18Y1xemVjPmoC4H9EeC8/4MGpBnnyni77LmZ1WjFrs8gpvnXb1
mMNKz2mwJd+LxhCR7lGjjwo9T/BA920/9cWTJmMZqPk9PF+avGJuYoqaNmwVGicnsvrQht8ohkam
I3TgywV4psfIB6Sf4bQP/0Lhsp2DUJ6o8hWijFVVksShqEgdwbI6Npc8H0fZMbdmS9xBAO0j97dM
pJDhdD4pObwHuZ6w2/HKk+KPvI6tmsHlfTY0XMezOglK18kaWf7f4obHlj+V1YbH4djA9QmmlWad
d80ZLruVZY0Z+M+dBNbLxCgHf6QI/yE2K+2LCeJ5rfxi/OQFDRMIgIJLi/Gs3L/rabaoJge03teF
SbMx6f1YJKPPrpZ93eWPT9IcGEzJ4yE/3CPpBFn/TkD2GC6fxyUdpKDeKo3jvyVhcO8gv8PpTkoM
wLrt2tN+pi7egLuenZpAi4SkgFZiec9x9VsAg1Ry5XftaV0k33Nxu5IqjxMCitLtra4qO1N6ZgDF
Y8pQJzMjHLWt4/pj5e1dH8aRBrlIBGFRMdtUqKw3corgt+dLce4PB7i3a+RZziAUQAPeWWcZ/zb9
i/eLBxzNVe64e3M7G8YvvEmEd3dG9oPRZYRib3PsIqkOV1QPk6eJMHnk6gUtTFVV4QEYwCFZyyfM
nQk1TaahME7tE087alOTpjzUJOEcVpsxzJMmrl7vX7LqSy3lKjFXKIEKKuCXfbNrTF4LK72KMkOp
jVN+seJSrWStFM+BRUWOE8h4biaHB8RXUSe3qp87rv5Yqjg87RVQtZbnwX/wKz6rHGeYhOLDoE/O
dBIMNWecpauUraw/GxJ6v3A7y3I1uLo26bSTOzJ/HIKuORX8tFbpfJsRfgGT21XjGcKBG08KrbM6
UN39zsfByZPcW2Dk+LXj0vRzMuWwakWUNBri+gOaTsHu832d2zMqY2R9hxNT1xk1/ZJ4yl8IFOHv
EnF2wqpLb+DvQyEcaGbzMjdGjbbDA+J4+M61VJpTFzplYupZKANiQ0BmC4NZ3PR1903GD8neGdZ4
zsYkln19WvJOeEdrcUsy7HI9smhoEdqnkDvXgK4mjbilRxO/y3F96z27WoAYQt7w54HJ9daCuJR6
T467hrNFnOCdkg1+DUsfcLfjFii/soTmkvJs+jkV/gtPM0YrBaXa86sZKo1XoLCM1g0tnJ3KZtfa
ZrVZ4gql7wRykPsFf5u2ryM/A/DfN2Ijh0x261pKZkWFfbYc0UcuERkPv64CwtxBqxMzUoY9MtbE
QWtYxt7lp05CRS8Ywd2DVD3GrIIt65s4bolcNTMebTIvtShE4xZB8aOdbJawu5hO5vlLqYZdKfo8
FCpWAvEeTxlVirZoKpKLatg4FXsEN0p2SNsa0MRBhIK7i4AbeLGyJt8CaLfU8jxhf448h/8M6h1k
+DD5LnR8onGcQHwCQR8HRBAZQaNxv7Tz9AwPHURjRaL8AM/TAcmumB/4J8cN2YL0JqHzSBkBkgWv
9Xpfsa8NoiatwcovbuXMozMxXqc7iEI9L0kmklC6aXLwhTV7ndt2XfaWxkeZ+HQTh59AyGw8M3wp
jiHILeF4j6VqMMKZv/KYPij2ZpYkr13gH+cv18g51X0bE9Ts/dl3EixZVlBJnFM0ybnal7Xl9s4h
7G1w4GYoaRrDyIauuOCzqhefvDtJ1rxCY65h+GjNv/c0pstKKoozkpEG+von6OPCx9m6UJSLkehy
78SrHVzkG3ixm3ikymPenutxFOKCrtGHFqPg7aKNyuNC4PBlN8TSQ6UhHmF4ZkyQu7WyT8wGn55r
+yzTYUutEPqMVHwb7WKG/6fX3P6nt/WE+J++LJqtiYHA7yKJHziWlmcGbDU8O7+j7rldfkjjTz+1
I52QTlSESv36Pg1S4RIC1ncqJC8E8IZq9tfhGy6iMWPGbTPV1bZGIQwQTeywIZ51sahzvli+LuHx
fhf1jdfJ9vpoH+3y4GlIMVEdRvwiTxWqc87JhI/WobvTFgLwBv6JPnW3bEke9iHg+M6FP4U9Qkmw
zAoiCENz06bmRoSGzWDv1cmUTFXYIU8KtIPCkrm/79VkF4gg/GQ6ZNG+yH9ZqOHBU1iAIMzgz5zw
g0VIM6BNH4XRximSwmjpsJ2dToLkiwgzx2ZnO2u9ehkso1ENMaSfuyyXW52h4M8DojnBLpI97ha0
MBHVWsMmRqNjhOUSPX8eXrAC9DLKRzJPbkAVUL2Q0W0BJNBMTMaXDLREutPiD0Le2tTNtWE9SKgi
3/CzvmQkLj8ltIEa8b44OkRJdFFJ5rs0igXjF628z2UW9FOfpmPpzQUT1QoeTVgPcvflgyG1Okrg
BPuRGM3t8ymM3MdhQdtZa8nYeOYnV0Ss0FvhBCwmiSwJp9y7ySncKXFOZU/dj+EsrpzVrtkXoEPE
crN3X9RFEd7Da3Cse+cr2c/9gedNMIeFBnIcCNC8urg85w3LgC5zS3lTj24F7IkKPEgvLuy167fv
wpNuf/egqXAgxaR3b4cUSnb74orgOTxIv8I71g5/FHNtOG5Q0tW2nYfAqYi+jlcD89FBBRXZBG9a
7IpthJabxleLgU7mjCreNsEmPXoXdWCgPagX5T48F/priV1Ask1CkhX+KczIaBkTXNyRsURu/1dy
GsJuOm+M0iaS/vZsFEmOpnHBhK9vu6IbLE67GpHuv2UUUv/ABVjvWBZmZuYqwJ8SHvja1Kny7v8n
GRif4sJPdXRh+OSSWZaWzzhJtT37N9YflxKUaOnWFLTAy1X4eiyyLxf7fNIkXyarhru+TRCKT1+y
rV8zS5M8pmuHSWzR3fBFmIsMb+su7chKeIcEIG7JLhMzXa9GYTbgeXDvE1IlyqQtKVhYMo92AdT2
7CthjxcwAB1TJxcEkaYWBP+65Y/sMnQctuJyDhE0dsKCJNGLFXzwtbPU0U7R88/G8Q6cGdu6tTe4
pilIIWKlqPO48pTAXXcwc5E2nk0AedQqjQU2u3xY7Bv8La9Dj7I7u6khhYRBlQvjxxfA0EYvUJMx
2XX2SpX8z6UTIxGjJMeDxHDJZAOpqpmrkSFO771bSBgUXuv9ysJP1TAOLRcdcnANs6NEZ9kz2dic
KuAVw+4jHwaxGf5gQN7gEG186H9iLIlCVJpFa6KFlmqad8iek0OTeYSi2YJRf7vUOycYaD366Ivo
rmdU/5ai9kN0bV2/YLRptCedLT/HX2FHXAVrguaGS5j5n0ItzdfrugQY5382ml8c8JobWqwTD/EG
WHVfKZS94rNTmAhSo2AK2+gScRA02d2PyVeRJnKltZURvvd76IPzY1GQBUTW4QIXARSIhLlF6hAa
OLSiFFi4jk+d7yt3UFCIHsf9sPqUhl3kE5kY/K/vHInzb2IrwKDhK3iACSlMxbWISUD49LhXRiYM
EKqzJToVMvq8Z7iIQja41KFxK5iA74OLdja2uhwDUn89W0+7TKY8w9Xt9pm0OeBhFzxk4RQX/3+D
vmXg9KT/WyO5zzZs9bq2NSXGGWX8PFqNwtx4mvDZOso8eV7Vx+OW6aWXx88Bks4e0D8A6bjTepR3
Urm3qQ+tf4QwRtb98zeRQ39zcfG6SEIaPvGHi0cAOjfwTxRe5jIkKp+psQQzryxVg7+c7Aw5Bo61
5DiAeRjWr98QqfLxxy0zkYSGdKVEM/zpCrubh18rS6yIPtJvTDt2C4dTiWQIVFhkDqCdT4YXjEO1
BChEI/h9T+UoRnpXzvJUAgab2w9aRgeHO7wsb2cTlL2xgzrtKG937jSWf+2KlGmzX0nRdqN6PwRG
7p0UKHdwW+z8xolSZyWzdS1R/qq+qZ4B13HOFfWeZWAY3rU4EJc+6HuWAXUt1J0lZ4wg2ND7eHCH
j8OB7NfU52t08VYvUvP9NlUr6Od+jrm5aHoueiOqA0H/hqyxy4L4QiP0d6FxFVkdMlEV5BDdK+Z5
sVlAPZ5Tc+w7rXs1f6mcr4t/t0y1O4vOLaqI+mUmkrRUqBftWch2IU8dyYJcKunHT34ia7Oqwu/E
lDsoY9c773cGM8gNLajKEYVgJnAOHNO04OOhQocXy4evGjCflrAOfX7kNhRQHe4NyHByY60evb/7
aFazEY93UCpJ6ukFAGIXVSoEOWyW22cpPZ+ImJG7jyAckoX7EgKT6t9Lz3N0U1t4eopkJhnpPiUP
Eli7SEhjUugm4e4UPRKicE6IWoTzVZ8h1TpfbkorNt/no/Xqrh7JFd/zrH1TLEY4pprqhKX4ma1w
DFisKX5YuN/06/qDyqy1sS+uN1j+wy5V6nDDZuMbYQhml0/wh1IBkSbyrncWidHn+csolUOoklgf
IZCybGwLSYWDTWKXtar/CUcIV2UgfSBIbWLhbY2tuRpRQq/iJlJdNJim9Kqcd5aWteb/Lg+rQUuT
tV8eG60lBCOqInIcwg0z/qWr00XdwxQ5+OcevNkBD81xh87RBmgKjKRkCq9oNGlBHukq2o9+A0EL
UBC9vkegHqJTosFZx0M9RO1e6ftylRbfHSplSeSd2r3bPJotI0x556p4Q/QFZpfBte6pTwAYxIi6
LqUp0cmNwfmIOm5h3K7/SU1QK2HrqBguOGObWQyQmumJ2mqM+kTPvrfBOroEd2t8vuhMV9Ymc1Jf
wfckhcm9yuyt8Sc0tU/qtYlqiHE03oaB21mSIKNeJAtK0ZIZwjrYWlcCZQDuj3xGXCgWjwFRJegh
YvF12SF15lyE/sO1SwenrfZqfgSryxtWmv0xEoI4CzMzgU9dGgHSexWuyRMYrOAgFmC/sR8G8Qjs
/zDwckWAyANgAQL2/MqCrdpCuS6mZhPx6spyPIN/b+bH7FL1KeHc9umNV1Si+NW3/yL5Q8bVpX8Y
Xrkf3jAFiJwsEUBuq4Z5VGEG52WGo5i+DqbaiJv3PJtK1bTuHoMVH2PjEwkAEedmML7QdlVH0kb8
IAQczGvrJmWtlzxRqArA6MYnE87WVlenEBJrxt7+HcOT/mz0KQZFapfPwcwxMUd9WxtDdWVfFing
+jRA3tty6VQFmFvDMB323F4eB2AWOMaUCHVGQKx+qvfqIoKKiB5+0Zs2c/w3p5dAvM/H57cHtT2N
9CwE3EzF/vKxWEr/rB985CyJi9Mg1BbhYy//mg5q8TO5AfSpujpsqMUQZ8JL8bEEZp+oaRhI+wDK
chS177mK+ENWVjfu2H/4NZy2/+EpW6oXQJU+tSbPZJ0s5zP+3F863cPHSbaGZBxEiIr7M6d2TA4u
EuEVgTo/FdUOwYJpKJxjwb5dNWZWXvguRCYmmZBmQDMN7Md7tZttyPvYor/Ch7bCe025thOjF838
su6YaQ68JhMJm0d6SrTEyS/j5eW6BeoWcgy5xzU4xa/vKw7xNEiftrzwtvEpC/co4XiKwscjvSau
9/rzZrm+a0OeLQxXMhmlaN6IwMvPTUjQ63SIuGbZ3F9NVB1qFgZoly01Oja19w8JDieARzyIDpqI
8qyiO3w4e8PFWfdhGQ8uQgTNxuPwxiaAA4L0kpGbrnTd/oN6urtbPWyIh+G6Niq5A4t5T2Kf3Usy
bHsjmovFlJMhOFqMmyFKvTQSTsH6ZxsHSuasrsvT4ojxIWr4636UHcOFDM8L7UyTZPRULnMWljlD
xfJfjmtd16yAaAHHbC+PQb/U0uSD69bg1ImzqujZ1crghg2J3aGTIvRSOxQS/7YiIQ0JBdhIElBB
QfmyWbRBzhC2AkfSs87VIuqGu6cFh5tyn0nZW14f6eyXVEVxA9+LaljCPAGHW9o92KXQR9tlEUXd
83lrZCd/Qe+5TjgcIyxWLabYU9w+mfreeEB/2Iv7BQTFCe5dnRyp7oKLW6pcRhH39T/2qMGukCgz
KdZSKnNJM6CcN7921y5iSdoCCRP44tmhlXc1Z8+BaCdmOZOv64/bfKaySjvr/qTrD6w8dQrE3Xuj
dIr9eIItSCcRpZUhEzHlBLdYzh/kyx/2CwFT1bQ/MmjfjiO0d1FQj2YbQlVTLWKGhh2mqesqQ1na
luAOEjVlGzP88o/vDNJ52iTMpADmaXWyuxc0SLMtqGYXpALQUTbe8t5xHuVXRnYFmQNEF2MhRtus
S8aCe4jiaIU84QVbVwDVYN/H7WSZYZfLx4dmsXH+tQOMmXwnv3xezVAhUNTG5uuMStrppXQmonH0
0bFWB83ur6NWDEDjeXRrBiV5tDS7TUw+fO5J6QHSAVDHcGKvofrSfQ8L8Unybvcx3EUGYbTrrWwy
iw/cBs78csnsN/ly/C5B6XWw3D4ORX4W8c3AhceNdA8XuHsaI7qcyvPRSlt+L8YI5V9o6u7DcjuP
ozoauY4DqjVWmPPe/029zoBjud+pa9aKSOEvZ1I2gcYRA2SLFGwl3085cfS6T+nrWFx4KEVuc7zf
ig8Wj/usbqsWGPywNNtFfmeUzX104i3b27mCcx9GRaiMI5ngybwymFC61/rX0LuxBgrvPg4yzOPI
TJZaADh3YPaBTP0/M6hSIhAJiMoMgXykW9QpVzyOwuT7I0sYO6hseqp1hLNVHvx1QuOf55oazr59
lWtYzueOgFryCkLNM6FVG19v5n86H1mmmVu7Az4i+2pPlQOcj6ghMw6pUirYGTM7e6L8pFxtJhaD
6CHcptNBdd4ONJxG15QFqGTKZVkSwuEIMvk4tQ8NZpSjA+BzahVaU9KxgxcMATQjsNwqONGbuUNV
QfXA/8s1GzKeSbhqU56LGF9JASLykxl+uLC1OVZm1INfqiz65DU+DJOdREsjfOQHd7OiwNXb3neh
P3UrHoWfkzwUWGIWJsRYAm6K4wd3Hd0/Fhkj3jq8z1Dx0RnYvDtsTCYUkTKUV2L1fv6zm0h2xYlm
CWfUNnR0wSJUBX9uzpmMqwIr+PogBjH3Jn9dGJGK7ASTzE0ZCLwLfUlte2UUO0HgM/vkEoued87K
xVpTgcjvd/e1NMPnDuZaCDeyN1M/iLl6iwdb+FFLLgfoUIO7OzTGkTHnubXj9uXeQorBB2xoWsIt
9wlpiHV3baJQdGUn3WIEUJuEP/qB1DO3dniruNIKcypVQ8TQNeQ3JIb8zQOYPyBdUA+LDXXTVPu9
musawxQGSGioJNbGP98IIcuznxRrMVfPU77pL24+CLSzxDobQVlBIxLJiH5qkyn3HsnHPTcfpfzC
QLp/pA6ouj6RbJ5qpp2KrhBpRziUqn+WkEyIZTdRA2Y9KjNHC+sCs3FHPZ9+e6Dki4FUNGxhdciY
9LDzX0rTbtoJLLRTX53+nc8O/9lylISbbnmqs4aPBe7Gx8yBVdswQNQe+XsO+8XAZXm0es4DAGvC
QWnRs9S/6uCe+YYlY+MY0I9K2tu1ahz0m6MUcEdDhxyeVe4Rc76oRY83EXB6HQTtPxPuaIeRQGBJ
hQB5NfEGw+/sg6hjK4mMen2irbFZfm++SqL8fJu01THonA5wcqdRlDgKPRF2WWReVr+FQQhFk4C7
m18dy25bAGx2Y8+yt6g6g0BbW1cgI9jg/+z8iWF+sq47n9l2K7gtNldF3V5ydr0w+4ZJYp4CqFKy
AgvMJNdcNbF1aE72KcoW6J2e8JRik1eKP5IaT4uxuqabi5VxAYRVMu4U+vamHJAL5myzgU6dJO9X
KEr+c9h0Toxc9P88/WZ8E6lA+a6f/Kic+3UTZEOVH9M9tDt76VVOkzgGyou1vimlW5SrSnf6ZM44
JvUhKS9oeGppGPVccGjLOZE6g7ate3rYQjAx4vBn+EL2qM1XplVI6Hl8kKIFv5K8jsL6IVQUfQLn
RMvnhPSfJao+1j9WnKtbB+4AhrbxkNeVticVtS13e5EkN3fwEQKXXcCYDR1b5tFmDXmBRf4RSBWV
E8B734zhz9OUP8/eoBC66ukB/qgxFmbmck/o0svQ3k6hAy29JHcEi2AUsFETBAQBN7aKMnaZS+VZ
nKdV+brx477POVMav8XqZyN4v52xeWTdAK8f+FtZx8GvOQXy855D4rrb44nePZo/G/OYRzLxGJcj
TvCxZmqmjgKdEyZ5SaJblTQ98shzVpwydHg0zmjr1thhDD90XlupcbWSG6ZbzQMxajOL5cwDBi95
/M5Gh7R9wxaFg3k9fQ/AGOgoxVI4Asc7kqe8lEy31EqzppLRisuwxkVP078YsfCmCmPeY4Eelyeq
vT2u71SxGFEZ9E9OpuxOoIucu7LAJa10NWEB9n3dp/MKyNHxypvR8BEfrjCIT0Dj8VerTxrbfjzy
Lgy4laj3FeoUmZjOtUFZ0GjLSUaQaDYmSKxHRj/Jx2HCIYrT5FTJscrNeWUKDf3Yoq3qhe9Km/Ro
EPN97f3o8jSY0gTcCQq6MZ4YVZySB34eEm7ptneR0/Oi86QE47QeqZMFG7bQ7lDlJYOJl2YzAKAh
+V9/RN2un+26etDX+Pza9oz8Bsr06Ab+ippv9PGW9AQ7gPwgqitjubcUSCOeA0ghJpqf9DO6BeS1
o2lnhfUmgzXQ5U4S2Bcsv72CWFKZSy9qN8J6YhzCWWQ5UR/We1EVwnQcP1WdMfJPjC5ONazshWsW
uAvMuNUFHYRNXLdU1YMC0vnJsGoNyVrb2ARK3CQYRbpN/FS+LIMr8fNbQvGfIeQrO0eLeEIhvSBU
nPpxCtSbXx2GMm6wBWCPn2v+j6+2Mrew/hlZTYC5OswFSdOyebgx314GAkGJJ1F5TABHCpzro8Tt
yPjTsQUxGydJaAbm0J7R4Gt0SxpUV9V6LVIq/uZzGSglgtn8tLlxluwtPcsHGPiAVgj2NJRcDgEV
ZqfHV9oacQ7tSj1tJjJWegvGUSpYPQoopUy9cSLBZIzVTlke+5jJrqyG42Nn6831N72O9QZLeIn7
YVtRvZ0Yel7lW5X2g/5TKKQSmEppbFsukmhwJSnZBNikbbZ8EFlSrtGXxuTn0kUVNa03GHHjMJ1H
D1OgIg0lu7DeKckSxKnUpdQ/cFid25t+wmamP9w5+yiUk56PB7kCi/cQOV5B2okWeGm0mc0f/0dN
VWsACj0vQgysFBjnxm6q5yocomuPK6WOSQhvIO8ylaoQvqj4aQJi+pLEx/0YSeXFaW/WcD7oYuGH
gTOBbStv1XF1VRnX+rkNwep2XLG2FwYa3AdlECwlYiYciPs8PtyTCm1UbrILHLkZIaaPui6me/Yr
xlSBl0kmAxWkbx+0HFUDp/CQ4Jtkd+8lFrZ+lTopQPCjeyohsvyPLTbpgTweSDzaeEoIrW7CqsGo
zSurrwhnMaigufgKhgu/jzeGxGV61WMbKU8voXACrBGV+g/vJzc8QkOpBjd0rw0mGrViD15Ik5ta
7RCHkB5OPNSGslhMwmyhlzSbcuHTarhvF7dM28383m1Ilcgy3S0+R1IOkulS+hsg2WJenz9IuXno
ZUUm/Yc89PNcBDafDSGWAc8Oe0D+tfS4Z5Matg6nBU2BmgWT4ZGgYlB1mNBusuo2r7+QNOnZVxux
UODwpfu9ThxmS9bLSrIe8RJIkIsmIUAcWQqX4qsGneXUDi1kQ64/p/Wy+vyp4GbW1LKEV7oPSljx
oK+sorIoaMYyXQrXNARPLqBiYeXwKbIbpnEOLrtsXNbIphltZOUWqmLJKbSb8n6fwrigF+lJ7xDj
FnAYDh6v+vJe0gbAIV00rgDL84noIVlcioki1isvNnqkgfPYSxNE3YNENKarUSV5UgeGePjoqpJT
z+Styu1cvtEYGh5Slp+dEBn8QP/Ey8d+don4EoQEJWt7EcYv/pM1/hsRyvQ+98EAPUcasSAlmPGj
T39mJK9lA52zSsTSvRpGthoSfCSYaXrUhyucZnQfuP//nUb/21oVxvvg+IJky1pgMllYBxbUKKIP
oXvewF+i2Hf5X6Saolr4XrjIwwaTOyKAl31/t/IrQ4Yq2i+TnD2Ho1d1EuMo1qhWvjsWp8bPiXCW
VQsmlAH/1aMz2q/BgXrlKf1d5Cr015FF4kl6SHDX7QQVqFOB4C3hNUIUmIqhx/LR+A3qYe4RoyBz
Zk+W72FelhVQn+I4q6qCsv4aP5V7B0866X2U/USdVl6Q4SBg6AnM3NFmkR3WkPF4DnReL8cd62oi
EOx358BLActtLVp7AlWAP8ZTfB9F0Fo9JWetknncZcqSsxT+6cJNCGG3+BU3zcYyd/Q14PvDf6yM
oIlsf1LhYXvhrWgMf3Zy9wlhT+Wa7pr1TrH7z3Te3Ha6I6nbkJ8rIE0UD19qfXwtu93fEsZQursS
9Lw9Sqyk9MefnXohLGlDiDz13mB46yZVq6PSInz8hbY3pdxOfJY9K7nz7VAupaoufnbKFI2GmHOP
aqfrltdhkG80jmxLb4qUz+v78YAQJ5ylyPAVRENnmP9QO9LyIld6d98KsPotM/SDh+ZYsQh62SCc
rRFKD+bxKkUC2tmA6xbARsy5n6KqmfihPYH3C77euTcBTctCVI9I5A/LkJ1TSHZ5bsA3KutqFVk6
W6F6zDkTYvn7cksQ3zjaSRk/R06SkRCjAcwTq5dk5moNHEOEXin3XVNuUTCNvrdwKjByljS+qXPo
gavQmPBiXcKTh/hQYaXzGxLL4UtrWKN+bDTebc1xTn/iMz14Ddx+7xP7zTcErI6SJd6sEq/qd88N
gtXdLVyqSpnsp5LsCkAKtVvvJTd4Ar2OuD0tsCVT8zdQV3MQOBMdMOyEWEy0+w/CvCgLGoZ41rwQ
Ch8UPpTMbjACSig2icfbdsXFGrtp3SvRf69xamyXHUn6k+65JbEkvjwtbuqeFmfO71/xZ4LpyW8J
gMj7O5BKlpY/59WWZgPgbgMnoHjukitLqvk5ic4McqnETb3634aoXT8Jl9E5CTAJckM7OOC9ERbs
xicH7HLpGGeHzp+btzD8mZpQk/ZU/Y6TabluqNHq9X/BuXCd/sDwX9ApsuV8DatcB0AjFqN7ko60
S5zLqVHORvhUgsXmm6VTQZCSy3ukWDuY4LMOsleeDMKdxWvcvAnEKt9wrA5Z0f0MIBytLN5pPl1g
r4zDdZp6j4nZhvfB4X+0UWJjM2l8lR1oBDKu0U8vtAGHlKoiTyTHIGVmEMCNgvbpfd7hi2GQl3Oy
OWa0Fv/VWamyvfI0QhF9eCJYeCZmQETOoIJl8WrOm57cU7vCHfKCRiozd87GiLg1uPAcCDZ2CB6m
zJr5MLOFOB994YG4zFE+j9PwxDUUKLwGqEkqXITwahZPfqS8Ni1UywXpPPNKI9LUN6gcSdroRKWz
YTtdjB/LebPC0ATkeiKKdzWgxoWjd4OH9Ccv8i3ispGPZ22CyGbCcDQhSmFNqugi7vmDUfxq5b6u
BW4V3MCcbaqLSOXH5WE4/liimehzy3MochKB5PMdJS9/noLCvoPP9Voa8iV0/WbT760kI0ujmhLk
GN7XRptpOZePMCCwfDEkCEHVgo12rKfC0BUHIk3OWXb2JHBy+ly9KB8c9ITLNtDgsnhgReIAtom+
JIKG9SrQhYQnHRZULnE1oCUViP0CDAMgExJDI90KhUmkKsyKTHcfdTWrNRokCpROW3YDVQSLPvAl
4wyLYY5FdGu7WHwZMbxfbwXoe5+orjJrRCMZkpJG51ln0OucCGsq7AuV+YbXYHAq/jWClkQajK5L
2Z+Hp1hQUKPZYKYO1XHeVe/FmQ8oBthK/YTX6vo0JfkmrU54oawBZFRX/7L0rcJ2b6btXJLAv+D8
fbkdsANPVXQgFOOhTMeTiPsCwiHmCWdURof/BS9SFBYNPgE22KfD46irFfhR/ambgaUo4h+5moZD
hBwcrkP5Ou78V4CGgVx7N7IZIrS8OxUXdo4kumzJBrDtEdQc3rvJ7g1wNgKnXemRx2iiegNFH2/S
isuK1FpBaKLx1LCcmBG23wFHDlqAIpo1AboUxnESgIAQhG7hjOZuSUocOmwVP7M0kvZMOgw7//4I
alh/t8ivzLHsIvJoWBqAUMGPe+4sQezJJXcAraHVmO4Dgwpd6/PSZ5TPNkTEFz7BROrVZj2GAeUx
X+dBwiVjwXsgIcgAfq+13x9LOWuJ4ZYGmGdsIO1+Jnzro+Rs4AFPPZVqVE8PAF+4yMcHSFIinPr8
kqh43OigGMHNKnCvvrTDU1YQUlu5t5hCd0clr7ZJVh5c6cPtnGhxAvtkUvVN2vWaKyC3DwfGcLTd
0jeFCGHuNOdHDERjgbslJ8auQxU4uMwU1V8oX42/tA6XNZN+v44fJ6sBsI4tTlfMKWzwhqA3+/S7
o5RpwDMhYT15oYnvYxf6jI+4AowS/BnIZ36CZc6+H30xhljG6huO/4rh7EAc+dMOYWKncn3Mn/JW
QwC8HjdKvInMaR2m+06NFOC8V8Ie/6CdMoAemDzFGArYbrkfWSokvQr84N+6ioqtfIhJQ0Ha4qul
WqxGCaFXeZaGEnTHkUxn8kgq3ijxl29oQtjKZLwmPL4BjJ/Hafbe4waY/03XV5sxiO9VFkTzF8wt
OhMmOYYKYzFkbRDyMQU/2nBF0JH8w8TWvmYPQpEmrt+wFd8gtmXAGfl1I3GHP/KNYv6Z7oFC1xRF
/cDHBxzg6OEIVFz395fqvs16zl5eGa3DBu0rFGQDRK9GLgGsPgS6AtykTprDJ81h6QhbB11GaZNH
6/38wmZlCAsJlqjMQuXJY1TbV/wgdN35tthzI0rXz2hvOSCwMV4OjaC5cqLRCOrxViZbBCQBoFcS
lIbB3rkhmAcUNwxBoGbdvAHFOuRcA3ZeJVM5fYV2cKAGwqJCjUK/6PkhJiReXfaJF0kK/0y+RRDW
POODT5N1CswVKsnr4CELdMWuiYq3pltsEi3SkGnhthBRxmpTB/oCoqOBLxw7cMO/Fn+jpOyDjFYe
sowvAxlpw5xZpo4D9572yWPlHqduE2OJ5wUDPbZacKOk0oC4JAdLJlFpzfT4oZ3XNFaDUvWUmq45
jXz/Hm9r+NpLav1crUL1oUX2/LDnWxsT6OVKNHusvuwvW9ObRqBM3Q+5l3J+iH+YaNBNprxIGwYe
v2p2etv7jZ2YlFbsM04u1m2Zlidz8e8hOrK0FRRzItNhjKoCJPPyPny3YyVqx0irvgr+12Kpoori
uM5Idm9VfiM4cjWr4GHOCdjAklaUmSCjMlYwaJkwkzzfmKTqTR2HYY/gYNjqYxH5I2qYhdtChHmf
ka66P+md9hKrFI3cj55lb8WYIXO7/lCyT9CdQlU7ZuugD44TA1aqjut0JcuCZUWLYFUKyZb7SpiU
UH+uukmlYnh+DGCBSrYv0SBrOdpmNmobOXgT1vZ/C6DsrhnieHcGrnOCGLEs1vsdTa7i+LPgs9PO
OSH1RVJHohS3Tl47JcFAvwhx1HqVVrLH/SZ4Cywq8N2eiCbGp2oyTBqnrjqxJGca8YD7xKtgutv2
oq8AfwoxymaUa/33qhFX6pOIM5HtRu0W4iO7nI7KHHWGej523zSR0Rl5Y3NqpMizd5Fnv1baM9KD
aLSATNB84fgWsAuZphYtsvuFIlESWqypK80CjrrKXem7dBd0fIgl7x7fYowHY/rI7s1p/UEpt3O2
RrAo2Sa/HxSB4qb1xxP/idRknftV19B1VZd5lgdLOQSpk4DoWu6Fsjd5S3iEw/MFHDBmxfv2qDDK
PwUiLsEikvVCYuVn8RHQvG5OSFz3rGNcXF9r/m7d0dS5mUVUzR+TL2H1UIjSnx+WMOFjc0XR7N6e
26hGyVmsfN7g8tnfln7eSgMvt0QFPKFBOd3XL8sNnJgnAgpWwGkhqvrDimbp95c/WcRCTv2g8Cp/
AKu8snIGLfNL0kT5Q7WiRvzr2ueB1sO3g2tUaCjbuTCqN207i+dNpK3TUmAcpMHeDDZXZTxukvrR
XYZ1GpLyA0TRfx6FWcHkrjh7LPCH8pihRkJKwVDyrh2Zh6uzYW9WCfL6ll5InTzQnIJp1UrEOalF
NgciW1+lx7q8mDZXgdpR8Pk/evfTg5G8vQJ/hi+w13mLhRBThcEdP7oC6KrX5b3ZybNEMPNIYUw5
v3KqLLZYc6miSatV/O4b8pAt2w2HAAd5HFq+uWQ03mKyjwEtCPgh2D49xPvk1kVHVyW4xdNx5E0o
aRLhCZsY8JXxVCM8ESMxm226tj+FHOVW85L62cu7GG2wox4ov3YjRrORB79vkvozXDqFIK/0CVoe
2C4iY8GU37yVmPkR6MuhGKmU8KIm5tRHob1EDELlfDSbNUev6mnctnjw8NTVcwIIKtQat/4rkfo6
JtFXjmihEpGvmA2qjrhNoLw1a2Af7QQIv68vlZuQkPHDwT1X5A/Y6gw1EaFcVm67BLDplvEeU0VS
jv3OT/dh0Tn6X2PcZgj2TfbvvGl0cFseyiwW7I7aAGKmo5hXnLtU2xTw1enPX+4LgbDxDz2kK/+1
gs8eOlk7emzaeFnT1HVja44Pd3ucaPItX6Dsa5caLuJ/NLr8kJLRpf+Wkdq+lU22P7ZhlUYup3Iu
UsInY+FnKYIj5Ju3quuBh0IxvzyOwi3octd2oSZesNE0Z68YjjNF6/UNYYlvgLsg/gG+RHaI4hh+
bsPuHH7bRBlpu1y7P4VJta+OIuY2LIbHuQAInrmDJzwG6q4avmCNyLYNUaJ9RD+v821Ta/N3+83J
AkWB45YPJmqFI7ZYcYGsIRPAvD9ajEB9aLUrM6Tcl0np/Aef2EpgnPlPZZKl1SQHLWUHOnqtjgJs
fF/veBHMK86N650paxg+/vDUuDy8mh35BQ9hbIdRwn8xlZniMMHy5bKanyxfialDFdNOViQvdleJ
1YXiX73XjR2YSpM0MJ4gp7lq05jA7/hPS0W0iH5/n7XfOoS1IKv3y8U1hPDxZTTMbLSnGB4VvHnM
z8tI/HsglPI0uyC4P1BEHsWQdTgTjkqhCZiiUayC5JQAWJksTS3eXV1mexFnc4vp9ZbY4wkD+eIO
6uQW78gnR2K+hFLbgx1eplSMl0y+UIi77C8H5jfrxg17xqIP0N/ZxQJCHG4m3AvBDqwIwkotaq1k
jP56ETG81Fmx6FsPhEgPNFvxnYnKAvkBvpljOlJwTwxyyijV9wtiUspQsdiOEFz1Jq3rOe9RHyqj
H11T/cdsb1fmMrtPEJTtmXYD5sYoc5uQiF+gHxIDVnWxqOu99Ft2T1NEhLO1xPa6jBpyHK1Wjp72
waD0iajIrpnqyRx0aZe/1GdbkclkepPWTRwXcU+zRmti4csLh+ZbvO+2/cR3qu5d5m3cT1dD0LGT
LlRO7QeO+BD17566K9hTH+RIUuioLFLIlv/KEKzjENSopLwOBke8KgdY0057ZdygY2Cx+vjiYP4f
1eU2Zw7KOUrIfuXkeYHGU4j9/rV3XnFOFOykfL8iXdP3H5vemw31DykwqyT+xlx8rBn1AViBNMzX
fyM7CoLSbAFw9mZp2/qSjv48tDZ0EuQKwPxuCletTfzbRDSvKQFcHStpKwQ+IQadEKIVoZl0hY5G
VdmmCYM28nVnR4w/FqnG8wXz3zlfRlgS9fW18S9SZJFlrqBb/yv7fKTcVduaOK9koPvsbYj+vPyG
G69N5oCjotQc5cJUXULdSyWbPW5FnficnwTWIMuQsxytcwot3YIbw9d2y8IQf/QKPp2ytUHly8fX
GiS7UoctyNooKqqRhXwvQPTy0pDp+AlHYJg4o/ucNHrUeR/z8flBM218G5hbQWh1iP/w6fpKY5ay
dAA2L5XyHgP4xUraYQAXJms5vSW1MwFgBa/43yIcdUuuqOhE3WnLNj+gC8F5vO8cz6mPIp2u08n7
X7PrdhnS5a/dyQoliz0vGi36+nv4XGMe6J2jRJSxsSMxmDRBUstcN6juuDw47hBs1C9kQt9FwVNd
ivj51ZQFwG9P6j+zlW4prZ/jgv7koFzztqez/s6BhntrAwTxfIXqD97rCW+6FQvw6l6mxNzTTZIN
OITWoAt8beKtAHLMe2u0XMOmZD9iKFgPP9vnt7MQ0duAEH/9PnjKP+ZYpDRsd5q8Jnti6j7T2qJ8
tl+4yE7p/CeaxBGaDa8NvjORraNgtNQWjuM4hDlAiGMsH7Aw96QYk6NjacrOUvQS20g51P2wNAAv
3ImI3NVv2Q3wb83oKFtL+k7r3S2TQZRL+0AZUqYZaPZOyby0mJtU8a1am+H1eBS+seoXO3Vz1vr0
35nfeNlwUuQYOtOAaC11kGr2B3Zqh2kT5Q6UiG6+cnvfGMaTKSRxDkXnvW9W9Bbcza5gymwoPeD7
zR0/f4oIKl0vy9L7QA1PS/woi+mwTWdVR1w2cifwsIgVbHhvbQiF7HpNkMKSxXAEMs+lrEVfhcu6
VaHo3Og7bDbJj9hJCpiF18dt04qRP2JOcKfKhawWGQy8sUW8Gyfn9/04FQ0GS85LBIxqZyQxIfWQ
z7bA4CiV7f44zHYbU8EbPa2CDbBcdyOcuUM/1a7jbhWleDSISpOXkBQvOkjPnX+R84UHMRAw2CPi
VMs98hPy6anunFXykeEQlGphjXg1VDyp8vUrFh/jfkeF75PsyrYUtklqDeSMRsdA+49cXFaBqxbM
CVT5u8+hl8sFmyIMkhtvU0F8h/sH6I4+GCwYQYiRtKDtYj4xYCFspBH1wofycOR+oXJXHhkMdc3I
li5PSy7Ds5No1WKM+De/0HAT4neFe35LxcEPFnqz3JcvkoPV/Z8EBvoU/JuCxwWk8S0xRsZyCQFk
7vH8a7fjpUuatDmwyZ374wczkOpCFlFmK6SYaRumjsmwWjcEyY7ZRhMSOiO2j2ReZCaASGWjeZKn
DSnA0Cd1Z9AlaUXvJFxSpO/MBUXC1hmHFozX/OEHmyXfSsdCAbk3Y5udbnhJo90Ul89VLC4YkMIp
sOI1nGI85g5uV/At9ma9ROs8JOAdUzNwIscDcc+DUhxuJYEbWXB0oQxu/GEDspB5wJTIgY1f4uOO
YD25LCnHGOi1BT98xEHCAcHXGvP7NqQtyCtc4U/on21/0d/7b9FwgTAD2HrVKfu9YJ04beyQshat
NNVMFRh3yvcAAnGsoY5RRkMwO4AJpyy5RxLoivPI6A3ZhnqrO9PCF5mTioc57VEOlUY2obpgFbFt
AykYcjz2MPrIaZkOSuZVwN73hLEiSpfRXx2i1zR/QV5QJHajdiECi4vfqRTSoX7GiLL2zVnwHjxl
uaKeD1SZOW5Kk74Ei8zmd24yz0Nld4wl5zubfsUsvQOkRK7MBq5o8QezuAfWriVQV3bbDhJHh8Yd
XsOu9PPWV3uJAVb4yeSO/jDvJTh8INE7dKm3EGMDW5b47xGPbZbOXo0XaTes4nbo7bSKCi/63OWT
b86aWRdy620BvaKSbhMChWYmtrjk65EEAdMZMtH9opmGI/1T+bKpIND/bhtY3bhBfrol6mkY6pei
V/6iotjQf6cg0XbaT4AfO0ezkysNnJOI1xYB4w5Lxw+tnrawSTAzxX5/o9SYdcU6FM+2NDnbESMp
fIeFEWkM13/ylAOm+AWNlKC4Zl5/R2Q3VauZQL2TK9T9KRLQDIK+Yziu8R1m/1eqgxf7Z5mF6S26
Cn6ZGJOyHFIgL8aRx+YYgXMjBEW63pd5r7rOjX5q1Uh+Cv+qmna0F4eo8kcBGsM92RZlowuK9ewI
4XHedu2xeWOrzPsOMcW2FjC1TVIsAsGuBXr/f/ZCGiH9R0n2uKD0ZMviMooV3mJav8ZLD+dcoJ/v
pVsz8HyBEcPaGRPdkxb6Dj9vgrtR5134tt9H1vJHudBtABUZ1vs7kFBSd86H7Bp3dWcvQie3fYkN
4nYoXT5QhU2PQzgyReGw122H+aTlzj0MhVnBynk+S3aiT4HeZD6oQT5JOM6VoTtFMO5lC+PFm8D1
hDfpxORSEFGqJ89G3ct+n5Cqn5LAU6x8ckaOe7ggmPRj3Wv4iKB6Tp2FS7HL7RcXAQJLI4dE37jS
2QNA43IAKsd7I2LDrHwPGubfpTG7SEx8PDrbvyvZRA5hpyi/p67L9lrd8y4qjOmFUBhpOs8MXwzw
ls21IpKQeEarhoOY78YuYIOiMPMlEjhnYXfrCFIa01dvdeXkxrVtoBBpWcHfrUbjaLVznTmyftxP
lY4V8Ud9P52zMt0Ys0Jre0Upg1g0EjxlSCq3RUgBpcVNsxuNyX0wSu+sPUhniyh7BixPEnNoh9YT
y6ac1llckd8ajyMdPhZ0k2pUMfYltK4+7LlAsTeSQ74XiitQX1xnzsQGviMGNef9t8C62jucYNSq
fBPA59rW1wz1gVdTQF63XF+ao4buuYgpvG6fvuQq58aIUvy1y1P5wVlLIp4/OQQ+yfuE3cMcoYPt
OD021tmMmOLl/tr/0Qd668tFLC1V+8TgcR8oK65mBbmfVZVVZ5jJDCv8rD1UJZ0Eey1MKMMixHPA
yinLkMBO5DlcfHgI3CCSHsyE38bKj5KyDknETidlkYvOcbe4p3bHj0qdfDDXqa3b6M5IQ+7YZpDX
lVNU2p1R5w/DJCHpxASEzA0WC+Biy7KahzbwYtIdIAXKyCsJq5N9MRcxPCn/96lavA38XeiCPcFj
R4DOyPbHk0hwKiw1M695QMFqVVjLDsmQ6Qo+KYEd1wOtl7i2HpQrrvc1Jq1WrZnp+uIUwWVBPrH1
+Al9m4F3TuKgfgJF1MAFrG5ifUbKor/+HikZMa51F2YV/Uv+yzhbDNFskfslw5qyx2GqoT2vEvCS
vquk3Nw2mejA73IdQuna73GS8J3JlzcCTSWvygpPufypZFnfGTPQ8s05QliwdJ+fAwpVLMZcqcl/
nXo22vcQGTlqiW7M90abG+Kt+6OkraIvT1GT/po5D47JzjupuBIqPqTn0aUpBmrXJ7kC2/LkBK17
pskIMFIPly9YLNoKlLbp/E7euemVMDEBG5QdXpfcUc7VuyTVGWHtCgnbzJYbGZZ0uYflc6YvmZFg
WaHMSw79wqOUkw9NnIRtKE5reSYUitB0S3Bqj6PJwrltSJaKMJiJXhwn+SO9YBsohKZf5fofwolH
FBnyzpeQQ8ix6IODZhmoiIOdxSuheTHivu21UbPFtUMHOyRxXmparC3GMvjCUq0yz8jECQFyqN4q
84g1urWunSpTVSOnyBmNUugZHMeQlDovoIfkxtUBwWskyAz7JVYi0PL7y3eusG4UaDRwFv8L0xWr
FfxcrOAJyvIYGl3K1zyv8fzi9QYypPqTF9AosC7iC97HnywRjO4UU77nHlCEJ4GowwsAQfsyzCEB
KqNStuFLKhzBACmZ4HtHZHOf1Nn9TL3Gq7IgG9S/ol8UoZ25mOcxLISB1oLgMgMOrgYxMRg7h6Hc
gxSGK43PXznaoZJe1M8VytitXWvq9AxQuaU+eWuQlrJOsKedXq13KuHEmjsOsBzmiMxvAZ20OwbK
67OYht+SMLvUboikrnnqReJhSqSkLyhhUWWOG4CuT0/+IXvEjeMqQSam1YTEhLMiK559ZClgoByX
eiENMv9Mqd0cDp6gbxp5/AAIf7otijMsV+lK4li7RFy5rKhNu0JeKoX3YibHDBNFYNO9aUD/XovD
HooHSI816VUs7YwQaBBpS3YCNTO4XHMR9HPGS12xqlT+iq/ymIt0gmbxsreiiphovfq8kjaxRnN6
XG/TKgXKxCUfp6gkobwUVFo6gHfnNSCzRGK19FCqnf9jB39sOrVLxP1l/jJHTc6yKXAtJCi6+neS
MmzopnSyH3hrpL+vqYy1bFYCW9CMfzexPB+XaqQmaXJrsmUA15v0Qs+ezxZqGN2bveJAnZU9zfHd
bBC0HUQR8b18kO41tXbo0GR9lc+JqREiefLFJ6U5Iqy5FllmGqLZSdsZyrPayPl05l9QYku4Ika6
wfAIW7zbkneI4fcI50M9UQYLF9YhtW1KT3l3c1+j8cT/6nJcpLPoZJFUZTw8NMpLOI8vIPk5Nvnq
BwDEDzEJA5/TddqLv1BGJ1glv0p8wWj6qIsccuk0j3GueRL1GzlRXevTOViY7qylCtR8BRPGdaz0
zkNJK1sdHXGJ/um8u6puZCv3r1XADsd7wn5SYkmIDzaDi3woansDnkl7ffVAKOptu4p0UOvtrScH
lgVYY5kwxHZyAlVIW4eXf3bJ5WNuiSJvmhDUQ53+SaXQILeI6pMPVAEQ64icoMZB1k3ewiKMVEqR
cNGZjWAbjU7mR0odbp4Qz4uiyL+HkgHoZdXx8J6ALRKgtzhOdrtRMcrthtQqNoKqs4ee+oiyRMZL
YBBVrHCiV2l/S/E1EQzQdlGGSLcdZs1p8A0jVpRevw1ZhC9t6fLUS1kPz307VtHA31x9gXp52Gri
A6uj4VrqULihqPl1nUfQHqQyTUhQwiCAoK7d7aVOZEYQdNvPGonry7+0c5UYOwWJXFv6M4eTiZwx
JNG6721rt/Rrn9grTOV+6MZNStBxCay0+nr4WIBtqn9UhCYXDBHOWuffuQrlrzl00bsELZ6Ys0GU
Y6DCkOAL0DzLV7jU26tgzAUHooTw1XlmxKaqOefTCrDvpI4Jj/+qLHxZT4dhuxrQFoiAJFG9M2Vs
fsnIZVaU7XxBhmAZ0P/q5pe7yT1eXwgdB6YlelPp5Inxj3i0M+iDHxfpBrCR6uB7iRmRoyyHz8US
ixDGdyeMaf5GEXVkNGJEmi1nAsOYM2M3uCdaBYUYFkce0bWpr+ubmeqF6pKxLKNkCDNtIY5GPrkV
agibZ8NXKJRwOobo6t92d9Nzptdz/nsi49qmscXc+6S9DLT0Bxqk4IaZ2VZ3TLAr5dnAj//5LDug
kF7zMDWgSgcMlStlGL5lZFbU1dUuBD+LvUHQjqKTlUYFRYV7L93QMSTda7J9AlsrGxK+Kro/+XZr
mA/XfBb5K4MLMMYrsihjJi+F9WZIHNHSE4JjTLWhaY9wFm8S878vkTtFRTWRfmV7dl332jp1WYQJ
674ExrkctWNJ+kROTKIfOTb0/4wZl2oj8uAWlErqmhi1xzqY0cp5gF1b7SBS/X9HMA9VewwCr7+S
sPHORP5Sb1oShxjl0+kuFhL1ROHy7cSfBFLGIp0e6J4LPhOFVX+VU63oEQBlku4+PMu3GOs11V0g
/gwqCJ++Yov4jvZB0Yj7I745nGLKvPn/xHkaJ2jxtE/pAw6WIZ1o2XgdVnPa3kYOT5Hd/7F5XnRl
IMTQ7ApVG1Th22q7wWtncj84cvLyPqXNXIJuysmJytD+cIUSCx7wN49FfWryGJvHmDBJt83KdXrh
TJX862SNNlmiOr8/c0kyBNF4yBeTj6Rl1AuDWdpJYtxUrTrUjFoKncRAFA8EWD26kJ6hq3BvK+Vj
jTjQIYKTpcT7PvHM3AFMT6enKPjEBNSsPDX8PcYSZbByb91IpjtTShll+5WMNHH2Q0cgLL8BQ8cU
4QaxPjwqQOb6y3Qd6HJewJo3cVy1lja6RsuDiad9cRYjobkDyOmvwhXGUgosPj98nFFoknefgicJ
2UQsq5rtJInN0YfHlyXW4YRn5VLZ8ChhKXpMITRpMdMpFQmkrou8tu4fQ9plgn2q4Yp92I0V0yQs
MlgVKL8Tf2kZkaX8NV5a2upTJZcGPeW8BYAJE0q7TlZ1VjCjwthGxmEONVVIrIPWTnbzRI7hIzVh
1Z9vbQEvMiRUYzKY67cIFuRXwNTv+J4xZpZmPbjfQ03VivRhoaI/FmzK7Fe1cpdWZQlgXVEjuFl+
cPN5O2KfkIrpoBMYDw7OOUUyDw/uIOIJgC16UhSWEl5lsrmgs/UV1tcJ9CWkkEAAqCkqGqatVUMB
Ma5+ml7UgGWo9w8BvyFq2UiyusQahpfr5XxVhK/RtvZG9M9IGQkEDxiIJahWsyhvZpZbL6gjrRty
6f74eB+aBbDyaj/IM73FYQ7WqtmQsz9/ki6GxOUspiuB4E6w/TN4SsfXnJSP4aJSgQubodr4jMnb
hu8NnpWSRViTLGsrggjACrbBrxdN59VwEjdgkqB8G5sxXSmACdgLXH2TTr+5MRwMbYR3u5wKm49E
M6lengRcLjKiuWJ1D6/ud0TuC9K3psHmzdnSxFwfRsGb04fwb0UtDrjVpg275TLZTUEKJY4c4Nqk
5zm59Ust00OhXiSaBNP2CdsQsVqgSsDmW7k0LWLF/EGncb+uhrvp2ipqjtoSu1BiZ9GeMokK5GBY
LqxeY/ljYjRWQf9QgbhbfNFkpPkFuGlyNzk5BnUpOLSXHPRgFdh68MR6HdnBxH203QYiQ0M9BHcA
yV9WkhtJRU6kawiZA5AdCAiIVyV/GIUAPQz31OIoE04W1U5S8AKH11P9nVAHiyfhp4I0J+cz0vvz
sChWREESdZIWqWmht47o2gvJUXSAsCYs2yAImFN0pt5er9ntU66t1yCwOVbuz8BSnqtOasnn7Yzq
MUdW7dwkoH1DLE5EsZlESUbdfFK7r/qo0FeUeYG/AGq5txrH5e1LNtA00sk3OuOw00zx4SXqHbwb
gy1v3vlZy0gvmH28kdPTyjvlCx3IVoPsM5VB1Tjd4AC1SomcDDY5YwCSQvONrHqnNyscP1/2ZhZ9
zghGGaPY+2mItJZk8iSOWY6hnwv4VKpYeN1MiB/SxX2r/JxJZ/7Iqb8qM9i+gOzZs4nD+bQ55aYo
u20euJ+pHgHACx7vGMHwXdJIYxDDTKGJ+UrOTFbgIx7ccsQhpuPu5FZCNJkf81PCM2Pa4AlNNgaj
ac3g2zk/XW6XSuaPwgn+HyIr+l+gX0sufMXkuuyZviwjhR3FIkgF2X5gVfclcz55QidZClVJf5WN
M+PEzAaTA2AT5LgiE7Of7AodiDfG37OGGlHw0WDAMGlZu1ihiJTYNfM8K2atoWFqWQKGoNsnwAI3
qCJIth53zwGJJbbnhTA5499q+BwLwHoeXYuTa1NPri0Igm+JLCmjgICQ3SE4o9e28/fV06Uj0HCr
OWo0J70EepNhh3iNxUOON6z3ltoUezx96/D5O4F48MN4yNmv2fnUZVUzfEh+CPh02rC80oDOCxhH
uySC2m3KZc4OYlZY8n4mQIKFnzqYKzwK1HErjJTXZQ/SgES8p2B8QFqwb+yNxjFQi6M1rGOTFYKF
QsUCGmEd8xS0fIbPp86QtIZjg05FUGYBe1juttea6VBRW8WKr90iA1wZSIWCKapUmlRoYBnFaO/X
5YZ6FMLADuJljm1tcSc8tiohwvaCHPUytlS/zqszTcFkgRZnzrbx4hf+5Ul69jqHr9dmXBsL73n0
9C0L9AFc9V7qGJD+UV2CvGB0UIYOVfEXaEFGIlpmOhnFG4e6rjhcKDR9VBv4DqA6m2MVK7f6n4NC
VCamk3tjHEPDLWnUAgrckbHy5xgxD1sVZ4PEeaB+iXwXCCHYU3JkAVgWWFSKFHnLcW8jW+7R53ZJ
VNfLhqfOHWKHV3xnGx9wSPrdDX9I7CjOyNJp54/SFtzQM5XbJqYffF53yceDX2iLuH54keyATtiP
5xDrWUFMP0hAiqP93FHaSatf7veTUPpbwwylaZUOGyz+nGj0cWFht5t2D47UcTFLIMqwJAbanz5O
V/DU+qeJEkIYJmCaaERJ9/23aGpS6V7hnYLwOTHw+dzknrPJNsw0ISNCE9Qmmbfs42FmN/gj4vph
WyVzzbUEltOCAf6pWZ8CfRylyJ27ujbDFVw+y0TWA1CBggIvW3+aLH57SNDMsivXytwhoyN6Bwww
RqFMELu8nPpcCqBRQkee1MnRiThI69M/nI57vfgMT35Uw7GiwpOTeIwD5KexT7gKUIg9S2p4ky7U
mLsxtbDnmVfvC6IauH5MnmBbuvfZ0GsWxDDRbhRW0DCyF9AXA6ZYdvzX350Nzwq1eBoANhP1GNUu
ug14eF5NUkruHFyWaEIrzwMT2azukJst7X2pfOfH4YVMusFkwkys4QHrW9AfQUAkU2JFvgrX2l+4
x+Z0GAcAeF5WQLC5F3DZDl3Z/5O6Xk9Dmyh1HaaDVwV0MtXSFMAO+eIclGUAoKNvQIf2E8WpJWtM
CdX0shJKdrGuZhPlK70T/zycN/ZBswaFO0x7S9ZaU/LrgNb8cpvaEq1VNUyVrJgeF5V95ttiuATj
4fCQCeoIvstg2iDDZ8F/pj6FwqJcRWJ69sG46pXesOhFKsTTGuBhYgZLET3GEH5KfmAfMJEdSizS
Jc0k/FS9yKQlcySwZmKAr/6G80YcYHp2zP/bBmBGOahG8EfcTXaC1t1Kn4pc9eRrKNx1uiDWjVPD
avYrRvW9u39i7OHoAWWp4Mg1CNg+khy/FVTHBw9GBKtKYjDsx8uo736VTjqXtT9/8FTstjF/Ahvm
AUghMYF6W+6mbklIcn1VGiQkl/zWVvWLgDBN/GW1WxPnRk/OaUzeXuOf+6wshFCeqk4fla7pbAOU
QekT+09x1q1wn4BQqaiVTZl1dZ2CTwUGQZmvysEMlPqp4esfPcz98lZLoQMShqjtHUUkaIKgzWIW
WZ7w9j1vAmBZnosi65huvUD31Pwpfdvv1B7EAuRzbSq9cE4Nk9UrGp+lfHh95RMcTKlIfv6ACRLZ
mhwMf7+EArcSxxssiOUszdPRz1HHaWxorEBQMoQsxUdFdC5l1lJY1Crhw59qCEm80QeoazY5WeOV
h9OvFX7O8mP759zgglXFP7VT8L14w65iDjTxeHobJfrk9h83xGUoJ+uhxVA7cWp+WPKl9XGX0loW
XuiWukLwfDkuPQnQayusuTXk1du1wwbHOgydKcGbf2amS4aNyLAfx6hv8LF4VacVhU6mJwS5B8OP
AF+sTWz9ndzezgYyJFw8U4YuZj/tgZ4AOIB5wFhrpzg930mGf/Jp5/H+leXbrcWc6cjWJTMa72iJ
suuP4a9AdtLH7IqQHBN0VAMuU4X+gY65uS4J/F00DT8RuXA9CG0KX5TfXtA6eFVxkdmEAQXtHq/z
mLfDSBfXmAMWzObvzNGsrntR3kyYlj51f5as29ElfNCw2Ds1h905K9Dk1H3B0n8WunP7VeGJIGwn
9Ep3o+jtTQjhf/+bH0YQGsxwzkqOBkna+nZlcai42AJnE90AE6LL5duteZi6fwnMnfiMb8pI/1pu
RwvYbYMvYM+CFbYagAXi8cxmNAit4HCT3YnoiVh/Cp9THGWAR/j4PRK0o96wOKOiJFc2NE3LN78+
i7btEoeSv8EMv8KDrI+H6JobTlKJB2Eo5NfMFs7WU131f2xV9ji9S6KnZdvE4BYCFrlLviyPrqS8
c+Q4D/gD+PwEBnBmYdhvWEpfZbV7xkGeI7pBAYXnq+LeF2b0Ci6PZM1OGVC5/7Wl/6TgsmhJNteG
xU1y2z4dGJYL+OH0xcN+40sWh+NSOkqqpEIjLJqYTsmGs53mopyHUMKxthRPsg3NVAHL6Jl34YO5
6gJYzyobFn6jvmEj9QbFogWqbSfz9GWe5rR1CevTl7HWbCKz+31XDV6rN45JghRJR29BOsdxJ+OK
o9bPK6IlGZLFuvGi+Rk01pbgIWFwf3v6psZ0Xr7Sv0OeOBdYCnpLN7NcKppE+Nf77Qxpq3gY42Tq
vKDeJmtEG6vRI3OfVOVvvpeqYDCWiWvFlJrEKXgwL5i6ugiNGExzGggMyqfK39hdWQR5UuftNIOp
eiB9+C93biofDQKiZqWKiJklZnNCXa+TCoA7InRUz2ASryvZG9WDnyaKOabftTcEOb5llLQKSvdk
yxDVwgX5flp9iYHpyTbLBMasRyTr+h4NZm7juWS64UZkv6HX/rhHUESuvPtHkB3ZEwL/JkhRN1/W
miPSj8otMvc2yy6cBXHbkVaMyqVJAQn6ypa/OOKKfZslqA1wqjlMmoyUK672W8MhcHqln6+As/FY
d0mEGWB0ung7mNRbMgQ2gIYALFMWMqnpsAU3Vu0QkeJvzMTmTGEQ2aBfDBKS0dDW2nU3N7NsNzRy
de8m3mVv6P/zN8MqOHcpPN7Ka8DN+AorDAgBW13LKVCdDjQB+FrJrQfpCunUVBMPRVsOPeqCm/kn
6BpIeBU18UWFcUsWugZq85uIAXhG16UvCY3WKeOhgKnv8sg4KDFjMuahviwSAlRyAayBAt9LKnYK
shIo3rUp7eSIpaZPRqNf/nuBOvgmfuSbkGCs9EijnI9Sr4OPkus0XcrRqvBRa7vTTJG2cybeKReZ
cOEC4/nhPyE7AYSEIAlgrPx9C1ZE2v6ZXGT+l83YbJkiYVSAuGGVWiqJozkUWkLFZ4HCj5iEjXac
5OOQRi4Ml4hfJ1hG3Ja37J2wcVYgmBq1VFCY4GYxv1iZqntrNugS9OHPhB4KFpen71hiFi3PtoJY
1k2pCBX03viN9VA/nTumwN5epo9tTOZFZxHpWLPJHlBOvxdYHtL+rFuvAaIIxq0WDDFMueFKk0+X
mHnzqsWCWVLS3GrA+kbdOJS9nzL2E1rcBbC4pVRrXOmIwCJPtsEw12+t5XltnpmCiC13zya43Rxz
Wlhl681YiRQShD4benQ4KdzR4g3k7X4+FckQ7dNP00aXMcq2RVtL1wMLjjn/DjetGVjNMcvZgOsv
bkd6I5URiwYBo6MqwyHjtX9msZxVlldRx5YsejXPir7Srb/mp0l9+AsxbuNDWLo8pQiTXTIUa8zD
klbQW/+CFqJRhXu/vuNaCy1C6vIrHqdqMdVfrOOC0fKSInHVZ5hPa+Xgd/fSnJDEunF/O4mDPzIa
CleY8M9y9OesMzlP+twUGXtQ53m5Z6aUZt8i6rkMa67UJEYrdx+fSaxTmN31g7ovRpgBGCiAUORg
S7BCgJ7Ix8gy7MQgAe8aga5zBTHDXG+JnpjdTUX4t6NCimBHMR4as7Kz7GnRA8xBv48vyUxfP1aT
RqgvMqbjeyVP+BGVydLkHAN5/n/KdxY2W43NBavHcckZuF7I4rH5LODMkF1kR+cU/IhM+LW1Iliq
O8vi6XjQ93BNN2BZVy+jIbeyeCL0t57xmw/U3rCn4BU+m5ccSLPkiBZYNXxqZuxpQEh1P0xkfcTS
Y80nTk6TGGlm5O8XXwucwz5xIsms4xFQqJxRWyntSi4BSvMvDmKKs90WfKacusGzvuhRqfdlkeSh
+EJJysvqcG8KKdmmRhFgkjZU/v73QoKEw9vZVxlZn61Ms/0iGplm0o4Xq46G+dUwIl0WBj5GzzOW
Awo1g75gC6ftdd7Ptjc+M9xr6het87g7pXV7GvtOAtwpRT5Xf2rLODamoaS5O181rMOfzniUkPU8
0GhJ4RPyZISde+MC3cHwdW/GwXyHcC8RXdN4Z6tQRK1ktbWfewSHf4IPMi2E9nrCK94okMGA5w+a
Cm4ZqdH2fJr7c51Lk9srwoZaIt4K+sVFqK7lEQYo3ZHNz43vJuEYQRAONE/T5SRaL8KheWTKhVzM
oPV+P3I0RoXfApxMefM5ErtbohT4cM5SFjzKezWZwr99kD9izms0uCZNV39Z7veG54QRj213gn5A
wgvOf10yUWLQQ4XPWZU3ym25ls/XM4b+YeVaasJTqjlx15IbpSffnJ79uLQ+EtVkinA/xeg/y+sm
ohIaA4JRK3/VXPDKq8mQdy+HCex3/eMZ7o14T8uCRTwQHYyPML9LKhMJDH6PthVsGGVTmwN4PU1U
jjd97TJdjzvcGXTtr4ZcA0eweBsy62NDnI6llSwXLSRf3YBR+xh8YWyx3GyHNhZEPOBUJRj3MRPK
0afRpB6JosrdY/uAejl+YE1VJn0RRqcL01LzY4C9kHNFkw65VUFs1tQ8FZQCEQGkUF4nbMitXt3H
JSaFyOQnfhMOCrhbcfRjxfg7ysVq9DvH1WObWh3eRzGiI4XgyzNHmoboGQkcO3ui65pDEJpz1bvI
9CDMJ9oUZjechZ/5uFyl7fgarmp2Bze+GZF1M1iJ02w6BzB4tBpHgeS5CEd3H+iE72DBix2mHEHL
16ZHvbawfcLNJRROh7uAA5byr5jVmlW2uA90yaj+LMWG0EQ30Qu9paPxLQIZ61hBd+QhmtFYwgyX
CZ63Of4NNUk8ppuvkG/a535eP2++VV9Lo3skkMK4hATpfINEm0/BvZbShWob8ElhmotjK7snqib+
64efxfNqGMghr3Xd1nTaWRvUTF/seKRiT7GzGw/RwLy89uRVmWv+1tmfYBMfFT4D+vZFIRpIZ2rP
L8S2eNGMIIRZwvVhBbtlQ0iXkKB1UJ6I3kvPdQ3REm7Yn8ZtSqJawvv3hL0ASPxKJHgz4t7+4CY5
Kv4SnM90u+HsKUKi84gd0nw1rV28Qc0WuHS7LqGDRYENqO+tCy+5qTA/5E6NVGopcCdGHpaeUdcU
1s7shWyZ6K+BcJ2ZwMTtx8PdMlccwCJfz6v5q1f4h6jdHcfEcGnfc3ucipUeFd82rgTPygsQN9B9
iKKN1AOLPSigYY0GFMLIw4g3drAO8dOQiKuuYN+3M1zeR5Bu+oxc+72JJj9ME4Tp6uFs5NKRFvlQ
C7rTYetjkYOgNgIsejQ5ScD7jelRuwWklNR4yF2R94hgBrBfFLY1sYca7Betsmt8nFFoFkvywr9e
MCtHEL6LIqXGfPoKeNXQuc8KqqGLWsEaocM/5e/qHjxSEJjxHvAKZreQ/WybDZiEvcjcC1BvqiK6
fIqm+b5kaRozLAJFzNBELDzFGcofj+v9QQ0Kv51AX1ALosZ64N0cIGAK5iBuDPtm49rcM2BtHN5K
sE8KnVX7t+AwWHPp144FdVAJxt9FkJYaxKwdUMT1xUZ/6FVpQebVdgm29y4dI1f3ylt8+q69Nwnh
aowJnF219cZ6U9VfueOmmrqVGAAH5I7a5zJFfzqR5D9zTxwenEtp80+4Mgcf3QIXpv6TmZ6e77K3
gdw7zz0LXHJkPXdoZWb5H6IoA+/YugfVXijBxOON2qytLE/vmImJDvpBLqYwXQByFduIPiG7MGj9
dfT12L9/vSGThnwPsGI6NXHCck+8S4J0vSPLIhiQOVa6hTtkIZW1oKL1fFfTTkxzlaFg4hCBXKQ/
1Tu/NI+f1GtJKksHttGAPjHyMGZGGanuRE8M3vhfm2/Bn3WTk3SwC0KEwCNOssYc2QP+FSZ/rzjp
x1YUVOAeoiG1caLb3bWHTxfT/CJlc/mmz/j9GHiux3TxyGXi9fv3Uz0fpCu2BS1gu5wGuVe1CmMg
IwgxsbU6dQVq04elzVHxzwqMAP2Ia9R4BQXK0VjaH7km3hq8et6t3Xkv+3/9oMdqctk9VDlxvLrp
qT/RDPEqWUBC24bh8P3POluJpjxTKki5g8uZPqsXbImPVT7TzQc4G40QF0CsP18h6Fjf1uWJD62I
yqcs5BHiL0ukUpPgyhDeBGh5n6CtSYlcVdVnN7FbNYhc5PME2KJgi4rn7YvwcQA9OAI6hzrzMB/B
165sziP9jEdYwcRxX9L4Cgq99dA0l1we6FswHlTOCWdBjTKy/p2gQFO8eymX7Lke9rhHWqeBZ77x
8qz5mI5Goim8iK42Dzyx6UgOVCsrgWUQbP/TBsyph3SumaWlBjiFbMbKfDilPUCbHcX6fvVk/y/+
aGDJ+uVK1WMRb+slZPCbVV72WDDWZUdPrMpsM59JeSWFMj+bZ+IC5/1YmHRzaFZqmLu8xEggMBEY
dLPkqsXa/OnkjdF1gl1NVA/4NyBrDo6EFs9dsaiiXEvi0+3LQn/mbRONC0paCd8qseMfLkocALju
w/MyT9fTa5ofPguj+726jQbKAhsjas5SJSZAp08ddupKEY84ZzozGnUruK9ouv+Tc2JoNU5JXvzg
Ki2fndMwx9pyc+5tjMdBdKbD31FA5FRrPLR/u43P/pNPtJoFiHaet4f4+Qe+9ECMS5umdQ6tJ7i0
hifFjBOUQHVILFoylnGS0KUMKdMywBwhhzSprxVTeWbdpp8/57lPakn7fByoVrLi7NF7x6eD0mwy
Gq7XASn2kXBT6AD5GcLKe5QBi2ZETMtdV4yUG6HSOaa6vwl0CJD/EoYjxTf1Kj+5wXhKYn61LLm+
p21pOYdWQWZoOWunUR60ZeNTt9otzSQDRROaQMdcKfwiP4t+8oIauPjkOawIsYFyz9YbCoUdmxoq
heAUbCZYE37SzkVvKRU7NLGSRLutpIirkj6dD0m3m02hKD17TKltrIM05PtKJZIxYF/Z7C59MtEE
oP2Ac5Xa3AzGYpslVyQR3OkqVfkr5jzdwiH9o9uYR3zzm37f4sn7UYvji78ggzPX60RJ0wkc6eDf
rkVZiqO4mFbtDVyTrXlTdlLb4uH3mrWFnBpbt3KzIrwhrLDfW1x8bxF9Yw8irKwucBbs6NGLCpxv
L58M4MvDUEa0t0Ok9PLTAmrQmJe+sXm98+7cCeqPs0wxOXij3nrfdTe7rp56AOL8WRvbA7Ip0ykY
0PlB1OYfWhIZNtATeDMy6BQSG6V2KeqyGQj7jwuEhHDeH5AuKxmRCREQJivA8bMxtZNClFm6X6dM
UPkrs8Kx3W6P+sdsYTneSx0Teswt31a3/1EDI1BZWQMdy4Sn06GDjp2kkhkurbefR+fGZHk/8IIE
1DLbeKGJ0QK//AY2VfPbjVZ+mxHCpab8Wp6gTIMcu84c47sTnDbxMMUtMlPMrSascf9Pi1T9Da66
uDzIJg4fMksG3v9hSKwgS3BZs/VT88r5mGhfKtLeCWrNwGe2FF4RTwc+kjhG4sMCLXwMUzuI6JKI
z3Cjuy+qJeAO+sf4AAjyVs6pGbTQTNTbuJY1c4iJkRWTfBQOGQHeckBWwSb5cVc3e2xEUZewfTOW
0ALW0oZmmvJUlfxzpBEzhxUMjDhLCsDxWBA7hjR3yvd5M/9/VMBGy/Uvlo9nNW2a2aMOf67d6cUf
+bP+t/sXp2ZHvDCLRXR0OCxwF+IbRmyrP5vFZIZTXm8N7qqRWZdIspQulTzzfAG3bGlrHdI6o3q8
vdaWd3Dry4cUrrDyqhJYfcs2LfeVsRV75ZqdmJitLuwbKxHSFHmmVWWO5YRZ/904yLAL0KZ52Uw3
s79vqPmbpBGe7zivkvLyrl/KOAM+V2KZDEZvH/bIx1pBd7Quqt+HbXoL/wQtT3WANt9INY38Te5Q
8aVOyryq93iVcZMSdFvZnnzjQWuRYFGeZx6n63j/opRqB6y5hwBXsW07kIgd75A7hvb8mTQdl9YT
146z6NcgCb9x+laFV1RSvHm4fUUXIliU809r/B4vcJdxb7uAAWswmdPJF+UNTbvxaeLquCFodimp
WGsStgL8zQAQJfencdd4zph37eDxiB7j8LVovOctpvwtZ7L3jWfrun2zKgbxW89e1q+Yz5s3lSjs
8jbe6/WMQ+ORrGTRrBfXVTcXfmFqjVFyPpR6oo5I/2SGkIEmxwoEnE2aklX6X9qoo83n3KFa9xtl
xsZa/5DiuJcKiUxy/6Pf1b+2lRVUD7d+dKsVMq2IhJtjbVihYmC5ty+Hw/iHTCk/oquBQD6Vzfng
YU561iE5ZslJIrUQB8Gmdn4PliunxLKGUmRKiyOKYm/9LIB207LElajAnB7e8EYlwCLM+ZMguUYm
hAt+9ySxEHFDQGZNU1eiSzXYoJyRu9FhYoCt/W2EpnRMlEKEmgJnk9KGoLTnVQHekykOc8Yk9c4Q
2wbrthVFk4mdkW/sjHtrv6LyodESHWAGpQoYXD5K5PMIcXFM5USE+HWWlICP5ZNK3NYtXaX1xPVt
bnWYEKPaiSIl3GSmjCYtkILfRqaiyTtDYDfCsyMYg65OGAK0AIRbZrtdYpndhMcPIW26IOjc9ijz
pgtdG8OuDZoxU2B+WsIRb6aFgZRsrWRBy/raGUFhvUJwerLHL5C+uec0J4CPaC88EZw7cdFcp15x
sRDbFZGIbGAs7dAyi0cpNVKKgkm+i82fFOBmEpzL8LxA81q0yZBzNHKs2hLzLd68xHaSnGa2hYXn
Auk2L82zK6kcuWdCVqlb8oLhTfNPt4o/iCg473JnLEiEgNvkeJ1HP5olQsiK5aDbrLAigLOdXlzQ
YjBAYvFUnm8pehsDBOq4TEh/exWBQWnzqi5nmxjr6okZOtxMRv5lriKocFk2zeo1+2LBUsBAWTQG
ns/PeKWJ4Q3DJQ0WSBjgD5b3NkJ+E54WvAQuq/imBQYNm/fYCfYxXgUdYnIKIS3jurzD/sLRKyKj
3j//QD8+54j1YSw0DYeo7lKqNm8RQQFytHgcUkizwBzPF6xU/T4HP2aF6/nCCeocCrXhp71dHa7V
fl0uN2UwkZw6oh0RluAaSHs9LyiysdUGhkxQ016jt3OGbj+ZjiJFw9LRcW5h/kjNLBRp+ZQNQoh/
AnXL8ix4sVxYPbiEDuDtSTngt2k0djwbGK9iRsohRbyhIT+ojePXqvSze4nnze2A2ojQK17hi7Nj
PTyXMHzzwsF5H3bZC7e9oA8GJ4ro8LviTd6pVHi8OoYdmGxnFHZW1iNUbSH66wB3EzKY7/UUv2ZD
bGoHTD8qZIugzxdUaTb+t41uc0eikiZXJAJlEXPMcxFIfCDQmeDCfpnhSx5jw9TedgjO6Vf1gwkq
mt+YbUw6euEGf0wSCTcaOF5qB1X74NHy4L9pE5dH2RROq2waTLOUtsXpn7zZw3t3BDfypA8RpGLH
Rv40o1LidrleXyUjDw13kdR8sfeyX/pxgZEibfz3ywJHy/0vUKHwPNnunMzSNGRvXRYsnTyx+sKa
TC2nyvkqdd/CID6PNBEjQ7jkkO6bfP82u53T1PTgTxd8N5uWkffkTlWSpknM31UKA5T5kZFnPfyL
1wxCWYu2yaE2PNrhKZuQpfZrWV+aBODZ7K04m5+XuwgP5DxU5VLC0e2V2hPaXkmpdWPG5nQ4Bip7
vHDso/Xqiyen8UvX30vnbEJEooUCAj+RDPLDOT/TJdRmhaE2N52p9EyAqGGlEj95tlljlV39tir/
ORBfijH19gHqfNmeZYYMRnfBBz1pjkjYOgl0YAyhKB2qvvEb3zM2Zdj8zI6rDrglDgF5za9NSpeM
7ILlNjFrdMxgvNJcAlJZHhYWOFYf+GFzS9m602U2fl92cI5jX+KVlKCmVF+2TUjHWKQEdfqeI11j
8va4z6udQUGoxZUmHzc4hmEqMvu6RBBiIVv0eY6Htf7ew/dXqJ+OkxMVzIPe3INGfp4/UTfwNyyr
FXW7JtW0TS9LEqWvsE39j4FedjbWKQkJ+fYp7il+iRNd5d2QVWmbAFmsbXoGzm8JpdwJpGB6lo1s
LAK9ZD9batWLkQC6pDnmdNi+mym71d5/zoqY8TWUzuZD56UYtgsy2R6qwRWDKopwtuKFtwGWc9kk
KNkVDKOQLUrSKgNNYCkTl5b0IBc0HFptTHPEzZ8tOXBKDmwTGLKDrF+tweNu03JNH28rCOCaLQ4i
vhg8OsNd3ItFVAPHuGvW50cYcbvAq5I0XeKDh9rcLfZfUTWxdaba/qFuqKyYe5IAaxeE3n2f48Cb
BxiOJUp5S97GzyxlbUO9sfsLt6LHhZ+zlwGp1BZRYz94bYrS5sbirR0VUZ9q1RBNiSFD0jZM5nuF
KbyWwwLNToxvXx8ZPilyvyIF4kbyk85Wjx5uhpXSpp31ozK2JwYaXgv/xw7hFxljcUJl/uycez8D
oMI+t0m0hlXMnUqcfXNt9E4IW3ht2NkFNJpMWOtpT6pUa8Bo/0tG7cHl6Pr8Fo0YNXyZdzsmAyas
dtcClSb4oy/wMteB+uv6JpV79gEsvwNKoR5irf6lvfPlPOpEzwOypouIynz8bBX8Ssqn02m3g0Fa
IsHSiQ/bIMz35S7fnUeHOyapKMWlwYXK3l5Q/bTv2GLHHis1F8fy9WGG9Few08G8PJecVzzySHB+
B8LSn2G/6SxHo+A/F/BlQuMfPPUZhVyBBiQ5BCDnger13dKrscE55LSPx3aFCestL1r8JPE3WTCC
oSfLa9sS4s7G5PxoG3Joyv7+FRmlSIVk3cs97uwR2KYylIu5MejjS56KCHEUOw+OC4d/EkE/pzju
c9oZeClZvW1t3A30p4YKZ3eJIZR5C4jMyDL2/VZNpP0JJS705QlwJ6mU97h5qwKl1zJZrNAHD5dK
ucpnNtX+2sxxX6hNdICLvz3F9zSrdLLTaWFsS8Jww825bBu0yaVUeohzS9r/os258+quuZuxHz4Z
EenZnSQJWWy+tSX2q3798CB2YrFTpMM9jYGSF5cRfljOc8JqZP2ZE9F3vLvaXE90Qq661tLubVXf
UeoFX8ylkipLbJUZ/IBEfoFtz8ULfz0Q5tNkFXA6bzcWeiMO1MkDlXUMgm36GhlYqqlKPtA784gu
MgUJYxTRUy6oHhvKDBVYxBNnQNPS98qGD995RP4sbKg/1GCUNbCVlKx8iLYt1mVzpeiS4EbMHtLU
C4Gfnasc7TA+8kXS3RroXLoPUuxfa164pF74rCfjYyNTa9AkarofCTPMv4OldlGUkmYV8eYGtNru
/jYw3B8vmnDs/y/hrron/D5ISmW+hH5aO7YPD8ZnOGeIJXL8/A6nSXZUPjglh4nG64M6tlyKvnwr
/t2t5/40TE/UB5z7KaDpVbASDFPnh8H58e2TSeVsx0Kb+KjFm0/DWeCEKPZ8bZtcqcJFh556NR4j
YqkyITs5rVuuf/So3MUTnBW6fs6peSN0okgQ4/lz6mMhU9iJWj+BU+7EwsJoV7REoMuJtNG9uMF9
bw5SwDYfMXa5P4bILQ5jXmxaDIw8TUydTuPuUWyiwmZnOnXgTaLWhVzUsefcHageAVYLNnQAllyu
EXkClXlNkU6XoFaB1DhRttgvWtn5gnfVqfYvOjifmKer5Ok0WoAisuAvj3j7r/V3HgZ35g5pdulW
gIQ5U/42PlucHAGD5Djv14mDWvIIasfghrm2zjQ2NE0cace6Ru067r/aqsnzGQff19s6FdtHZhUD
QqkjQMVeGuyFaVzXbn62pkEefNJnkRqL2ZpLZQX2U7jsm7fsTa8KznhG0tJJLfnPgF9XyWA8SoEd
JEjaf1ORd5jUHe7gLv4wajFMZ92NRhpV5twevrqtQcS1fRrQhNb/X2AWRY9BtyiVzSfqkqLJn+8O
feF1qiSvDjcAXUK7+i35M0zuAmHKEiil7hpQkOKavp5tC8dqe12+slNqDUm8h2b75Ibzp9KDZHjE
C/CUB1SwyltuM72I3eq7YXHaIwWHwuDTDOZEd0enp1qOXOI0mPkpy6/AZoVYxCGQQKD3OAWFgye+
rPfI3MIW6UGS5tNmu41fdTvovOUNQqPqRYQXuhr2aQpq9+2vxFC5YPJEim32aegt3cuRMx310Bev
GJ5B7uspx7sLoa3FIexoCbgL4UL29B3Ba+VJcVKzA6Og5ayjFBRGnFmrj8yMTc6jL0Zdyr8KPyXl
+IZN9n66EYUPgbLUo2RM2V6nfYK8Fu2iHpyQnS+rPHGmL8//2cjY4J3bpzV2C0UIC1aLZihsigr6
UUL1pFWGv9Tes7YqsMLZ1sMWqDnkDSAfdq8NbdFkZ9aWolikgzFH2Op24BFQfecL5N6h3ufbX396
dQry7bwDZnV3qc0yO2znP5fuRNywsFuWvOVmpy6StWKNtiVGzd7h/SK+RPkvgg7cly2pgF0JQxZK
h8QnoMOhzZ8DPYiEYsKO2jsmYjtCADWg8r+ETfYGnwEnI4ZJoQGpBwZJ61Qc/mBHCC+F5xYE0sKl
GhOahHDZEMcZtnqbdXumkwx5Rqs/g2KpUhE6156Z1gpN8ATCwtxqKSK0Vfe4UuauMyEwQ53Tn2Eo
IFYMBGzMG+O4jXwoSTslDM+6XZafp2375+IyIM9fNpEY2HP1N8WJtDnsbZtBpbB9ypYKLokGoknX
+I2DB+OQ+evZhXlUXXA7ESMi1mH55i+dAo3of/2SIEI9ySFfbtlTy5QDekauEYt0d9D4Fv/HqgKl
7s7Rpz8CuI4cZup23MtTeeVvlk2HcZl5XjGYn91guOMW3Tl4KgCIp2hT03yYCXPCMgQbUCAAUwtB
KRq75fQAykFJoMPmXOJdHG73ubkdnUuK9AbXtnWMkbrfAhZ3fTE+qFBeY+Y7ireKbUq+/KrQvuEq
hX38r08Q1KA3R8b05cOGpg51XA5ssJfKyN+b5n7SB3DT2xElt9+bgPoByWAkuswRU2dkVybpyWPZ
3Sc8HJwFuUaJ8d7xo76zFIEITPqeZ5+IY4taHuYA+GB33RrS/9bUVJxchWD95MhdQTTjwUZa1ywN
pka8hXoRoudHtYZMuT1OcAjZbvAZK0AeZf2a60GAk+AnMxwfTH+yhpnbaF7D0zCUMToQq+OLau/u
jc+Dii5/razbXi4gJdYLI3QnLst63KMZiS/xjsMumjB8uFfDry67ZRGAKvE2UkVbiY8zlZOxnjrv
Fed8IlrywIXqlKTURdUsGefuwOlMkTg1LOxYdK9l2GoQvrR6zJKxIoeIYUIH7GpE305Y25MeoFLY
sCPcfuKHpnHzvvv90zocO4lTzczgi3TW/5o6vvkB1o5OMyKkOWic1GA3N3fzTcgKl5Syd4YV3N1S
lxnwmcQip9aWzNHX4R4gQuCtW12M/FbpTNpJFrNzRwtQ+pqNj4gwgWQmcx2i7+0KhTvwxXc0oDFR
F6a/cTWqBOeBTazUMI21ewHFY3ZeKrIGGaM09OxrKl6a2wKAYvDug4cYb9410Xonzng9TtNr9pAt
RFKwgVVqCCtt9APIUggk0zHCGNGtwJXIhOq2zj6EI5ppIqJfs7PmTc3gOs2Y63Gf6yRUqjbT4nQl
DkC7NUoF6Wax+x5g/NxX1KHwib4GJ0XzYVLp0uf69MKLH6rP6qXWO1AO3uhKMf6HFPKWRxyhwvVy
4xTxDR1c0RYp0hdDyhOfJbFU9f23qNJ3i9ru80j5lscL7G5KFNtBjUs4VVuodEEbaXeDS9p7XcOS
TXi4O7Fr1ZX3CAP+xKKhYlqCFSk/N/swnWfdu4tiNFQ8H/PvNePJfZB6sAyXyIOAumLYfoC2Uqhe
9Ag2iEWg+D39BqjHqDahWeIOvl2D7YcbJ0ilGakKv+fiZHtXVbZuLv3r+mRjOBUT/Kx7ohDQ+0Yw
r8Z3X6IvnNrQMORzRfJ+DmpG5XMG83H6xhpTQsJpZp3d+ULN6EOVthr4Z4t63whEGMlV9jzgpRKq
ODC5MT5oB4Jw5UDdEbw1P+J15Pems5ZFuwjc4RUYtV+1UA9rsgWc/DfJifoBXf8K1Mi+kW6QM7Ul
WCbqDnNvlRAbcuQ/OpSk2fBPO5lk9of/Bgwnto/KhHZZ/zia+Xy3MH1+ZvRInMJ0QzwXtikhvwZE
MoB4NSCsjNZzPAPPdCDkuC5g260+TUKP9jg8W7RA3Ev/kKoe2gBTdf3wEStQV3goVmklvxSR1PKJ
0FxFx9E9DsZkHwvIhywdLXcBgqZ/nc//lZMvQuquU/vUYK/3d57vcxfFiFVOqlAqPn/HnXW3Hf/n
2f0Jp62gLjZHAt76czBLzbDrlVyAqClMMYoBCu+HR4ag+9rD2BJEvMIVuo4kVKJBxz80wvjD0UE+
6SJhvpu2S4Y2FB/3JlrGAJaLEL+bOrdqj7+NDkcBTw46Visvvvi+TKsJdKIM7lTy49Cvfi6EhJHt
oDxwkiVAeZzmVxTgRSdgfA+pAq14hYJxeCsRYAesaRVFN9usTGGyf/hIJNV7k+Ae7H9LRM81PO0s
MZ3YASSfoZ5OD1DVCGLmdHz17HkJtDs/bCHxMUhBRJumDQxbhwNK5EfqzO0DyK+c7Vzvmbbb5GeP
RSQw+sgWGyY08NS+7r3/Y7UIUfhbcs+5WIodhT7AOFitb02d3oPgJOotUKYiZXnjVOCdLB/4cy8M
7xwgAP7V0ckZzod377GCg6lBTvt664aUwCDlbnsWUfCW4IDeY/YDkjU4WuW9+Q0v91mI2t9LN51h
8gzb4d15JTJ4X1XpTdu6jmrkqZz7HgO7t+SeL8VSlXMv35h5OhwW1I/gltileR4U463RJnmwUvtb
CVgizPeDeXppnSwMdQLidtHyTKqHFK/Jgw1mPDSPNNrjoZeD3K/uy58RU/w+Fmi+67gEl1K1d3T0
pNdcPkN6Y4Ac2lNaBr+rXhhrYUWHOeutY/9rltQfjIyfH55g7M9O6S0VBYrUTidz0hEWA0HDtFcd
r8QetJivBkKq/SCUwVNLIBL0cjdGUuyIaw3IvudTTeBVp+dfCkXku3yu6SKAtMXLscDhAsy6VRMS
Btw+ROOsJGo6jozIS6M2+Yl4epjLkxJqoswMRX27qh1+CMQdvcXFLHtfRu3TQP2Yhs2wgPPdtcrv
Ks2Hwkyt/tUCk321xn9myDlXDYLRiH4qjStvpWL63/CLhph7WFFugyNII+wugft59+HaLOXuJap1
x//9gBkhwZIZmpuzPHgMC0P8XP58e3hIYuMSFRBLjVN4dHCb1vWDqIOjXukIxWR2wyw3f+huSBh9
IUOh9BlhLZyLZEr+HuHvIapnsDSaL6ufxp7G1WmjbKtn6N8LzRCc8j+4lXRPvHvLRWA6IRldc07J
BFmcJ+DR5nKDaiFzhqvT3Ad/N/k7ArIKziawK2wgaIphEDJPjIZlZ9SssbhLb7LbRnEb48d6KI4c
KEE3/3ErMNFP5iibWmikD6F0i5jpBbslRWOj4GqFgyplF+XUuvs/SQdltLepFNYRcObYVHVxeJ/l
GWecqUQSTKTU9YVl2dC6wHC3XMwv8zweAVSiKgvUfBVTsn/QHT8xJZkZqwNwp5mF61r1I2majU4c
EbwkZFxS+OByTiUHVv3y64euQYYwQt1c83hmMWtc92xnPJqjsoJLzHwG5FCkTh0HexpTr9zUSQjS
iluTf39KOcKQRcXc4I7xMDGV31rPUmdK99/YSvnxYS1gVZjWGon7qfb+/hAXsMtSzxJq2ayXQUf6
uhOPNFmeLZQcGCqXfb8KnD0L7jI7xlvycjicG0cQpNekWQf9VmgK1N17ZIIiSaVhRhpt2Jo9Td9d
ITPx9yW4v8Ew8mYg2AClbkA5ffYCkWufYSYuWilIrmZRKv/bQrCW7NX53tcCru5RYdhkDY0L9fE3
RAagj7dp23/b1XVQNzosWv/MjkseRwt5oA3w4KQHtZf6p2bF+46gRsIQqgzQzFelAXU16yt/u4JE
wBih3/AuBd+2/Uibo5KiqtmL6jrEryJKRnbKP32eh/nysLw74eC/UBLtaZ7HkqdsIEiM5I6wr98A
qWA9A3QmHXE4LXYgUNBbaSQm9MZT1WTVdcVH4eP7wDHzRZbq1WH70+e3EEMn77BXI1NMDatH1dwJ
pV3/PyNauEIQhTZKRNT64QRXqV+ooNVRXl/zrPmgcWXKY3fAMgkMkOFCVIgdiTHVb4xCtBfzdvK7
72fdgKljDmNiouUJBJQ2HyPD/ZcNnHc1aSVTUKnaH1Gy2huJuSbQkCTqRtXa4aBtLxUoXl+yesld
bKul2ewkSxVVZds45TbsV2x0Gmg6eakAIaUkSxl9JPr3FERxWy9OE3yq5S+5rWqk6bd5whxLD2t4
M2V02rd+ZszlUg1E6u442oume0WOyOa6UT801JbZndAs0JyP8k9hkz6XDBwAdz3HadFpwTREt9o7
Z8EIjJGRZ906xk98LD6vfNeVLiVUk7aslCzGWEvJCh9hvWYKDtsEFLVOV5mrKHx6YHNDHHUeZmwL
xqCdIUP9nrQSrevH4v0X/YnABj2vU1m8RV2DRZibM05BGD41IwxXw3x5bgb+mZQhfpBrqNGvPB2w
7hHd4YLinUdtVz8POMVAe5pDj85DD5bGn7r1t7voXyyo5ymjofJjod7gTalXI0pM21ceQIE/42kA
eYS0HmhBJL3KCmh9sSVgOG+viCJQKIC+zUEnRrwJyJe6U7zDK2CCuJYgiAYJTgOJILX8rPMAJtdf
Ma5o00b6ZkXEj1o52ojE2PayJ9TkbgTIuXnyYx/8xdQloxkMYMr6rNoNKA/XBeeYpKRzbRB6q7ZH
Np72kRq0J8qHSl6gPpagSJMsejWjA18PcwCECL6YttSRoA+99XDq5K/NEkaORgubDxyJ0/ksBzj0
iiDmI5OyNgTLaEHF4smM/IaECD/vtfPzzjbJ8toOF7x4GVcLlnszLRmBgmkW+69oyRqX9dlaNAYg
X3GxUrIcusTdffrE3i7hXNAKNCZwLUoUm2I1SQuBQIKSsC4KaNpYqHH6NHZDAoJBTbTC7q6q3ziM
+UeRYgSY7dxQyKzCSs3ksihU1jyPoC9XAuTvxMtglDjtqSytGmPlBZ7D92r72gnni1Svq1DzLECY
04IbHCLMX6N/zXqZ2PvWkQvTIxws4vNTLzMInJXFALum3vPpdVQWJc9hm9PScOz8nP1BTewlU47R
IjfMxHEiAQulITuoydKiQwUvj7k41atQh1U/d7k4S0EpgRbr6K5RHGXOJMX2V0S62fv0IIGMjA9p
AsZqea011uRPN9IKJ6K5qzv9SxmV1az2u577NTDHa75KLMj8I7E2PBzlWPH0zevah76H9AbmGHLm
Fu3d0TR/CfceoVfJlQoVz1HLlMBZREwaZG/7OfeBy48qGs6vbA1xCL/A1Yneo965z0UQmvwR28+m
vLgzG5oKmiytYN3sqbUFaNORmro7Que9mFdSppQmgp7wsA9u4DcCsLre2bR8ppN+GpOkhIyEqQLn
ksY0KbrrVDh1vVEUhoOyXMrwV6iuw7s+YrpuehxiSVwFmKYhwdc7pSVA/kQx0zfGFcUIU9/3llY0
0KgMTU/7nvxJCYpDZctbiMuRlJPzhN6fT2lDdE9L4x6moGmOZuCvGF2YtPV8GRL0kEbBnwoGn5tf
XfLYNZs2ycHd9O7MNYzAYn0CSjORJabC0w8MCKh6g7lCM1Tv+RLEfPOqm8n9qWPDLFYAKocH0UVw
MiMk2oInyor9ov0z5L77kvcOaj0x2kf/3nZNgvTFNjKG4/zvKf7hof3dSYhyMLUxQQqKVDEHjBCH
Kz39UwyEe2gi0et/9dS25FE11edMzPL3gDT/h2Buzr6idysvScfT0kJxyFTg1GJoq8ly/xIqVcvI
5J2MGJ4GM3089e2WbWkjpkA3qiU+b9J2W1yzKq2tv75QY5DujkiPT4fIQwg2CBsesXyvjwbCX6/l
bLLH/LqigXnNQQrI8cpNQ6E6Ywd+Pm7f30Y9m3ckR+nqFsso88TsEvgr2oF0lO1F+DTMSMO8PabL
x3YB9q39KtCFnPgFevzBIGTVgMdyeEcak8OTAmrppAQ60Hxkut94TgiLHko6CsMGJqIuvEPnYMd7
aVUqBO+mDrU+Jt2uiVm+6Hx1WqmF35/NZ+Fe46CX0qIM8DDZo0gM7cUeeiqTfbhUrBzT3WrE/coI
7HrOGED0f+MJgYO2fBAITdGp6nDtR8MqAgbRajsTl/y9p/YUehS2JNpR3uS5W5D8JnKV9a8i27Bi
iWigF9po4EodRD2QiFgul6e13GUaG1l5vYUCJzSGNdPHs5py5VdfwLTToZeL0ESlVy0Nop3UUwWQ
fFX4055Hfy2XeoxtXe3f+nk2qmJ+fpgWE5P2dXbxe1fkz+C0ejMzGmAVmbT3AKrUAJVwq4v9riSI
txP/oISKBpqKd6c2WfocYmCQHyQN8WYE7Z7K0sSS0R7ry9aBY7EweKKMpaWmxunubZdHM5dLoxZ3
EasP9w7v3LBCdtBDPDlQggwbU6dODtxI5i5UJIqyl3PngrYBzQjZOpwAgkOW/4rV4UkzS9wqMuBX
DxYJORocRl59b2NG5gHocdLmJDS0iVRe2NuiuAphmdpHXZqlR8JuTikP+OV1tuaBZsWmVszXUUXA
dl4NPkM1VsB/6uMqxaX/gMpTruKi5R6x73wGs6HlnVYQrrVO+fvvST9SJubchKjf8DoT7PBruMj3
uUbXZrC5ETTfsAVrrjCE15F/+9W/rYmP34UD8RBT8BjrWj4sPcV+9tipOdFIVmYHBQ0O7pAHkARM
KQUfJnQ5vvYcEkhqsAGWyWW/A7sVfp+8OsgvCokA+oen5THE/WuR19d1zZZR9T5jTG3/LHWBO1os
ro+5eSxvc9pchmjGUsq7uoQNDn48x8fnzYqi/02glLjzS0vui2H1aXd9OaaTIr7sbbh3N3dv/w5A
C7tdjEfmNBl7W0ZACZOGlrTK2zOxNTwYmOxvzaC12rWcy+3HLIAtZ4t8YmGzmh/6YkMWHJkDk+WW
HoxmRVLaXcuipVy2B0fvhdxo6vxiOc1fg49Va4yHJvZEc5nj13Ng/GmiQY+QspOf/XGU684iUHN/
Y3B1G82oCp7IOVN921M7k1NsRcUP/KiLgCIgZjpz+tXlNQ5OOMGuiS+Kr1qtlyDAtdjb469sIZTT
yXjEToL+hG32h4D7+/JfulDeF64j1JREmgcpV0BBZyEKftZpEdCwWTaIlzNJSLggUufvclLQyIou
H/u+nfNyzbVuiXD8cjYPnqbUZcRkxGjjQVHBNFNQBzUhmaByzZ7uH1vrjYlPelbtHEbCqW004SeO
f/8rM+oBqZFOuzKCoj7iheEvltxkbHayUBakbDNwoprno7Kk9dN6dNwlAbFW0MgofzNSpV44nzkZ
DB0tKAqqLmSgrZUr/w5xR9RQDIfa8eqK1k9Yo6p1H7YzqcAj7dSgRUt1pjLbbYUrBmIlWVzAbqf1
a27FNZvKm69zOcZY+ic5ixaYS882BvZVq8rXJA6oyzjCK5ORiY5pcIKxUJwDIedqlH1pgnyWXoZL
OPRNv4BoGuasG7h6nXrnVmhexR3eXhmu60uqhETIhZYEv7JElU6+eDnpJcSK0/w5QxBYaFK9Ssfw
ucQjQ9okylsCuv3pj4Yy9LXlSe6Ty9U2oCmXrr0Xkur1J3ekjOu6o4ERV5NFNIWbdvthUPRIESA/
MHK7HKfbUz2ni+0kTK377rPTZ/mc5SHIDLncXBNzLcXs4exA+Nih0SeIKJvpyne9O6CKqHKkNh9j
bg6Eaadec5UAeXFmagFP2J1Ksowy4Vrs/xLF7SUwiuVY/zRfgz1Vm7O8N92NEf4Yf7+EKWmIV9FO
eWNxdTMQTNkm3ti52G02kzonSinXD1/1xTyf0yX/m7SzmKQ61dkWdQt9L4gmVKR4WIvuFEjife70
7haVzhoWRoHPMlze80A78YN3EGrHkj3poqnCXElfVWsJeQBQr/yGwSbxNqvDbvcLt6ic+UlhDrM6
PLMAacOmJhmeREenC5GsvYkw7nPMN+euAqVqUSgJhD7pjTXgr7EuvIHH7Ip56afPmWGpfq64RAbI
5Sp0Rm3tmtEO0p2I2iHR6OPedSGTy8F5+O9z984FRqyLIIYKFh14GrQwVF0wGhLufcS7kVaMn4x5
NaohBWmSog/SkEV9DC7DZ7fF0m1aFOtTLvUc9atTytY5ZdwdpdoFYZxO8nfLSLjkzRzw6O7/KwjL
bVK/doYwS/4fZXlHANalQ/22UJ0Yg5wWpwuMjETjrHfirMkhlzy+8kUCJbduOcciCJGDz5WOkwOB
0r8GYUhEZtHWy2fMtSDeTq94TjA7AkXCdGCGNChqZdje19vWtrOlfvt2IpLAGDzzOCQvDaPXWIuU
l1Yhy3iwyKLFLwvWSOlIQD48tyayiuTCP0ZnycroERQnlznbRpWcnyJJJwzzNMTRLYLYr4Fc1eVh
ILDo9hl9bpw9wMISwEMfetEwa1wCO1ENn45pNRXvP7+pTPJyO2NL9xCPmgjjPMED5bNqCrXcyZwR
j12v3ZoexWWbnrvBEWCk/fyCZ/YU6kAkPyjpQ1tkHq6PgyO/deIwF3HXohFATYUkk97FIF2hmCI7
rOhxdWhtioh5Jw0Pspi9id/mIkdsE8I3n11hPtJ/g8jDoBlerODlM7uBk1kiwbgq3CfoqkQqvVxd
ytHoOuQrQo4+u6YHIx/sYD58zdN9F7b4UlwRnLUBwnRXEjyKeraVKxsRVMBFMWBg4nlABKOJbpyn
wjCWM5Cv8cMmvvUwBNn9p6JDLR5GsmlnRjpXy/mCSd4NeuAKGSRjHECQvlIlRqX0j8nZdyB1qnsB
ITYx8f2rCBdw0n1Rc/MRw/cyVo4OKeqMk4qYcxi3YPLTzCfvf+xVeYMUnDjjwFHMsGFtsGm7Wdf/
NrNdORWLfnGf8ocFqesRHHWEBVfm1elybIpvPfEErPXD7ieOj5nIcNvD3J4AHdMgOaR36SRL9UZV
1cbrQTQ95RQSj8gmDXCDuJXH9RX3ICsgfSZaCcgryJxf+aKU9lYEathkI+kqpYWaFbuH1wX3oHpN
FJpLqznGdubXyBp8hJt/UeP4MOF5/zVZ2RpCzDX8ti2c8WxnJmN33Fos5TphP+ydhdk5tSJghn1E
QP2eVD70G86zAWYWZ8qfP1SvHedvv8D+G3JCiWPE4VT8NXUv0Dofd4FSQOrpap/5CmX1M9VqVlLe
K7cKOXCKWdcIsVmYW65i+j978ual30FIqXo8DiWrdkayGUewd4k4mrL98uEwgyeBdVvqqCbH7oQZ
BnrVNd0JShLb7LrVJr51FWM6X8djymJsn5SOFcsiXJI1K1E8qBPYMg+r7Ymt7jgAcvK7YB+MZD6F
iHjVIHcUllFayLFSLpqwPCe4s6uO++unFZsNujQaowr2ecJcfgQLVbCtDCHdzD+sIrYPmaXDR7ML
5FmzN5pmbA+semFeCA+v0Gb3cK+C95shJ38o1SPIgHpIZ0MTOXa0yhQczev48bDfisYWTa58LCQE
yI9o7s4I6Q0JZNhRlrYIpQOmFhnVK+CpiAhPfk5dFi/E5HBji4UJ/nZtfQljCb/b4ubi2yv9jNQ9
4PqDPbgtG43n3uwoXsFdB+snCCObV6+qL6TFqspKCDjJkOuHDh4GEYrZzp4jTaVCPQpHiRJWvN0g
Ekaw0UUQpA6MrQEi0FNkyY6bUdoxYvOQYzbRYklwU8PsHni7gWQtlNzD6dJYoxgvTiG3fSjyL5wi
CkESqqC3xBphHNxNfipBSKIhmsgpzfn/zFr6o9OHe2lFXfZvKi76lWF1CvpkOhG+UPRWfv6dmO6R
KmFGxhACbdvb8Ic2Op3Fm8TtCsTf8dAWHPsX1Mvi+kctPXT5+8sz2Im2gjc3EVxOVeJL9lOADGXq
ushZtXZVsTs2A2Qi2kheFg7cVWi7Ei6NFTPa2pZdR2pozEspzBTEsZHJo26+sm3l0iyktIa1ADjW
BGX9zSPXcOWcVLMbyaCl6EqvlAe2Pf7yPVY6DLihBPALS44u+CpgBiOIiRxfLfsORjWZIrzuDTOT
yX15vbviaQgwibjmKluYKay8jNzOi8dqWSCBddT8tKxNfPkq6Bzn/sbEY6/mpyCXIucCgBs9SLKT
4ErL9g9/p9H2HOMmnvDpZkKjp2+rPVGKAAH34iPATsp5ByKr9oCeY5KcnilSLWbi/u6+tKkmAzdV
jozBL+eZ0RlQ8o04Z6LONsxbous665mzsXKZ5oKA/ctDSi+hGEJEdxUmIb1pe6g+hHV3zooj33fD
mB0vS/GpjoR5woxjAY+G1cOxOvJWBtCaXeVHqPWq+2b2YCs1OGt2v23fMsyZ1XHJR+jt+JUF7PXb
Vaz5bBh/3fEoXWQ4FcPoDbckvb3cqDym3WW6yZ3oJPtDEayNUv++Vo3HhbpSNPF/vCtZbCSmdjbH
s+yq6p0wnN4LPWzXsuC8lH59yo79dsnqb1AFuZpJSCEOPF8vtFyfIHpOQBEuqt6urXz8CSyeUteh
WUaga8sZsoDhoxKX9Ra4lPR2f9QsTFg77P9DRgB9hfxbET/ukaXAW/nHhWPTDyuo3074HeCuENqO
SOdOcP0900lWGo+CBF7C+qPi/9/EK6J7f5GJg0JHyCENDwnH04hDHgu0Qt1dzxyf0gDja1dhsP/A
RQuAJq13dLtHMdzpmh5Y8Qs0MPLRnhwit2FChOZpgwyuDEVlkoh4Mqr2Q/lEIR9etDBRvEKlo67D
r9m78uTz350JwA6ItcGQblh7BtIjnWN0EIGA3MJufqeQ4Vp021xU+DZCul4vgwPUSMXmhK1hyOOO
nI3aDEw2DfSa39Gvak5LQyHKo2DyFhyCkW6Xn9TGhqcIMIsf0hJpfsDjF01VOL8xB6FkVf6kmvo5
2gpXPEqMYWnpCR/DxtKDMT7vmu42N8BwMqyvaMXE+lz+1DTHb+uKUNYp5ZgQE1OBX1AKUR9+WFN3
LitYyvNd9VKrvRussTvmJlDz+XQ3xzqpHLi0SJa5F2CYn1XAyfLYscq5pw9xIc3wMG53SiitE1xe
bx2lgai42u4cKGoHBQYt3ttaYmKVpWRDirqyW0ZgQw9J5DWbCqHbR4jRVnVeQCqTc9yQY/AYmgXO
CbHEzTBGo7eCrxJ290GasRz1Idy3vyfB8tkH+FvM/DNAn28UeeWLUaTmrF81WfuiHyqZ9Sq0ne0n
hxgfW1MssGwI/G3B6JxbjZT81rGb0yaJa9DzK9gBhF32PNSpebT3t7sWfcuwyO7kdpKYu0SPXE1Y
3gYtE6F9I6ZLHjO11G0I60cf1W3Ty5nrYuAQUpNhhnsziePPP5f9h04Tau8kDZlKGigYA/k27md0
n4lIsoXbeUxZ/a2gmMZo4kW3TeCKOxEx1d0UsVx7RWNzAybWr3c7rInbSpxjAUBnSOU9+u7dPVRl
WFJQQ5MVRT7fGyI9dRqDRsIlZBA+FulRRF+3F0wtmJoeh0oEh/Y3nZY2l2G2gpuLi2N5+n2sT6hc
tbs/XJglLqp8orsVDRJ2lngCWcDEIX8SyJk8o75XXpaYSZ7kCT4KngmPRaM69hCbVS2MF0Wu0mJv
YW6bLH81TN5yHSF3UUfYR6bDMscR6iBBdpquTQq+pfhuTD++E1A0yw22vIOtr7JawUmR290mzQJK
Hjow815IIRFKXIMqGL7n4CCP0Qg2KfaEA0Gm4eNUN8UKuWHAax8PmXeQJVZ9K6PDEIVEHqROWBz3
rVTrjsTGPvnNWMVWXn2nF0mwl+4JgIXSw7YEUsZ31l716OfiPAkjXp8+w+X5I+vqRIhMxHuWPgXd
wetDmcGXdqDcy4o1xl1b5sMK/ORgj8xmeii+9qDl7GJ14dJC9mR+Nxah1rthTvUH7FjXE/103QFe
4DbqmZCjI0vdGIr3jAmo+V8q90S/kb/LGSwYW//fhLTzyq1k1wUj+vtsujyLhlUEib+t408QQeZY
kcAT0BgDmLA/nSaqKYlWw/rL8v4zyjT9mUGOBcPbKdNBL7MJTLr/FUO7Qsrq7J4sPl0nT+J9tLx9
GlqGVQdgfbUsROxmwYIme6Po+6Y+2SZ9S3o6lB84tYHDJxEz5ANLjfX0LXosNiItZUxrZhxTvMcE
jhcr+wV0jZsT+rgcEydvdOYUf87EyjBakeR5eAufT40/Mhoz7dETfTZPpxp3jJOr4j4EXL1hIJUV
/3i9ROOOJziEsWlib+cgREEkgg0F6E84DWD5aYVf2WnwB7Mhyn3bNwlUUT0uww719eGgRGE0ip0B
5RPM9cwLMxiVVhNOLfueqnGp+ptoqMJekSOHBinYqF54+XZQ6py2T/SGYPz1i/S0gGdu4qiQjBoY
oaJyftKszDNC8iAtZ3QlwkFyOEfiwo46J0Nm0LuIT6aUWI9ea+F7K+b3/zj1G+F0gsJfefUufXON
y4ub0ZP+1AJcDA/XLW5ITMRdwHdEe5in0l302hUBTNeqAM85YYeb4OWmTE+Lz8dtQR4U1AxqqMat
DBrj7rExImfegrelU0N8DxQam6kIIxUFQfRQEAOvyjmMf5j537bns+WVVcSsb3ZpC1uNi7E9hNwE
Whrcp2h0FuibvpVYI9Ly9kFhnN0IbrBGGie1f5i/M0+ZDkv2+wSB5ITIZBleJ/LwQ9gAghBiIbW0
5Eio2JodxxYsC/lnbFLZtpZCxqKj7fUWO4cwyOLcqMS/JPeWCV29gKK/sH2VJzUt4ohQwPty2o4I
3ldJihRSbnBb2rUdzbibD3sVxocnw0eNWYhuso6J7U+aclLjRMBVl2CpD3MgzVTZlG3mNx/2PS8o
71rnJv/9dTQPNo1jwLgZ/JxqQoSYrbIW42bsZ/Wt8pYyMv5bCoVDJ6qs3FpiQ7nQq3cdbxu0A28l
WAzdswC/pRKiJt5SAqq92bXElimBQIO5PUJL+4qkoypTRzJAiGo3pja7eq4X+MT+fQjaabqdpZXY
8QCwRxzFBgVfoPVqAgQ1OoxC5F+sxv4HMgvt1UDrF1hPUsU+Zog2fWIlA5aHxalREwe89xJS1aW9
740Bz97r32K/xjG2Lw6RQMGRGN7CvA6BUnM+A7NsEgPzidvPACTq++SEg+qUMfo6Wk5uNrAgOFfZ
lqkcQpK53immaqTx+wdToQRySsH4tXh6X263Xyf2F4aLZne5m8xcPabIhE0/PcG35bFRwFx6trl8
iirMBUUqREiaRiHV2LqMVxGTECcbKZqx4C1MmOp1HjjERQQBnmQh3GMSN4nSCe4x4lFKbw3dgXEx
+Zo15u+apYaJssq5uw7lOeCO9JJiSz35pTbGofUEcY8A2JCtskT/iMka4ey4Hj7XS9clJyfSK/cs
j1GHGXYthcwplp+fwNAOTJRzakQT9XafL6MZQtKo/Mca3oNgkXj0Mn/2xgYMuCvkRBLoVnprLdDx
SrAy1uttY67HOrQzJCgaErwK4qRkO+reH65s//BiLv7mdfu5q+T1FMLK9SSRkwQBHR7Nb+v0A/HD
zjx34Z9lKjLqtsOtjHD1silelhx9Zqp4UH8Fsvw71uX82tUS6ACAstEyBovUA8X3hhwuk5DPBepA
AYzhBgu5PoTwbskUDqMfK/ZhSr7Afp3GfpXn7pG0rZRLB8tV2h17VE5QmF/tF7tONqw+vjqxU42R
hURfdkRdAcLj4cCVI2JlRNuLOPbSJ/yvY3o5/qAU8N4wiPy/ZzjNZOI4ijnSrjX/A+AtzxE+ijEU
3pLnphQdCtkEcBJaHvxVAaWWHMiErRayAA38q50fTpLH4d+aTibQE29ggZJwVL7kt6iDdjUJ843S
/XZnhJmHWXw83ZjLoNj+P4FIh3BxxBq8MewT9whpdt5IzN2L8oRTOCh51hakaGJ7jY1NXORxiE1J
R+aRbkDTkPPGuDVDoXR1Rqvz/FiPzyAh7surNB3MjjPqfTZSjt/heEHtNSr+HSjhfEbjtiU1hV9+
jWzE1WDqHimHMAZL1B1pq8jItn8AJAmhuCPx786yofQjKfjfIyZ3nKNuM063FnrCqVCfo86lxg+C
DcXVwCDZ4PXIHsB9epHLlRenA6n8RFsNKvY2/RVjl5kxpBbiBXox5pUakGietAliHuoz8wkJBqaV
lO8t4SEhFXK++Xh9qAet68OebDsiErCBfyNnNML/YQlXM/GQoNc6OxUiVegfIGBz/sG96Lyv3C8N
KOvrvbRMBkoZROut27T6lqrPxHaYQmyS0ZWyy69mwzpaD7qZr/DFftVx8GX9PJzKsFVteQtFmwej
c5PNaW1pFD+PqFEENlQ4xLlBjOO/NWJhHoWk+xFok0o4eHZ6DytmjA304E3lQ3MT4ARAXJF9xslH
soVLvKNezDsfdotMQAC2hG3y4OmWtJXmuJ8oEy7xzkqKgzXXVi51k3ZHM0a7ByfZubRaZjBHgdpV
HBiajISW8SDarNODtUASMkHTnGdxXRFLLcnEPKeU1srbFhjb4y43+kXIhef7YCQYytPtKCUH4FZf
yY18VgyVxTj2tq16VXjT3jErFMTGitzrMbouKa/Xif8Q9ksLZ31Z84wDtTWdTdRXZdcuRguHjhz0
OtnJwO4suwTUCTVM0zgGjPHDXKhzhmyG6Zs3qQf98NoeiA9LOZuqyia4P0pwRV3cm6kzghrmeTyR
CWz4o/uoz7gPHfuW8RpEmI7aCMK1LsrbR/wTX9grNnSYb98zO37JQjYEpsTB1TDsec6fckXRT/c9
OTpW0ul/MyvIswwKqhfLv8tsyjy4YfmJzQZqu17UDftbJPk/Q4RG3q6V7xXFmouAJg2WAvWi5idB
/f3T0busSW5MuwGlGs63opcSWyXreosq80fDGf1g0rZVUy0qqlpXmwszPrDiaylKj0NOFkqHlQXA
knT04P9MTA6/gdq6QIZAyLaY1x4J9YvkS+Q9QgxFWYPazyPZXUZqsfa4MxJEvfJ778LJ/2Z0prx9
3EriqR3WEpHB6AEDWVhnDuLF5CvF+kMl2ZqRdBRlOMDS0dDPYSdrPvBqQFumIOmhI4ASXAQ4rCIe
XdT1BEQ9sBc8w6hRSi/pVaEVSgv43sr2M+xjT+Kpgq4P2FCbD3FYaydIA/i3u5fexbYuC1pX+Oyz
WjBkqyq+R/NZeSpP/CR5PSZmP7Yn6EBEBDOl4NcNjgJqd9FhgdBGdXvdrWBbFyNVdQHTrkejgeyG
XZUOz9sCn0I/nPIEWp8szQO8kHt3SqDZiMCzE3hf/1M+4+s3/3DtdeM2xH5O2Qx5Bw6Z51LaaUXt
4ZIBW0q5+4F4lvW4hWKGMnPxqS5bufipHytReeEMU2biWmaZ0B6bcpJelHO4+6sB2ZRYiaOdBvkV
61i847XZU5q1E7hFZ4KQarqfFmuIg0af8PPKsqsVZQtf9yjNFkbAPROxVQNzArzbghotvt2jN3DE
wdCXHjeJHvWrIB3+e3h04xVnGxxdfiiG2YylRixc7g8oDlVQ2oH3KmNRU+QfSLc5/AoLlJ6KiplP
Ktbin5/Z5G38dOdtG4BiGO8zQdmhk3LcCEiwde+Vy3tbxqrvIIQkbAoYlnqCEL+T7F8kMS6EN9EB
3VtKig61y+2iFbFpbK6di9ukpCeWgw/VwPl2RUD7hvtqybmFsbumYVfi0wrKZQyOV45EE2N1lnie
+TDyLu2EPMUfnp30OHg8tUapCAhK4rDIV8audqxAiFJUWYeOq/C1uCSi+qzr9o02qlrjiDjAEi8r
WEvgQMmp7cnouyZD+itzHwkz54HKV7CgPINSlLcOyWDgvhfBGYwRWSNexK+PBXUpPVtXhjtsU/uJ
YGrpb3LNLAsedJ98vS4LuBCvsGvOWKpoUK2A82cbDBkgkAQDbgi4wXhJEBNgC0jhrsylH2QU6kyt
5KaMLKVwmWm5CFmj4VitiGSBD/IT1p7OnHyK6xoI7LREyiS3jRzueKcty92ZxHgDgGo+WY0k73oG
r5dF/HjZzrv0/c0NGCSWqtj7TEPlgOeqJgponWwnZOApff7VkLoWrcJrEx8ucc+AXn7RaScwXVmB
awotwtzgxZshNUXXKFXrsuxIxePXlSBk1BpCR0T0I6YNQmEiVi5HBBANSfFAH9JaDgnKc41fN1Iy
zlUpAhxTQtj8LVRQQIFemXZnFnNP5l1qx+xobUJdZJtL/NQzANFHJIz/15AX3pm3MThmoYiuEfER
fyVlkjKw3zCpRfr+l/R2yVRk46WmlJAxqQ0WXLfxYGEKndQ+8G96CCW87/w69F+yrrRmelfyLZ25
wSuVptSMh0U/ZpEL76Th8Gk05wWRC30y5D+ALw7y7yKmA+EWpHCDnZ4mMv3jEcAKdMPNdy6SJBo6
HWNhkcLCnKeTBgkvbjjOTcOW6b52XIJzXA3ZsfYEBsMUv3E5herZYJwfbyAr4pOExpXNHD1HKz3u
JOS9etu80jBy+kgJCTzN3jlgdARt3KayphwcJol+57LlhwoszTmMHmKLT6badY8dWU2ozWUoPUk6
WP2ojnx3M1DTv1iCGUmZuz+zBMmk8VOgSGXSuv87sU99cldiorxvJRTEXVuM0RbFoKeUh/ZUd0q7
VMdesdonuzlfj07PcJ3U3ZiBP3yNFESsp+YCzc0bHVTgYnM87ptn+DSHnd2s52w5YxTrGyNFqeyz
6R1Ly6WZE55l4TKvPoEnAOb3DH0v0xjrNZLktrxPurHnZOk6dGKTOAa4jH16K3lkuakGD+pFmBAe
UwYk05qJsvAApeOtN4lbhXYjkuhBAJ87zWc2IpFYuCYmLxreYdUUyIFJvrAg5s1i0cTyyFsugPl4
eM2SerFEmf04cGWPPTugOiCWY13jJ3LIJzEhQJG0pMVTp2zhMSeItDF7G7zwt3jrNRj+YpU9pc2p
iDCQjeP8lPV1ahvWofoe0dGkVZNy3Nj79nkaEfmSWd7wFwDgqoYaLNHLFJsUAu2lAuPkTOXKQ8Ay
BwUbFNkhQFaOA6l4PHN/IZsqmcxtuALMOpOBQEyD7THzI2JnWhMB1/57s49P18FBMavC50lGRzqA
zZhwu+WgCRaVv49aSuIZwq3GDdmQZBIio/r17Tr2GWDcw/R72XeIFrofYywbnmZgOHMUEh57kUxG
vy0dvg/RU6mGOW9sQIkou1ypT1bYzJ6o6rj2NjAze9eMoLg33I9WYCHOJOvhxLY88SnrqSWv9Qx3
Bw7GgxzTIqjDv/+Xe1WoBIFh0zzffvm/PS8sck17sTNrLAy+EkWudOn1Vt+8kmcQFGGTh6xRGhB7
eLF6NPEuAGhmcFCqAH7jLhYF8YB+od9WuBlJrKlQdiboHmKce9u3q4wdSpYY2ptrq5ng5JatLBRm
W8/SMsrCjeM1ipR8ETi2zyGJomTg0xBBBYUXMU55/7i/4N81iImy8dvEil7oxLj3egYssAKovKn+
eC85GywCcgT+IKb21txrFS1htjDBu8vi4rUVztG2Ge6xsYTcU8KAaz/s8hqnNFJPsBwxU1LlbgBQ
M9DxhfNkpglqPA6g8G4x9ccGahPPyIzRbH2s9etAmOGAJZU54cA+Bv6H7NMJTGnVcJ9A9ZGzS1bS
9Bhn0VmtFof9AvMI6RM/S+dA5pYvP+N91we5zUO62wNoaLEJn6t3+PRgB5hR8F96QCW5FVzcVl/j
l+vvlsMaaraTqoY5XKcfvnamIvCE8xMAnkeZj/wh5SY8MUiv0kpvJsmqZRugUtT1LMoKcTts7fEK
H4/UL5oS30w7DU3uTyNvb2FYviyMW4fB24kq2I3Z7aWJzetYidpz3mnaCZE8nRQvA36zTgOBr4zn
gR6Xvv0BOzuix4Lim3tDwpn9gPw4EPVhDtTb3hZz3jWCyPcg2PxRA1BJYOp1krn0JGdJwGaCRmYR
QtiohWednFxf+7z3ydIZmRLwm8NShWUjompOExA3/JBGrWpfPx0qOthUrfwHAtEXXsyGJ3vFGBHw
LPgK2auTREF/RbF/rbz+6TDgF5LlmNoFy941NaNIresPK4Az3A6m033oiWYCLqPSpA65T3ibMcX5
Ufi0mumZ7L0cZJTBVEeqNcZSty3tXhYOUCv8t/c7xw8dJLnfa8QPrCb2C0bb991nEWBG7dQjGATq
fXkquGapD03K/v3rhrJF2rnYNAkYZ+DxIM0MdWyvhVLACvzUMJHukvOXVpmlXionDvwEEhWhzYTW
/mTUFWD2SrUPqxLy8z6x9qQ44PT+Ytp7MUVjksYg1o5QTtiEltL5fcC4NIK4w0Sxsbf/RJWzCx+T
7qONSzAXlazynueeXgomWP8gd9+67ja99iDSjuoKHwFsVd6wg6AAiFcGxpQkDbRKnoPI1sGsstBd
jjA4PVKPqojtW8wSZTZUZBdxqXaxrrnadnQYTkbObXCmTCCGAUnZIsGYUVkt40MUD164L+NP3f2d
jJYXTcLT2d2qMmkeOmrNlNwVYkuJpHObMJExJjKa1QYmOH4ZymxKiUzKwmZZQdemAnvNOKag18A3
A5xD1H2SF+A3qJI/l/o2QiFWQtQvv9OzmFAxbJOnmGj5Cg/y0dcbtSdos41a2h2jGdvvH28IbgeG
igr6/dFPe/7YfieqDHvVzzzDOgO/Y7VqOM65RlJ1MbxelKd9wxQzdA8Eqy9gL7Vxzcz15mSibP0k
OiocUjbMj7B2yHnZOVnyqtV3OVZMbAF6U1tsILOdm8UxNIWuc4gVpwM2GgpEavN0XytWDr2RcPqS
mq1CnvWlbeyN+RdXeGoISDGb6wyZsjlP6MaFQZaEFXLEq36c2BkzcVhoBPw03gKkzuXSxq5SCl9X
SaPp7Beh57GRu2MJZghNgL1HfI/BGxefBiEQrDiLvYjaROHqlPDI494a5RZGwXcUk90Dta0C6mfw
nfomiWr79ieGia4lkR8byMyR5B2kL43yeBjHCiTIu1Bb5+cc1Szkj8DThtGfz8KjAIQzyun3zooW
sLedfiln5hDeqq7VciPqTCl+gYp+dXT8PvABMYvbcn+HIWOZ5nYyqEvDqwm3eTWdkBPi2xMYZ10R
2NbsRKb9GM7vtUp9LD8hAd6HVN5NpByre25+FrPiIfAO+2DQGJwqe+zuBPp7scgswIuSRRCaYE1I
jz+stFxzLA9RQ0Kc9ViSnpiiac2HmgaXG+wGHJHFP8f0M4UzcP+95xEbdj7ckj7sSIaFHgVcUpRo
yMTDSQL3JCr1U3iW+CDPYnfzK9gzMO5qSBcb4wrdm9XV74OCbRX42eOQ2Gr4aFrOLRkkFkfDczU+
PCTCFXFI8U9cqXo5PzvaEmWtpFZeNftr3VrbOeaxZgu+gFPYwWjPeaeZElwV4PAK3Vwtg0qWoAbz
dMd1wWn92X02A2F2evG3y/nLMarbDpMC+112RGx5kkr2G/QxLXeP68qcp1sOTVI/t18W51JGSuY8
AIwMxEEWilx2zm/AR4smj3qLcZjCnYLDHVKjXRxMev6sa8IgDOmHMenxq8noBtVy/a5JzXJhIa90
lA6Fcu5f/vzG3DSmrHBaLUtrDYMKtLOV1WiG0R0mzcyvxYfqIaYT8qRpCYn29wfO0Khz8Xa3XdK0
5+xL0eEknVuZWWuU83JqXOM6QGSolzy/jKxHpWmQCwM5vyPRCv3ES7jtt+VixED1htFJ5UBUUf+p
7twtnzJQOLCNvm8Kpc/7QnZj5c23aktbuvlHnRGQLWV/zhIcFY9wHq6ncydSEH4w/BLj9ZBDYVFg
DpLBjSrToDOEWvOhHaciJocAVfKWb/IQapGOzMZMDerqVOgophQrol/amGsZiHo4/qaYi3YpuTuK
36RhvWE4HsZvKvRXTUz3gF6Lw9a2bXfz7jrIIawmGVifz1FBFRKaIj7A23y2vRaAOFW6ehCSqn6I
4pp/VJWDJmJWlNG82h9odrPlP13l3xqXj2rQOjhEZShCTnL7f416MCuqOR+cgiR4Df0hLT+KrQhJ
VhkuBBWuXrMcICwpKyfEboLQZLNOyONA7kKhd+Omw6dCVvZ5/Mlj/E0DItY6oxZaEGVdEzv5GvYa
ii+bIjXWcpso7t+koxQQ8dR0wSBcCcYK9tVcWdeb68VHxWGIjQznSTWdgsF6HGwQzmXfxKZMPdAg
5UJTHaoZtGHowBx1R06OKZvAxqcJYDy7LArPaNexFH9ynjOebv6fg4KoI36CzAex2xIURYrGYZfp
HTADXj7lpOxYXZGaDzuQCSAe5paggqlW20oS1vXhII89hFTPpE12QBHxdgrv9xlewn2eZv/naIvy
hvMpwriOcB4XqyH/ZaMOG4WbKykh13SaRwxTNOqNTG2yncEQDHxZpb1TWcjNfKux8BAFQ2i/d31M
QiSHrRffIFvNsm1REbNkoEERWnv6peMzvcrXV/PvP0aAK1ZuhM57RJvEq26k1t1JVfGNM00YkPb0
k5FtknEOFgbT2M6zsX+hWv2AX/THZ8WQDztUEGrogMxV1+SqmyswmaEZ9rdu7muzw1ln8hYP99En
v2TkLhxzYwcFjDD0yVbXWdlKYkz1SUX2klCAu/gIV/8uKyh62L3tIVBLSzDIdYAyz8hA8mRvyJcx
jY6ST76NQthTnX6Vmn99kw4fIsjRA0ObJHTiu9WSoo/K2q55rwOULKp6Qjgaa264bO+hAzEgna/f
DZ/pHzznuilS5L2seJaRaD5RchbNsWAfSrGJCvuZeIRbGeXmc2WOBbrs5V1Q9A2Z7hsYwWjlYo2z
yFyVmYX0ub9p05rdpFFujir9GxeH39zcrs/zLBJ9YANeMMMOKR3W8SRt0oc0aBne6x8gd8rDwu6t
4yyhOEpkKVrd+DMX25uQit9w5+EPZ/fsGrMOKs0Pm+swoyaWLPO45j7D6KWSHpGiQWomgrku08ho
brjF5Dbnl0VRH3dReioMuIP3Qb3USwyMGwDj4DJp6PnZaQFK2bUDYchV2h012aFWEE7SMkzZK01+
vR7OFR7wK+rNlBByFaWQVZCl773sZbrcRprynu6NDaeCyU+7Tr9n5WcXcGWqFSwaBuG+/wVU3xnD
J26uLTwvfxJTxvY0uqPqK5tqNMUU8++uEqI1F5ziJzFoQ7P7uVUe9nM/I+q/UpJ6OcI3vkz3vMXQ
bosmExh1y83I0BU3SG2G7aEgm1s784MmBO8EM7jVf9tiplgZf65XERiShY0dxwpTCocTIPtBEIQc
nDZpYafEr+9BqLnPyjhgFoVElFFUIXbhFGGkkIDJl/ivHvokgXT5z4VwhLXS8lb52/TjVBGu/8RQ
+JBehk9Lsvh5kdCx5v7pVhj+pZ77AGbiXGnkQ6hj5NZCT8f5zqRc8HXxhRRGu7Sb/sZ9D3v85hLJ
LKYCuzzz7d8idh+Rtp1f2cYSzOfytKniD72VOPu2Bax2tTaQgNQZ/bFC7WmDh1tmk/Da2aRfDTVI
wb2lvcbkY+MUFZbNIQzEpG7NGlP9KaRVwHFTi9BvlGeu1h0yjkAW1F5xQvfSsz1MQ/CgCCj90g0M
EpeGK1Q6/JH65C0121bKccXi79LqnZSi9HxsLhQJfZl3d/LtggK/2Zw2HhRREpntiPpdbUhKhryI
Jr4i6VbITf0nX9jnsxZYj6fqW87YjAiLWYDcm3MtBSZAZZoyPnj8DZUL2SAJjLzLxht5U3zqaPHX
EV7zGFbqdmWczPlSfIUGJhVm/PYXnQ4h5rPZoHTLeb7Raz+pEx5oPiEM/oCtwQqVVwETgk1Sz6pw
/Whg0LNl3mzouxvWk8/ifSitxwlHVFQWJ8eZvUb99zqUsLhwYY1KsbNtL1YaNeQ9koJm87hYtXIF
SOmSr+NoThynN7pwYvvwHUf/Il16sbzVnlIifALYh36PvkXxX4/OuKHeJ65Lg2xUkFpcVZBQoq+d
yjAirtjcRkDzzLKw4XUGq+eoba8o/HOdKKCe2suDMlEJhNRx/tn5yJeCdQbpMQPqs9oSwOqSWUhm
ZrpOeH93Ffpd1z7ToJZJ4FqEhAbgRDz/9sVRiFPrwEKtwh4j8bSUhjjXG3tAvvUCIv40r10K7dSI
MH/DpL4/+rW0+clARIK0MluXzwTE+i6s5O6nl9k9e7b1E/jmCEwtaWBqll60J/WGPNwU5W0WXaNw
xFpjxKEqEsyz/OieZPuRuHCPTyR2gfrY8n6VP4vuWoc2ABF4p9ngo9u91Eqyjo5qtiQbc9IlDo9q
zrakV9kzJ6VnDxFV1tcVUX7CKIjiSadIzhrVncHIJSjLDkp5OkLIEeq3fxVwk8R6817AStWGa5S7
YHnjXG62DW7c3BMXeMQ8/1uQT7/VrwLWNieTZ7zx1QHABTanBEqK8x1KCIotjUoEOQaBUdvauEIE
0YdXhS+QyT11dJSi259scrFSCtb1K+nX5jPdko0IvaLn4s98jXflrL4jHcR5HX3YdgEkb5rK+rsx
0JsvLyPr52Zyg3eBikN6RGZD5uZed9B8KxZTd8PQg5wCjw1knFo6W7TtnUTU9Y5YxvKDv8f/aLMv
i8pFTD5sHJIYljupgQZzTqAUv7XJzeU+Nj2paNNA9gcNzBVVnaqOssGpkLTQG3wy5K+HSbFuIlYu
cuw19HX2l7bZxszQwJ5KftlDwjRqFoG9plsp91TclwqGNJhSJhnkWSNexzC2NlNdr7HEL/fHIFzO
LsHbCBXK7FvHjgz+Bjh1uU0RVOBlC0jE7sxY6hi3nh5Yu7HwFXMEv1aVtbga/mMm/bpkseZ3XbP4
0s38gH1RmhuF0/RxFZe5PD5pcdkAAVh1jxDa9Ec2xlGY9COn2WM9o7ip5sjelraCKM+ZLbVuZAyZ
M3eBhe6ikx7JLCZIL7y8Scwkp2pfpri6T//KlVK9LTZLh6lIxibwr1vQFU2agmZ4GvFNsH8N9oqo
yUV+R+pSAp2zkfUY6Q85nQkVSUfGB6rWYk+1O2PUNtsFbSpBBcx5ynNC1zqwXnu8Cbjql24Hjjjn
E0IrCuQCWJa83VWxK0yD/XPnkmOjoyvdofecCI+YWjOEnklxI/jyR2jzTVTzmmHNfuXbs35taXeM
d3qwvD4jiWoLpoisUze4REVUUfWkn9iNdw4+US4mQMevjpLo2uHwlQO/lHBwmj3CUrChqE8049kr
wtOFGOav2BTuwTcG3L1Eom66rMPhEuMnR0HIAm1M86j3pqeKLtoC6nSZVHVaCgikp1FU5hrXmSWt
ZFRTEGvrgdGSGU/xEOBAzR44wdOhw2kh0EpgjXrPIvwp8j38WsEPW2ECIP6EADY/maUw7UwgaYnT
m+zKNlPHSo9aGW4OddaBiGr0ZqTT83fVEW0NK4RX3YZeiUaAVljCeOQ1IqUHk/1abWnC14PnPy65
L+44omnUmC3+IZCNGnfHG7lpCym9/G3MKWJBjg2DvXzgpPfLMjq/u9fu320II6uWQ1EKu2fYjsDF
lCA44cIy1NSXHOryD31a2cdkDkzmUStKFKv97hcZ7Ukv/BcRR9hPpYd0Y7PEo+U5oqjI8OqVdqSh
ZoifgwoECbdTQZMLq1ZnuGzYrsyH/aSgC20W7Tt0IKFPv/JTykXAEaUCdXR/MN3sssuFhzaE/p3I
nn6lVbzSvuarzQb8hWwWnlNoI0vHOxoy4EKZjG4ml3iYtMwX5Y6PMRju3tlBmdPfUb6P7qi3Rfhk
LeWO9WCs/0I6LV71lnrsQi9iPZzLB/QzloliTI5MCwdF1UbTjwe/lQoQMJIRxnEhWK4aWQNI5Uh7
X0p/qPNCgicJAJZkXv3e19ZZbfHCnr7DJHNCOMf81va7LWWzfhS7PDRwjQ6e3LW11oq0M33TUtde
hTp2JudxTzCmQgHgkvy6MwP2OQJ1z10FRv8Mdue4/juzd0LgqAB9Ap1vXf3ARW9DlTyJmqYhhkB/
JksaBuM1UvInA+nTjUVvVrG9T2kbHuEICDQNQ7MJyoPRyU/n+G4CzACk3s0R6p74y6otlt/pT4Rw
oDKk83FVkGtLSaahS1Jv5dliDn95gi5P/txH03h3+CRpnYeY+Zfz/JqB1wVRaYPAgijh4Broe4Ps
Ft8d6YgDAlN+jDMfsG/XZH/kAtF+u3ZvOPiHlJ/tAsfCR7uaS0v/Fa1AEQnfqjyTur/kSfmKA0ry
X1PU2jFernt2wl8f8pTalO7U38Yb6rsNau+b02UpA1O9r2z0bJPSUSz9CaYkB/NVPlwayH3cYEu7
pN/JhoAIcfQCZfpz972GWZz1ZIbEBxJRgS2gwtGfcy8g2QsWU6A/qvOqkjD6MNbWV6wmWGJhCQH1
p5yBI9FFUOCQBD07I4Pn3jnmKk8K3fh0z2GWlLPuHXnQXRThfK+mZmqasb62SDWG9s3tV3UBe3yf
oDo9nSJiQ9G83QdzVgjNVyKh3L4KCYn/weGQnaQO6lmZ6p4NLF0+znBMlh34Q/lkzNlS5fhUmbTs
zOgQeW8aWNbTRgeeFyd7iO6RQAvOxhCcpD2fJ7Uyip1udJ50hmMajixP4pYzmgyUKa/U/6vqQ3Pe
KLqEAl9n3YJRw8T3TKXdH5+FCKIZS+5MJsC81hVARbTrI9fNnMuA00NSx3IBOQ9sFhQ9sBDHztLJ
lWmzp8OKrFGxAj4wro36SP6FkXS4RCmIMzs8sgU3cihJbqR04+kDwnUk5NMHKLCXNuDsdwOt82in
C9H5WsG7GvwBR/jKdt2HBTsPllHDeeWZpLEfKySRLuzipMlysKOATsTKXGO3yFzt4UcuhJpLzt4w
NZYUXkM46MZna0wNm3q97VoGVu1fdm30i9QtIqhxFzdfRo+fvH7JakzyxULMFVNihnkmnqPDxWLQ
wb50XiBzR6sr9EIpUJXAsYlaU0BHkMnpZAVqlQBAODzIKcF4MlbBj6W1vCvk1FSmEJmhnrmvc/iC
H9a1TGXOdDFxRBGCeoW53MLg0tPuci4CtBiUuH+6H4nofTDSe6ezjytqdpWZILToLQRdZL/e40eV
M4ZHxoIysKLKtmHHZCG1xPPVsK6Llfg7AmxigXdvSvA/b+Eg3zMYwer88NowjeyxHYmCkWGJIVnl
vLkM5WxpMK81ECWifnCF6JZHw0fxmlN5ikwf0tPr5PObxVDJ32wS3Yxu1FwwfOksDLAMGoRkqXFr
wB8Mlq/XqH4hnCcKeDeryPCyZ34vmklOUEkBqMI5m3GKRciuUzpUul0eVY+MklKFQjBynbfOSP21
5fJp01txRCd4Pq/GQdEnxhJTlPdLrhG3Jos27UnERAhaZt+Qyt0r9z15UZ8eTIovPr8EUz6UCyti
XpLL0J7TpYEjoxjGXKqG33U7TudfU9N6HoGjdaw2zFGl0JzaoYBkVIeVZ80Q7LECtV9zybmVWrgk
j9hhCbNCz2+CCqoz9SNV10HVO8j61QUpz5gAkl5B3Bmre1HhCKdXYTyAh/UecT4pefQaF0M1ZlEq
UR26w37DB6jvOEU37PfFurXTeDsVrYD3NOLrrMLS4ARVHbIy/Cc08IUeoEOouTaG+j7n2PkjzWyM
GM/Zy7elbasvv6Q17jEV2SrlbS1I48r+7UaBdQRTm3786vmzFpIIpJRAo13xu/RurWEJDqHN0DAY
78i+L/DelRIsj5pqS1SdS2bFeUl65tcu8mmw7NGeAESv2M+1uVMc3SGLMS2D1YUXwR9nQBRxqj+i
0+c1yH7nuOHzBZbYyacHISIHEwd9kkHom72PDqLX7NFbFI77mUCHgsviuSyXPGHawDBQh0jNgsH2
FvPYQnjDcsgWCTHi1dHplKru9hbfR1Z2Wa8BRW6GIde+4HPtxE2LJjbtp4xn4mhGVtaWvlA7hmcZ
leuL4/kkGSGPBcriyoazGEXb1m6vqZTiNBjV2bs28aNdIMBFfWfoE8t0QcmSCgHK0GGd0fqGpXJN
62N3nBFnlbn/97llBxLdgbA79wn1qcOBRwveHduU95pIGcn/UI1YXf9f09BAOyg/8LHMVq08oDid
afG9E1qQ2vFWENN/bD/n1ooBnzJh2bqQbjb+QHu4wnVEkBLH3KFcD8z+CWIo+UivHNHZ89qV/24y
/q3NEMAJZTP50sOc1TtX86lGgGMA58sk90lrqQcOe30iD2qBmX3bUnrOU2Es6H604kt9toKrYDuy
sH7YlYntCP1JvkMYsvvB/7dZTNdBsRfhC09R6hfatOcwnqPYxI34OquOiYhr4o6xq8dnGFCAX0kQ
JT/6vT5kmZ0USMQEdbjJx13L8vIsLaeaslzHK65tIsx52tCvfV9IBQzYU3RxbKgUmMSRzV2OvLFG
nNXlYGMLwg//4BL7pGwJ6DCvpzb6zxY75vGyd2rRrQ73g046aJ77Jp2w+q8bI20HopCDb3NwxjJQ
OqRX6j6Ngn2YuURLQiv8J7QX3oK0yHjiebEedN4Maph9WyZISExHOuGAFZ26X6a4iT6rcAAiQfTH
njLnE62eKyetRtAO0tBAcONZIuRHQlUvKt7xYYIH7P+hmbwG5LraPEJUyNBO2lxxefx848j20irN
GCFiiPmATFs8RGXiSM1SjgVTRmFvCSaTe8a2l0kiT8eogYzmNJ+FNf4U57nga1cYzHPf2brPCgAz
LW60+WVCLBvPOVPFhvqN+AV4Jox6r8X93vV04Z/5rue7aCRiSwUInhNKMKpTUM/esTw4fKSxmfEc
enaBMEVr5Z+XY1/WbgoM5pHqRi/SAWq/9SbnIYoD47PmkhAJsCAMASvVJwbzjL0wgBJdtexunZZQ
xllIjn8HRWPuzKZQh9BjejvzZjaKuxuLiNtlAz/ipUdQpnUxZXrRK3VaBIlyi3rm9uaGLl5Sf+Hl
BrFgL0Vj4HSe031Aae6mFIwFxnh+1ivBlIOs1OOIqosvSGB1mqTHi4oHz06sj6PLZSfJgbsOYo6n
+VZgHyUgwivjiGs5OnuBPdiV5OKHPamcB5UzT5GLD+hxJ9aqR+q/7KOPfgRaOlu40aestjXPERSJ
vn2cy1+uFh23ay+uSyzlkGDbPGfpkzS99RXA7gsY0vPrQsQKsEdP+0nAZZEwDtOrtqzqttKAeCO0
Wjvqi+tOVT+N64A8YnwPj1ZZJNhA3T1Os2mSM2Vgl3IFQRlhumdvpi13yttxA63atc4ByDeHyJeN
uHFhEanwYw7OrEdC+JWaFLF2k6PvlnTlZ8Q2OG9NT6f1f8uM5leSypVXCNx67r4ToPpST7+dIbEA
KtUEf0uEG19ArDEOMdf+nqToYJHHNKuWWFyIp5kk6g8pKmL5S1dGDl7h65TDVKZovEkjp6nR/3Rv
e/6eQ4LKFDE42tX2ypIb/P564p+oCbOdQz2TzaUNtcuAaDofh9IcACH7IgMFf+j47nqjBgN5+iYS
61SK3gy2PZWC/SqPSUVqaWciVT8CRts/N7x9HXCfmtMnfl+7PvL87JpoCp0vD+5wX+I2BWYlUU+6
kliqrLiZ/L4xq3lPKg9oSQnubnF6g2WcU7vddgFzcs0HBaPX5+vJt22ZAg2ZBg1u7TOqVPwjvBz3
YxH3YUnO9IhvZoVTkn/gnDL3pKYFXSZdUlurEAXQOoq/H/lMuOgl86ZmXHmWQj5AVtfu7mMRp/GZ
KmDsUE9GjHMccB+GJE9ZSr4/v2YsRvl38qo/65noYQ0zb0AXHuLDiq/o09q3JlLrLH0merU4aCO9
RHhTiPzvg8ujxHjRKq2mmHik+Otmbb8rKoeBY4Yi1IK8PkPCZEyN3TwHc5hmqKbwz++KdE+ywOXM
4Pm/4lwseS+tnkuypQ91+wdlWawfknGatpxSrNyja8pAzQJZKLrtqbxLWGccWmXNz7Gb4TN49rQt
2y8ijyYpDNRZn7EafmW4g3uoz+/9otPgibXXDDPOhANXMreZSLGJm+Eo1dZ2bBejOJWadqkxT+Xt
LDVKI5bu+ngOpLYJCisBlLkcRbaea2prLl/9UyDJ42FFfRoDiSAlTKNXKUe/pnmap9UO2jk65Y/d
fZF5xx1MUEREbN/DWvDffBCrXCVhkRkBQUn7DF42cZwDLcUVcEzCwdj6+1mk87LYU04hprFCYIq/
xHQBYmeTvgNf8C76/baYqZ60ic2um1hZfri8AJqQs5UFOe+Jv66PH5rU2XIeKA7pcpGOw4pWLjHM
d/xSuQDTD4gfX7ZSxU06zR6RYu7/d1/7FdBd3+ch3MhiShI1PJdHMs6Qm4+ZCsXpnHPFGQnwTtm0
jGQOsNYJGQU32hJVDeQc30+5TX3TrHlGoJ/h1179YRh6Wvs8FQIRcF1/KzuUZmn6MezCXSdkVoqI
1msJ1kNEULMo18wbOkZeUgmW9udw2kd1YBMWq52c48Ldf1rAYIRU38DRYVILb7lK6cYR7bX9rOiR
mXyexp9VlpG4HIchXIDOtSQ46/bR8TYrQfi5Wu7w63pTOsSrxmA5Fgnw0xrj+fDulAAJoj7Nqsq/
N9MlmMFNaaoNXEiILXQjLim94Rv3v8zQLK+UHRtlmcjKCQiNKslrepeC/R9NwoaZ6oUgDn7KBKOO
tvikLLJrWexKBpzGV91asZgRLRBjN00PmJpbu+l3SzjGw6dTEf5HgDtTxjaNKcn1evm4/4vZ1UFH
KZYIWTWWyWFOD7Sum06Onu+7SFs1ReKxhLC8HTcz+xpRoLeVLzSVsNqBfqgZKAPfXykAT9U5oJ/a
qPLerfDWMrINh5y1eZ5C/bjbQ6c6yquh8pr2Zoq/mBkIhmujn92tRs7J8ya9u2HKpskLYLyHbjuy
Wv2H4Q7wnsfDpswmIZzl0NIvygeRZJztsnhuUpJV3lZLwXUQQIB9X0FiJwFJJs4skg7nbTuAgffX
mnGFxAKF2vtJm3PvFvt3ZIzWc58S+Eg7Xc4mVtt8KQTDbQY/AI8doWSjDWHbvpIUDx7xYthqIgKh
5iI/TygEF0kXLZNsup27PRddXFa/TWOCdi4V6lWwG992jDrFX6xCPr30ZwHQvfjwG59SEXTpexTY
XfmQy9ruYgXmANf1JGex/10tRdO9gb4PuQ9lUPEI5ibQpXbBny5VVKV2qaIDUBKS3W6g2yyNywda
drJ1QNxMOH/tUc2TISqGquikSQjS8kYRkglxMI+dQEtwCh65U7M0qtPNF+yaGMaJI6Q5YoiVnd5M
7qa9uqe+Yz8XNNJBI6gK1Uxhshfn5t+vaG4FKzWMsBKIUDCoiElLQdtOMKzpk9s6SHT/ErzKhNaA
gG3VhbbXsFRLmttMUiMiFahsaQ0NfPOx/wZ18DiThY3KmnlWFapijAMetffPiprL+nQkRy9xo9YM
zFi8+i/aRZmKmxdkumEWfvLBQT+kCvPBMHyPHqUCpQpkle/NeOzxgiBOlOBaD+FvuSdNjW/fy1m7
NzqFkOHuh3ZPH6/+oX3LPaWdwrD/DgHKRQsEu9PSH2IGdKXUi2pKs+kibzFHMFT4RX9LO01qN2lp
CFl/ev9Ixogk/2W2a83duVU1pitKWVrhyDorVCDKnWhfIpoTIxCKeYHH4C9rxdNv4fz/uzGTo9bu
0vU+T/nKsvq7981XPF2hRDZ4qVBt6YOKSF8Ad70t6l0i1+93AoT5FSEeZi+Y/fDYt7xxYg2C5kY+
pWlw5SYI0grF0lCETcPwEBPTT9yYDC8n6D7xOWdpZSEFkiU3Ho0FfwMA+MDzplRbnUjMHOueNebR
+nsPFhcuz0MQR1gAohTABHNoDAoDkjpj0Dc3PhHm/mJe5F19Qhyveq7HHXrPJASM+6hZNJ1uExga
DQ2jMnvcFTOpoHS8vb7M+UT7BbNVJSPpWkH5Bh3Najl/pjXmnxBbJgBn37oAM5y0QkBwZA5fyJuS
Zb4/bVYse1Dzh365Kw3j8UC0EmP15TIWFjoywuZcQuFKTTqS/GBaD6FxZNtBacw4KHSrFjYEdROa
uE0x+p6BFU1lxnpIS+3gWFVAgajtUB8d+L/t6OmV5dS1HGpP3lOQXIizacNM1Cp1Z5DcTVydXxKd
PoQH+AG+qUyZuZyOz1l96M0NIgQ8MZNvZ9gvsP8ZrtZlKtC54HjwBWvKDplzZeP95wdYxS8y4r7V
+LaZlnYdV09CjG/U1YLIPBxkUFhVxxBNE84v3CcopzDCzhg/OUPAFSFT8okY1JIn+0n3SVNc76sI
gF+56wxpFe7ULEmsBEPvrQRIu/9rTXC6e78XY2DKsURcCfEKR8eyyHlpgMip9TxubNVU1hn2c3Et
RZH0Xz3UcOR2Vyna6padnPFsdEf6dxK2DaO68OOAP8pTma2AsrcHDIDuKPBi/rraGgjN9XxKlMqz
yWcan2S0weNvNdq2VYCSYSSGXVcgxmoLirRG/XoHCZLZqiJsZ1aJVfoFU8tM2StHxiQH3dFLj6dV
8cz41SSuD9T2y7lxWs8zOcoSZi3Kn4uSX3nOrC3ZYVvYi06q5ODKx60BL+3HaZ+KaZ/kHFNJvpaQ
BHnFtqhxzjodspH+MLeh6abGEimFuwC9ZaLwv71wdV6god6C01MdFcvcKoYn2vFTvq+nufsyrOl8
sYMP9eEgYnVtpxJQi8TChKwxVamvLwXoFNITvQpfmY/CnS4N3rDuCupVeJxXkXXDsGJV1h6+U82n
JYQKLZFoNe560Tr0f0gbvVwi1T7uzrhpvX2v8Y9+blWJKIPEAMSVFun3w6hvpKdJRx3i0OYvKkSz
1o7vO7AH/K3f5/0zJVUipGiqfMAAoX/Hl0No5GUvLM1W7+DsoSvYiXAHRuO02jpsHUhdxZdP7KPS
zh95obdciOEwDh5B5zJ+QSbYKCivhl8YBqKwgx4qt/j1LkfzlPrAdASsnxV9Y0zKX5lKumpJtCj7
bOJpir1ScObtGxywOXqbyxAmK553sL1nC1ldWfrVEd7YeAFWxrD9dfOqJy2GC+V0lhmEmk8WambT
3V/Etsi5XYztILLnkw+p7ESqecwUnCGu7kjMz3/YBszdlH402Drfx1mPEEAGLQEhjztzoE+h7V3z
PRxXVm/8KGo9r5D0IicijoVxo4kUkzYvwVQOhLUwtErb6RlPP39ErykuP18uMCxYUiGW3YEFq7gd
KxJPFmdZJRYkPRUQXfLWiiacNxvuXqDNKjvxujnD4vj36j+D3ZaKpBfPP3aWSoL75a1ChAnxGNw+
WZBhv+683wUpJo2erpmfalHRIwqut3mBkpwpZq8mq4foNzWqDMBb129y7uSTN6xbXPKoD3HWnCad
E4g9Lg3QFGjy5M9j1OiSqRXEWpMeDwMUSuwINHfMVo/WooFAweH8Hch7ILpqENQTg+VRWuRI7pvw
wzr9Suiq/yNDJ2OYL/wtETGhvzIw8qifMUK4Ajf6DPCn2Dle1fUjlruTXOXBrBJnluPwMJpHZi2F
Es61P5UKLNbxijAIH1V/T6/tjMlPa1KO92EADwtELbbVupeHR9BcBP5MWRaJBOuH8EqC+LAskEDC
PRAzYY0LutKGANXjHArwDGy84MGsC/R2mN4wJXI6nm3AdEUwfgOkSUL63vSMRWmGJJrr0h+lu93D
IU1tp7ILbpLmHE9l6/ZdXE7bqSheqcfQdNFrIyNy5/A9n+4QnhfpnmG2GcBhJUhYeHGrMtOXD771
B+NqWj5ZXyQoXPGIHPZfUxXLzGRn+SAESRdbFB83CiXeM/UlfsrObdsRyNlH04cere5rBdhwzYT6
9y8m1IPnSw10N0MJYm3P3kS43VCedMP5AjdH1MW9AGmnlj0AkiNEGRgfg0GlUMKzUxoUnUt8g0Hv
v6HlmkLu/PZ5d+8hTXR69eVfVUSl09cQB08i7C6SmZ0keCy0bF/5k1zfI983vaGfUZfJwMDXZra1
Q/R2VuTHXIO9eWTToUxs68Lfj57Ooxr7A+3OobTGFpX8zDTaRUeJrIgE54zz6ag6lK0fmsmujKZO
SGHcDyE3/kX7/KX656mg4ZafcwHjUEsgYG0zUCmjHAdv3fQrKsgbornXfVpPd0Y5bH4dEeYBEZ4H
ZrbgO5urJMvrRE9EZ+v0ZxzuwM2DB7TrHE9BNkw/ov8QMyY+0T4D254XMrIkanF8OKDevFmzvDoz
7eoK1Lati1loh8c5x333UgYmLnFsKAsAEj99xPPqMxHsymetIkpllcp45iDZT85zIySrWMga+lax
byuBf0uMbUTVDKYBuyve3f4i8+fu413jlFLTp/BWMHvthaEA98E/TgTZMKr4N+4QOE0/8G7DMRIU
ivft2vP4iFwsfHmK5gbjaH6KdsyctKz7f4EJh7ha35tDq0Ulrcciv85JNQVC3lECTllOeC1yok7I
k3wRKywaAPS9iqiHew6biWDlbSfyHfxde3zk0MXT9yrpTZY6eLxvI6lY4eXcr/G25tqM7iw9wjgq
7NIXnQXmyyyzTy3WKorkxM2HCtwXtHLly3kzI+6613cBonv77X5zpOEzHQiIyqCC2NTJU/lfLVmv
UDJ3rwRat6xJfI9YYBHpSimaec+Pzbv671+x/DFaj0MlTLM9YEE1TRArga2dl4Pd15FbhBeCdevC
K1w4TltzsWb+tB1qV6SVzw1RuajURLSvL0HOqfD32adXD74XYTspdF99Kv3h7EN8lsxhJiV7tkE7
B38jy8KPBVLwJ8PTH2nSSgVU/LI4x8IhmyRm9FeZr+VkZGoxZ3sYi4MG9PMV0m/Vt6WQd8oK/Xqi
Rw4B3cyTY1LoCc9g11zDNaF/wPjrSHxdDSQXmgVoryfJwLGUpFI3Bw8I5gYza67AAgzPQGAxIm2n
nOoyhBtJYTjJkMbTjKz/oIgYOmwsmsUafkZYtQ4tcP7o+a2RUC6gu8bmhd3nOTQq8deoKYRr3+q6
EcFv57h14GEavWLHzRjqE450y6JgqLZn5xawjewgZ75nObEEpWrfzLgvFCB4Ymv+tNkDwOBDNnl7
CZsJGBRPd3WfP4ag03uoJ60plXsSNy0ZTJpf4RSJb2Y8Pfz9are585qEiS4K2AHAKwEEM6ws5FJ9
VlPT3f48nbpJ3heGevJO6Qi0IchKNFK9j7fQAsd8YzUoldyRby7BPQANiNxCSfQGBKE+EbvKp892
KQtoa43MMU+Zb/zUo1ewSBI9z90vD8s8mJ/iJ6h2397VfZVIZ91/tBzoBE9qwPlXZyO+AFSSF4wl
2uOxmM3NZYW9N7HXrmSomYrFVgURRo0bdvDW6hWHf5Co802rznmuyF6vrjmMp7+FhW8YrA3Qbzyi
EETsDeUNy7ZZpCQYs0pYayxzQ1quSi+SwfU1u6QvG1NQqCucxsogoUfAOucTCkUCgPeOSZv8QnBU
vJiXEyIzUrRLKe1V488D4Zq3uPgAyEp5iNRFHFRvUKAneDDTjRQbn3C9TmM0Km+XBSm5vf9lyvBw
VDgSnlcYb/jgdYQW3p3PMTbzydG7H+ubwp5EaE8jLOoeAx73t3uNAeIGG/JfDhn88l+RDN8TSLCe
6SKBs3acOSY1N0Pa6LRCbAfZ3yVtBJAotvT6gVeqIzP0c8HYZZ9va/ulV/tuBWkOmwD7fBuT0xiO
eg4Wi62GfuUCPIaxeLisBZnOTAVe1OA4lBTII46eS2HqFcW+CRBxqLMZvwB9AdNjteUnZh0QqNV8
JsNcVKu48wal5J4RlzZPzDE0TcCAmuqIYLg9KAv4E5a3Xx4I+MNCHpsHfw4ly3DuDm9mZsn5Zhrl
+9sv8MpHgEosA0yQLuS28zqTWmevOGSNtWhF9LXrx4Xzxu/e0HO4Phou5LadQljCJDUleqdlKQAU
kVm/ebGGSjWIdWvTCn0omnAh4TAItjthnYaZW4+tFYhOTzkfGC7eFcjk9UI9dUdJSdcYv5z+E2DK
UtRUgEsP4BfCPpOgLHgXZ7yW2AvYPehyiLBhEYS8uaio2SNRMwk6p4NaMOkYgEqjqMooH/574v1j
zBN4351RlTfLSIBMKW7C+JpH9/B4eWU6hzLO4xFsCs45Qau+9P2Wvf2hUzeAUbjKad2zJhCPorbi
Y90lH+/PiQIP12POrqr8qVkFpCixQ+8InbSy2C5KvQz+jX3RzdkgYHlLMwUcB2EFkR4EKYqEntkq
XsOWzwdmneuuJXIDRb4wz8YG9/q8qIGi814jDzk3YG1FJIhlHjfsK23ZI+BW3mcRb4VWiXs4IgU1
07VzHZyVC8Vo6SaTJzicebNK0W+F+oitub0eb5zX7yCpvl0GJQ2zkr3oet8BSxpSAnBZl0wMu+7h
Mzw5wG4eR8p/S8dtm1Qfdi8hsLH+42yywPR1ZwQG8vek34ZoknJhafwN3Q4QiAk09SFmgr3Q5MHn
esqzcYku+IaZO9pnKthRJE6HWQnx8UtWH6GJ76i+0DRIbq7lNj9Nhzl0Y4HdnKNXDIzdvJHQ8vxP
HUlimn7LzPV/Q1snH/1VAIJiPdpLLuZE+hse+mOe9xrHSNSwPIrB+jnH2Fe+LONv0XKRR51eljuO
pOKW33y2f8FxkDyFKE5AGo97AyLHs4yIrYEpwBJzUTW8nFdXmy5ZL5x34xLDkcs1g3Lz/6lLOWQJ
BqbXVFnx+WPrsfFlpKr39ft9Xefw3c9qG7o06JL0JIJhTWhEpuNUu1uK8he3uFzltPiAhpKfC4OF
O7rVclrNZkyy4wN/CkQvGDLN3+/fNsc4pZsIngYdmU6yaNl88c7T9ijRuVF1iXjrytPWYZIHCFEH
ewOamgNSFNYRpDz+XoMtaeqnF/uN0L06nzpCHHXj6HFJLiDsTvZlYm4F8jG7vJdw9OalrXdU3siQ
Nrk7O+rHdB/6qYyipFAOLoECcR8uvvUODiUvYXSjrKh03BH44x2XM3f3Ak9ChxRCxwMzHtpvhv6N
jLhBvAnNS90jpprw6zfUiaD4Tzu0TY+fuP94hdpfPP2uIKMN4at8bGJn1ehWWH7mmyKat3aHSUuy
RpHT62RQZq1riUTfmTmZ+ccTrQPAywfgyDBJjV2eEfWByBi/0rafiSsbcbgGsGyqtbAa6tLvJL1l
JjPEl5UIuibWr2CioLH7+eidiP+a8/Z6WJe/FLBCeT+Vf6gAfEezrmQucgN4akaJ3dwvbOj1JZks
++vLxLycu3WORNGgb2o5PI4O1tM3EZcwd0S0dsg7hF7zBNRqLaEmSHIYZOgEdUYGBy0OwxPGaEmo
Yr/eHOwNvCeNQs4d6i0Pap+83xV+kOBzcMrw5vyv3NjivaCeaLdImRc4D62E6omL1nGEQzjifaF/
xuO3iUbkMGDSfeA1uZNPYYA3olkmIzhi+TFoTMMxGONn0jGzfGtOmvnxKBp0AoLOzIuybp2vfDyZ
qAyFcn0136v0V4ZHuNjW7q9eCHfQMYFNoZU4D1pDFJhsdwQz+4gZV5haK6YOTRoC7QBxGLQuDn8C
Gofv9z53LvR07pOSrFejLzR1CbSv8pLBIECBNpVysnPk9c7v5W+a7Wgcehx7FvE9eKSnDdTjTGH+
egmrSUGAPxZ99rr4sMFLiBJ12s/IDFQ6rYf3TMR7lxzYSV/12qGQK+WeeLX3CUdPFR07kbErHELI
GJFSVgMYTOAQS7bSkin5wgYwqqLLLDOF0XfyF1fsxtwPZh+QoR8vNqt041fqVlaLL2yiDYOuGRay
OQfapxLSK9hIbU8cg5jP7n9aG6MhAJ0PVdozwZkUg6m+zgedPHMalVPERLwbKDiH5L3rDy7BkewO
qLUO0i9WKVZRVQjD58BOaRKandCBII5Tu1FDZGLm4DVQYgwvI2vCthuSP677vafVOaGLwF8g+b+7
40RX0APlN88S8ZtYJNgRV8yECX6UrnuH4XS6TQyPjW000mUE9ALuhod0vhXAhwJTr1EzOkYsdGN8
w9NFD1OVxdpP4aUf9ffiRrF8FNU4ezzDepYYY1stRVArvBRFRR489h1Ts3CxuO2+wom64rQ7pHUs
I6o0nO2kf6/OwtF267jFaSjtARD4su2uLhWHFB+JE/bHkvdwMtv0nbFXZpDzFtencbX2NzbcxSzo
UKMF3XJ4Zof6AsjtUGkJGzZUu5Z2KnXt5cQBfl6dcXMaLCUZc7A+HGle/T50emzdlPeXa0RsWFJK
7WUO2g0fgjVdgCOceFZPyLwLjuiDOtafWrU9KKtPckMadnCcteSPve4jbJi8cn4nW36t6M4Lqz3w
fZwjF9nywG4J9at5wgPP3pPSj0IwNK5XgFqXzizQUIlCnr+V5fAOx60OZU+yr9EIW6lyGNXSMym9
XcnLFyEQ8RSOkG49arl/OFS5W1uZ9NSnQcflQci809rftLZFJy7LKXs+o1gGls5owcjYRx4FcI4d
U84sU/hu9vkc3GmLmnCW3JS8xlXL5Fya8x78l1iF0i1PrIZkAhoi6oD6WNVtCc5SZ+M/sEPoyC31
U2+Bf+wP4FXM8zKX+hP7bEFhmRJMtT4uXswf9PKqLxbksWal6iYa8ZM/r0Df4cYFkQjCq/RLaU06
EDrxGC8jHLtD9mgG97ghymI5uJaL19t722pudDnLBhLEMrmUCNmx2xUl03ZFFB0fZivt0xVD4sYw
JWaUS09i8RY8earskS1SIE8U3jFInTWz0F/SB4abSGqwzgiZe5NsjE17o9uw0Ez8du7au8le37UP
VtrBcv3s5lrYlsRncaTFlyn+wmoZXcqr6xZ9lasVFJn+1OvDmfean3Tzw91jR7MSA11OFEp14+6M
Mn3wOWw+E1n3tkHCLJY4iG/LNB2KJmUL+IK/OtOqyfvSZZ2I78sEejsHhb8lmwFcaXU3To4N4x8s
WGEuDP8JFlSBOGLpjCG+XQpEjBIsBUMa91n3JtGIKjKzSSsQOcO/83t4l8RiIP1oUH5r/VkmVG+e
fLsPNLkbqk1xD8zZnOVQnnSJ5b8OW1PvyiQOS/SpWD2JiOCJVdDVmz6NzL009sdR/0eK7oyXtHxc
OoEjN/MBml4FrT5fDqbesQjWfRDmlyi1+W7ZYrWA5R+LlfXzrR0etJ4McM1OAMGRwUj9QWEAOjIJ
SiV/883Jru0hz9Hg2JHzZ65QOyblXWH64z0DilT07wA009yATuGcSrgGqloyIVfAaYjG46PAuPAs
dKICOTfipxaGQW7ervREWpJdWKxcYF0dK4p/XJL3cZVVR1uHhfd74/7C5eruSb14XO0HtpZXOoDz
f8Z6NDAJMAzeMDG/hM68skXpeRgpy3vL9eHUqrbcETCS74f/oUtbWJstcCUHDqHoMeXTxModrS6r
/o49rCY4ciShsEngE3cKLMvAgYhwH9rVa54P3Ob7tvjmjZpsBL4/0W4jDF+58d+ISPSgV82ywPBf
+1wechfbN+Ofo0dNYpiEHLeTuu8IyuAe7VRguEiGeeluCKW0Li4R6t2JHJ7k8enwr5hkpxrbK6Yw
Nrgh7ZllQf/fRxEyLFcV47/yf0h2f8UDoquNGRkQY5GsdvuLY4PkZkA6ATaEmeCyKSHlPzW+kemz
rc2iT/WrqqymgZp6vsAJVWAejWMfk002EgiOcOZuMItu0yi9jSxM6tSqsCzT/mAZ+JimcuEt83Hy
Vm4EruzGDjH2Wpg/JxKwA0BSWEQU3az/3OUnzfgZV3K8hl/2ov/fHGsJNMxIl0Uj+lSZXowwLcWP
K3wXr5zqDBOZAKbNbrSS6vAtSrt1y4BoLLYcbP1IwAGjUkgBQhIcmf4+e0IFBp1d7YgO3r539hj7
dI4KpaieIFsHSKhkqKPGvMAajDEsYSXbBecbijm9dU1sDGXumivbOkJt7fztx9meoSeSZz/7svP/
5lKN/d8peajnMNZPmqmvcdE+HIJaEsDcWUgPCtma/cQlfCyyz5pgmXLoQI/+KiwCezjQR62dzZ8U
tcLKE908nR4z12J5EEakDKPQLlv1uOtpejOEjvQuMcRGOu4+3FQ0v6F9nk33iZSxrsM4du68NXuV
gkZXpxoyJDYS8PHj2PH+fU8c9QPsfu/Kz6OLQRUSMF3T3ZC/d5dvyqlkD+DMI8aSngAIRz62SNFs
Moz3X9BnWxIxnOmvdp41z49zfhBhGDCspqAUElQNG5HzcFMbaNIHeQptrf0cKJ3RvbAKVqd5FT/Z
mXgKA4GepZOA6z+d4o+w4SlCcvWkhPfo1JIYUacU7ZISvZKFJLPxeeLd45QN15rSKwq7xZSH0FLp
nAgUF6YrTqsVtNen9Ucq8HUPeuw+gJM/7uGjSN8EIErMZhJu7j6xNxEgxCADNVknF+isZqEjr1xw
L4KAmNYQ0YCgcg8N8lBTYKHowEM/61tTGB91WJPSBchJ8JLGbmLJM/gFGahlQs8xCzSisAljjxOa
kzvRidwXGWEFp6Yn0NEWrknyXVkGR/DkkGkFzMLSX6nGFc3VLp8RBoTH0C14JiKvXzFai4UDkeNo
PL4DCuPeWw38WQ2DLDRhso1/TkwOj5gZLcGy2EGSir866cVoMz5A7v8XKwP695qg9XS/ZeF9XDkg
j4A7hWtO2mbQl7m8sAERQmCmdCYg8+lFz1XLkpUYbGA/qZWG0am2q47I6rUvjpw0b5NjCLQn2tVz
noqgm/QPSbsLUBW1tM2IVGB0yjPHiUidghGaBJ5QEsLbFp/82wA3HT/8Hpk8XH2rTG8cjo0ImDWj
MzDXh/gnwTLhWfpHnMC/E9nChwi55o2zvF4cNt+RsdlywMyk0XXLGPDDF1omISaL9PAmlyQNP5Hs
3k7HkwvjhScP5HaIG9asauE9W7NZguL04InFMQWyTe4XcjEtyoUFu7Mrhwkf5dBad54xE4U/duDM
zTtc2TyMK7qHYDwOqVJmF1/jTZkP6e4nkbjL38cE0TplgvcEeF3agWF4SKqyK5KtcC5ySG0ljNwQ
sXhV44Htg7cNJ/DacrRLNlv8I+talvCXwOGUlTYSARuSWWwDL28SYq+jH13E/+nHMFrRsvYqZQN+
grsi1KLLCF+WUfZ1MkoPkCkiTfcVZdds0o8KsdidKpClyJ31Ct+KIfipBnByIoKBC1GKomU8JwpQ
Z/SPUBeDD0w4VAvWI7rn+xhycVi8rFBC4iekEjN2UXlBcNbmL7oCK+kxn4QjCa0nDdeHuqx5oB8x
Jrb4EuCTTe3u1wghXczJJXSA0yzgFI7o44Dy53G4F2D2xSwXUHaDIQvPX+CS2IxQWAcrcvuaAe/K
65vx9SfdhcrkrxvpM8IYGgoJ33Lh2yM/ZLHYPNa3vuZakxt/c3KWhr4BYqRgfrxB8Sq3+8aIVVrj
uj05fzw+C+M1BmfPQu9ECD2ENc211JVNSd40PgnVlzDh20A7JakYp6DL7MWNSHaFuPOPBDGd2R6N
PQU8w1ksMEklCCkBTzkKbeQKN+/ASS1uv3k/vUT/n/A8Bx+9hmb8/8bwFYGcNUTJ2lk/el4L7ed6
yphCMGRI2FRaifiLNq4oC/nTP7sMCVBJwzt7guuQbv0UBAFSUM5AhuaBV2d+yqNf6smA6aopbfuM
7tVmBFxQXOeKDn7NM3w9Orw5NhTbALruF+lK8/BDNaSbuNkR7rn7jb9zB6EPN1bNDAdlQXa/tAFc
ije2AF+60EOcVsCAdiPYUHbUZolTJ5ckUX8VDkb1czqJFK7xegNUmglD9VZUwCTI+69u3TtLl6F0
TngcUhJwt2UUIWnCrPGOV40qdOtk+2F5dPk45hERSfStvATe11RqmTTjHMNpx0J23+32sh/ywEAw
yyedmq6qh2sHQ/hSOsPTOm456sNEq7wxrfGR7iacHbxcrgJ/rr7+L6ChHMnkFWUkdefBfZx/L00r
BbNAn3/eZCgD/XwdB7jbIVfn6Yy1JTTH9OGeR0Fyhe11FfxIaLzKsvx0Kl2/d6+CgedzEJLfk0Sh
/FIAA/myzsfTFyUosrmPk3YLtKBFtxImot3NZckWH7AIFxvgIdn5cxRbLj1Az4J9GTZqK0Qkjcsc
6aJhLuzeQ4u7UMkEP3BHMpOTerxe7pFBePJlgHBsn3+ZAUc6har+Ut9G/1I4Olnr4VINdTHifA4n
Sk5Vo/wEKVZyJydSBAOaUckrKufDPlYSgML7EeR5w8705xZ23bF+azUp7KyE2Ry8/8JxB1Qdagc8
f5vIu0DjApyiUWRtOk+xNi5a4g7TMBpIKUKv86/8F+cSeTe8yRe1pu7JTcLZO2ui7euyki4hjBkY
uvoep702UWe8ygbv1+Eh+cJmMvxns+59cAjBYxqhxuz6DMCQ1CcJNAFKOjf3JfLVfxYT7195tlSu
DgzUEWsWY36Fv4x/u4kqhZGvAX4oTezCoLLfyAUjAcmnIL5a8sR7M5vJcdUVNPImYPJqVLMU5u+5
6pkKtMik3nwBN4MsBESPly5U0vo6ozeu1F5Poi544u4YrMnTpXOjMIua4EpaYLNye8rTN1CWxVBz
0htJACM8k74RdRZDzJ/4/J1TAYI32FWkZi/iv0aIm+vgG4XKMPKO1LtfHrI7pKzCy1zGQtsKOYtW
atKx6DPThiPZjsbrTKGiGTEP1bcuA2zi8LM6Y7P8N2buHbR54R5qXJ5bx6LaX/fyPFoB6Zlq81Cd
86oe+E9zsgQ8/RzYw+JqD7qhzHWShEuONznXJ0ctwwroL0Pehwn4qY1+jADGi9pcgdc+LygN6m+b
DHAs3tX3MFLcuoShuEVErSe5FNlbJ/xi8PnvsU+vOthR9Gm9voSf8K2D1VKQNOvIDxN4eeXJwxJ9
znEeu37Qhi/Dy+X+8THw2ZvOEoYkmpig+YqoRR2tmspwmlu7oPQbRI8tcViG5hfsgVCCuaut8Acz
DQPOHw+xPZVlGhg03ISfldp8UIXQEa9WYgMXYCAjTdAwj5bJNzMFdKARL2IQVNBcg8F5rVYDbKAJ
Eo66IeI6mB4NNo1/E8dg2cHI380855txRgSOAhiRsHnNNnyF0yRzdnDLEWesDT7hn7G2S3TQwiih
HT+CHvNijU8uaf80LuD0obvzYMuhhSoy60rey3XEUtk+mAUK/6bF4RRnpBXxQPqeSxoFUJ/HxFbn
kbS4QxLouF2uEvVLQ7Hv6k2oOvFUI2T8KyLasZtu+cQhZtrCA+6bdQyDXx74DbjQ0e4DAVMK4O50
kFzbwDg+1HZav4+9XHgUM1QeY2zsouBGlzkjBbbGWQppn8U4Lh01YnKRTzOGDRxV+o+6O8KDSnhf
Fq7Zx/14jRMmSLEl7bM01Xr3iFvlq6Yu4NLhrdRc8qZlYPcejcdHh9amUVpBax1o9jiFQMxel/rF
iLhbtc7V0HgSpf5zQj2Y5Rs48W9Ek7uc14olngnwNs5IxNKLDU7gomYqcnZF1gmvLwkdgzKTq/bR
uslZISDlYNkP2OFpACMhaIeVjYsmROfJ2PxALjDoWG6YNddFABA2iku5VDFv0AVZBrgTTq+/3dMF
JVz/4YrirFdr7qO5aKfsy6YseinjNoOAb/Use+17qI7v82TlVh0U+/58GU2e7Fm3MJx6nAyF+U5f
s3uuOF0v5bKt83pBqIJsOQcCgby8KCJcj/Ls7O/zKvIjKst0oi4T3btOr/I3mY/4fcpA9Lr8HoZ1
ovGwL48gMWSp3byDL6uYupz87nZzXLuxHdp+lmGS8OMm9j5Yteow7Udj01WxnYxNLUROhMsf5hbq
J5sk79xXT3kGp5JeEi+Ym0ZdcABFlJXLqK38bBsjPvp5dpS+6aspt4gqLf6gzze5/0AK4RyuzHc5
v0R+vpzg4O6cCY9ebvwRfbiTe3gYWNYwNghPTKcEOzi8AmPlBqwhkcLZtxh8ZRHvHnEhttzM7HBn
ugDtQqNf5PZdVH3K0FVm//dufgbgYUVFC7Rd+c6kDd+n+llOOyvlSrg3lIC8vzwjwLMvHOFJL4Iy
3FDs7rmDVRFDUf+7rajnLWqAr7JVabfbAo0VvniqzKW8YRPC1qg8EK25sVnQF0dq/WhOC5DNi9c4
eH5iP1g/C0MG5cB/wdAArErMLKvxgJ2QiP9hBdAp2Cwa0WoWO3AI07JCKYybjco7oAWMLs+/SQl7
cnS+wfdH69JCSsGFmKxhF6zLECF7iEXq9iuNmPG4cY/Z2hThIWtWLjoYAiY3Si9YZ6KXmpEDDCp8
UVDuACtJmjWIyJILT6QakWt0AiPipPCFt12tGh1h+qSfmTMp9MywWlRM6QgN5Jx1t5rGmHjEPKa0
sVWnwhunwlpVxkSRUFHLv/KmHkjETfG1uqQiEGzdUwCxI+Q+0J52dYN+ataCrrueNZe55QHrSVkE
HZLmxlNAgNkN9QkRlQbCw7bjJxdm8qBbxt9vMr7KGFKRDxJdsKEbNRLq11SiAg2oIh9wP2u+wTJs
/lhbwvSuXzklfOLKv6p3S8ArZRc6COiLoFylIJV09KTOw/EHa24oia78DFjFUv07jukTaFJRkthB
QrZ4ik543wzFD6zdbowukuYZEEfY896RUd+eo8510QpsJlN1UVm2I7UECJgzrde5bYZprCxjVuc9
bMpwD3m4wnCII8GzYSN4KsMg1CvZaqLr1LumLyIIgshQimOfGvXi0a8Dc5gBd8I04qE610+n30+E
lw4jEmoWlx+emOTGpRPNItI0DKiKv3yy0E2H3FI8kjA79zqVMbl9V2kJ2G45AGX1aJ0QAwjjDL0W
VhAHjUldWcbjyqW+6k8QjA8coxJGT1vwfHQhsD4PhKbAIy4HAV6x+ynKXe5GycBrjn2T712EJmZR
nOTAEVh3PyGzYnQc1CW0Xi1a837Lzf4Xv0Z8LHXxXBul85XKmLBmbwkQyB+QJApzEwvfN2TZ9Bke
Ld8CAijG98jieHTtGdDjrJ80O8jpzNoRAnkUYCCMMt9WmewprxUGCsMpwPzM06WxHVwGZoL7Nyb+
AIQXbAUiVJiyYNtvjCDgoKhutK4JohioWnSgZW0J/gUh7GpGLQkZHKSyYYiHZvXoK/zQhORgbwSC
2Abw3D4sKn1cEITmEnc6VZHj452ttFEAXZJUoztkwM35XUqcvwfhN2eZBCDPMk4mAnUPYiIt0xpK
yy6+XfGYnyaCTYqzUy460Kg6U0QtSFctWIAlYE2SpFzJ7QE/ZGQ/68PB4inVYxQAhR0UWY4rqTL5
D3ptOf2hgP4xxhlRAbAnVpW2Hi7KYKGw1CRoqn4MpJG5hLRMzL6Vn/i59/QDcyx+CwNodx+J9C1J
QzKxmsVzqjyiqjW7Zwo2ZsFFUIz/sTCYlmPWDWUvN0wEhMPHTeLtTGy2fM0o+OEuSyZl/sutv9tt
YRPQ+BsRWB+bLwnaFam23/KD0Tk9uVjY8Tidd6R5YD5QHT+byrmGyp+9I2/0GSnlMhWsSWRjmlbi
U8JGaj7vMUwCbPDyWxtdF0W/qsN7+Fk5kpp7mWQjyJ1AX1bQjqjE6IUlUW/MFHVK9mX7GT9RzMCT
9I1/1izHa+3NRlxji+7pmFhkZFYPjZOsX77Lfxb37gVbf4TeSvTdcoC4+koBnkSHIvtjo9S5rjYr
iqQkVzGRdmDbGIlPaL0NycCCAqrX/Lzh6BcAtbLv0x4UUHTFM3JnrMKw5t19Pqmn2eRexXD8wcc/
JM8BlNUxPPoLxhQizyhUw7WRPOyzQL3krjGOeqBgDvq+Ogm9hdXmN8COeUKVZieXJMBlpX4XR4Hp
v0sP1jvinL9x0JWX4ti9qOmDDXUm2C0+xY1tI1TQWsPH73QNsMW5BWNkDESlYZ0dVKwLyWcAMRUl
8I/nJdohblxSRG3+nU5OhWtQuWZP+tpbqjm5ciceFShfyIXyvYa5oUGh+hv4oQxmbGNZ12UBSPtY
FpXIy4iYfdQqfEwyx8TYlznZGSmGOeN0cDLNzRdGMu06YnJ7adsk/LdKM/MeQtDNEEn72BUFb4Ix
UT+foRqHyjm2T+Izn9PaSHpARhAX3IFkMvMto2tbxDWED6JRb5UG6qRS4qOFlWgz+oRw097+c6jA
QKFK0t6Ep7acSgczWk3pxRdWlpeuDSLOTCb5tDKjbgb15olL/eUukRX54MkjZ5EjiPFVfQy4xEdy
oM3eCKXFWvC5qU9/V0+An+T1QLB+W8076YlAfxrtPwxu82zOi1u7cxP0Urj0KqnSo/ynYvyM/1RN
SB86oSbY0UQH6LxOC7SHzIMKgIUDrA1B/wSzpDvDQMkFHV21OAtKlrH8S0F6g/IusmqtKlneLfou
gocP34Ws9tP5XXRNkyj+daKTMrQAJkJjl3flC3UV3YrS7VCc88aUWrnu1mtJxbHaIvSVuia3C0/V
Crc3V7tvICfno4Z5xcQjFbO5mrdHtrGF6aPnR8NiEijEzDblUDVchy/aVW4G28J8uR762LL53mit
bJzLEf3j1FzmwYLp9XxIqwv0BdffwCt2uPTivSjN4sDrBPwzUWlkkqd/38v8Vu5XMnajj3JYRH21
2HRnZr38n77eB7kJw9XXm44UqzATgcNLtNK1ikM+AAAXWDWusQsZmqyajSaRMaCCjnlP5cmCJtWG
ijd1xrLGSDj2iNuQDs0ueX1TZnmnakKDMAOhRduVCanv5tz7nOXmcqD+NHLiPDHY7fByU4+0sx1M
Ek6yetQjAJ1m3/WF2Is3N1k3/phqHg4XalBg535aoJMKvPr8tvd8V+7u/Re7ay9+7FyJnGIFy0yG
uWZxwx6iXuyA9QJ5lYr8FigSYINzzVRXUA51YWlxvk8x4rTMN/HknZKW6phYFNL8JzItlwVEf+zq
8IgRiavaQPmmC+/mOhyMk3FA9l0ErLAdgs8H72wCDHMYyTaPhePHDCavSQ+26yG7mnPNmNmkhuNj
aS3DQo2iORsfysvg/rNIGp581HJ5oK4z6HH/25pTVn6Qi3fbXT67xYsDWPRhrIzR7Psk5lk3YoMs
CevuT7y2NAgXjlTA3l9t8uU6FxerSQQxijJ0R0SB4tzDHH3emv72cPi16cZMAHGq8kbTv55ggtqH
qpaKYwsV5MrVivCpn/XhMRiFB3iQxROFcXG52rEjjiZakHs1bvtNpm1k4h3jCkqdkmHDJhmHi7rK
XRljQRsJHSDUHkdQ8nz56ncnqKEshTXB158EcoiFAi1XAaZucrQgMRSUn6Pqz8tXOs9UIlCcLh2+
/AYbFMuY1cMr5WexfSbD4g2SN3lXjeB9XIvDwHd1KEtCNqj9vWT58y3VoVTSRqbGJyLHcWHhW7yM
2WqRTNAep8AXPhlfBdInQYmXj8vD9us4lrXsSOcbQJizGnQJwJhxNque7TUbT5XNuLu32mOMxMrH
609Gn9BCSh8H3ITeb+fgwSsxW10DhD2j8+UvhMMmFNdnwt6DcsJp6o46I9u5NZwbvXLeilz+H4o7
EQ+TwlqmHSx95wPJn5/974pC2pZs4Nsx5mwG3QEeFofkxoeAGmlwwdho6HyZQ3Y31PRvsiGFEi2z
IpkJolZdc9ElDE7KnsUoGHG0ueHWwZNFQml+fPpQq1Y5N9SkAk47fXbjDAFbFn4PW0okOOyD8Erc
hS9AA0V/eD6oafSghX14tdQcKG5+flfx6zWxH8kAmeiPLgujGCSSWN/pMxg/zqbT3Yq/RZLIfjGM
gkiC7X+WQrFtqAGFUGLME9JUoyRKy+aM2eOFBneVfF8joDrdh85AKp8eYkM3Ea5I0LhXgvdjcS0b
tpXAawKns97LbJr1Gv4oChhwk5EV518lfPGj9mIBTfdAtb2ILGuaDTQEEV+X5e0EyA3GtTsGoYJZ
6yGM3iw3d2GYXhUpejbfwcyzqgOt3/Th8kGd/2hwNDfffLOd8Dk+ivqOkk6qDb1s4SBSrWW0J840
2AbYAIDkhfz0qH/Ee7dH/nGuavFnGhAU58lpsww2sKmStutrIN0kQf7NJAJ1iovCab9EBHIQGPcK
TL20dspiRM+JKLMpyiddie5zL1jBhNH/nVr6drDvCK+so6zMnRRvb6dcY1Q3cinGkLj/mbuETBvf
16UfDPwBG7NOH8dE9ZLhWmWgmNerpeslbFDFXAdBaMR4tF4ZCHAZtusxa4qwibTzFTDMw1wDSE/S
ifcSXuUCIuNL0vjQvdzgnIdFc7XhqEi9YHHJ0Z+sKJGkXCxMy+ftZWKdErKrpX9Mc6gXeyky9GJa
PhpcEYqkqUIf6cmcofO2UxrBzWPQ29qLWDuo8PeivHY1/5SucudcNzhxPspYgqBdTavg1feNLhFz
51y3jd8ICNH7BHhw3fFGx6JNaJI+e1LvccUcIjqSiYYAjgTZ1ebVe3ckRk+QukKzjipFe7u3vZYK
wCSGwqO1bR48y02yhXQNs7QR+bJdf/k/3CeXQ4QRLVVZt5WLdyDkiLZhSafhSbSLXaUh5Yo2xnJS
PNxHnlXnVTfHhe/APkDr9cI2mLcP7svLxAGZyGJrML8aewqX8ww35m4U0bWE58qESX5c8mM6TRZV
CtMwGOBP01CLrIv4fQOEycwx3mC/SIa4+70/62ebu0176a396lL6lKWaudNP3E5o1l7KN1z9+Tew
f1a945mrUAEVnkuUsuX3dcgTK9YhWWpfXY3ePLtBJgiqkT8TCaRFFw4NzylnCTlj3ahjrBmsy9GZ
aYXqfTD9vfdlUiF2zMpw7CVN+ESMkCX3UfGHf1M0AB/VsY7lkfliGO3uDj+VNaJoe3+XlcCrdCIr
rlY/glNyLrYayMYt62LN3Q5oepKk6cMjImHenrb+yj26siVLJYWNGOilccx9kzk/+RYqNI82OWfq
TqUltoBxxPLH7tYI3Xtdu0WRhHxXvd5gsHCi/lQG1cg1N9H6MqBWG6eWb6VMiNUgXvNM8LMJxVVo
qshJqvcweqrUU87TuhahNJtEbaCdnWD0umroG1di3+AneFWEAiDgaT7yJhVLeb2OJmQqvHNYulMK
+ao6VVzEr8snhF9TlUTGGOTCRgS6Ao7KjFIX1ndwUlg2iQh2XsOkKd37xe5E5zuAFPpR+TdJJNpe
OqWO9YAb4Ov6gSIar3ADVVWK+F4ttzhGfiVVLNuP/rtBZZRhBuZyS8johJHEpMrf0oegTbe41rk2
igneLWSNzm+EoSZkGEf2aAGzIzWrd47PW5hto19nZYLtwDj7exr7az1F7+r8C/OuUzQH0NI7PKjq
H24MblL0a0aNK9ZzPF4kaJHmgTFQGWzNq9cmCWsQvJ7AHhElcBNuYi5cnOfi/AS4MFa4aFJrQAm5
RJz60CkW7lRtlNEiQUAr+p5LBSGRR9kY4JpKqYGJIksTbDOO0Ht94WYnr3eofzSZKJhg9xChyUcM
KXu4i5y0d33bOMAxm4xb7CPQum1KxAhiqIWmenIDUu1kzB8KcJV1eXh1tIpUqVOI5zGqx7gHuSLr
MydYKddXHoN/eCe3jRvN1tEqgRWKb9ujhwyMfOHn5vw8k4U6Hu0YbA7fdSjyy6up7J452Spo3Efz
ZEFbc90Uxix4DIF6MHWXTNZVvSKVaWST5zsQS7c6SoGNGaQwmeXH85ZysOPLY4Piz5mKKOzzJNbw
0Iu+M9RxkISbHNy2MzcaDxbn3UokKFyA2ApRlPMt90AWcSXyixSBkB9slfkBBItExu/wbS36vQU8
5x/Xa12OpzvAVtZesXynEdHeFbeDZAGCGlJzy/j1zKZmcQFU2QTIlge56Bj1R4HYnqjh9pHE9gJH
1fks4mtle5FKI2VXnmTvE0YG6fZonvsD+inDeWTicgpN6fL0t4OrOahyT3u+1ps9kJs7+BxKRkvW
gctE2lBwQ7ZSI7dvb09UyGa0r1LfEYB08On7R1Ve5HEgJ+P7mg/IuepBflHmao/3fyEog0turfL5
Sg8B8AjvaQWhMS+8sclvuR9LmlMdNcaILMCvINQN3yp+isJN5N9MA/x+v9pDfPWrKSKgiDp8bTSw
/bW/YYZSSs8ZpzNifv7R0QDMmPAalro80aU8DHcZ8Th9oRXjqxTpsRXaqC3+IVjf4EAt8InyNrcC
g+HFrzMVRp0MD6oPUzq/AuniRpoPbSc4UJQMnyNqZEAXXF9FUf2iO0d7uSVX145b3z+FBsFIT5CP
6jvmdTq+RJoKE/Rq+lQlg6lzAuxIl1PhDt2iNvU5RfsIssISMp+54qPkGItTNStay+HNZ33S9KtY
GaawKyL3STtcrEzXyzTuapsaYE+rjVL6smzn5P0qOAB/T3KIZzYNad3xWdaGWCYRIwKr9P68W+lk
5iSXKL9a7WCZzZwj7Y8Z2TWz/xQnmNUuHeX3FYdgMyuzB4GOCY0RisIrL03ktzekp75FsYVfNhPy
tGx0Z3xkfqyOWSrI5MgxEvp+3uDxyCCRvTqDv/dyRJ+Qwb12bgIiRQF+tCecPNP1s58AwkIvilpV
PdJcE2MN5mRroqWx9EiwpRF3ctumnWolHSva+KGzDjWV3Wa1ATx+9nVAf0Wfsv93fJd1aOP7h2Zn
19/MKSIexs4mD/bj683BrXrg1rqxenefuNOfUt1GB0rjNPfBwg0TQSCzi/CZYYAZnbq1J05fENOi
yKTKXYUPL2O31imDPR47e2RxaVxDMrUEi3VXungsq3ft+FxhDTzyLPmH8zjsiJ/1jOCZOwHXu1rG
AEDOXPQMcbuI6ZWWqWV0k4bmUO38IPhocjOjvYuEuc4DlR9rbyFow5lgi3BDQ2en6qqRnxGYzSSG
GiEfE2XimkcjBV5lm7kypp2Tv3zM3B5jxdyKC8rWBwIm1Bp2SprRHfoPqSViAagNkwP+VfkaNVjV
+1WTVcPi+Od+ELUAhuMsqrKqihHQxZCye6HpO+QROLfCC7Qr8hZuU/Ocp8hQ1jnMx7LGvHNVCGDi
sxU5JtUcyWJoGJwNPbiPKr7qigkdeHz25MJgvBq1EMrc2u0oPN7GmuqO3olTmztYIfg/pNspQSpp
kX5zt0Xm4lXyo/+sT8H6356tU0Tp9Sj6tGZz0cUvpDZgetq+IkLzXsjNQB7RN5iVtxN/qxTkFmxs
UUx0kST3Zvp24pDIgCnFV7Y7kbWukCUe8Vvg++oXNqgf4V4DEc3MEPaQ3V9FaY51uCFFQ0JC4fsv
doh9k69sac6djH7a+bFn9rsL/TyB8worpKUeuw1r9VIZANI8C6Mj2zxBTWEIssSzvz1QeQus9nXH
qoW+PiEYir/l0ZeGsrXaq8pVM+qDhERaPtVT1fBKuPLkRh7gfmctS3zwGVQxhJuZCZ9JeUwhVxJz
lMQjccRZ1FbKD95gt01v64+65P6getFkws66ak4wbuY5qZUk0SFj7+YgYmgkbyp8kiPL1bELLWEW
2of9msHB+qcKJ0mK1wJMRJSeugrx/xT0JjY0C9v486DMCDGhcTnUMJWiA8n+Bd5NwMtl+HTjQjGU
zhRJWh+kEbUtCLcH3GYhXWkiwvHEfMw0NUypi0MO3+FY7VGHCJNpTYx4Ogj5DfdkeekL2LRSBs5V
6h0qhQREetxs8oWMf4F/EXTcGxOVt3gC6DOkz60+/h54olW9xdfxI1JA2E8aW9XLmFe9CaGjk3Qx
BThQwPawPx0f48PMk5LCML6pIYxyjgvLcNg2APKvJKY2jcC0TLvLGfUXPnEhar+T8VGqi+9Sog7u
H1Du/PDVL0qUVQnDvtkiEKnHv38oyORX+wgVMm7erxiWU5LRU4ZHfMDG/d+5P2Ib5U0PDoqSv28t
SE1IV8ouweId1M9I3WZNCD0BWtuStDc2svN5sYLJgkA+pMXSJRBwGAC94k+SW1f2Z0Wv4d+3e+W/
1f7DpTSnVrkAHR8rA4ofnT1l8DivprMTJfn/FO79QIW7yMHfeFgbD29hVk31o8j3Oy8rYKdwoXGF
15VQTy1HbHvju1NQ4zVz6MMNtw9SuUQ+cUx0r2MotAlvSnFF0dXVKQOTUZMpbFFF8BrBUGgXVAnO
lQ3ejpYO2BiCHqjQ9jOnp2hgIxoPshGHBlB1/5gH8/Q2GRF51NrcFf+Y716l2qIQtjSf1hGflENB
Rdvu0cDIqC+yavGqajI0TlcXYs0DP9b0rrXhr95IdYyqagX/AA9GiOlJG9hS+iddtNbPlLR1BHUA
wR7bnkpH5tsnXzI1jKLadJtWq1kZi0o1Of8wPTjMRl6JxYIWmmovvNkLhn0ytj6jdF8J0TdSVhsH
oHxtg02zUrg6lk+mehlYqw+umHeTFMGT99OTLj9rqpKi0fHIC6fePtNC4785v7fJtyRQ58m1u87s
qB5cV6KJl01NIpvZ8l1daXU8kLGUSbQVi9mG7Sd9lbbcx1D8G0SD+nkF4OCCdp5cF43zyDkhDkUj
+tfxM2S9BA/diGo/L4yGtysHjkF7USq0rLyCbsz55PKnzyaD21KyKwn5ONLHy3+4bbF2ToC4UDTs
1D0nZlLsaMh/+q3kEH/RRTcdQm59N5ieqoGV+BLd3dG0VbsoIyDY7rG0xMVMnZLK8TQdER52IQH8
MfpCkb5uY9JJ8UB1SGZtmqEiICKijOAwSRGG95SajuPhBAc+4mqG9Uk7ofsMt6O0oSzw+YyYcwVG
WkEf1kK1M2c1EAGrICd17J/lDzx+zRWxK2JHmmrU1XtnQrVGcUGzpL+gjksWEgmlQKJgw3ocn6Ym
qIRqoZaXjklhGtes7ppU8IwuWcHpEYaIICW3lcdsrHiY5xmZ0Ty0RPWzBuX/b2o4qCkmQ0AiksYN
m3c7JtdOaXnHMoTpodvmJfLcJy+l+7VQweVakeA+PJo2+TXlonRAaWEpHFSyfYZcl3mbRc6SAoaj
mzQoImun1UQxoBSE6NgmsTmRn4o0nBMDjcSd+ZXeReGTY5bHfkTmJkrV5i3eDCyXOToqBy//k5Ec
SCTmemCr03BJZHU2bSvUYyw7Cw7Ln391NmhktkIa0PqTBy9bzjGg0UIP3IQRobixwa0jhYH02IB3
F4I/vHMGJUqaOHzq8WjCk5siQE7cu1Hk+c8d5hXuNKx6UQNDGRJ1+8fcGOimMmdBo/idO0LYe660
zz+boPS1KJQmZH1aZVMiC2n2GYdr+s8XSBqtelx4nKyxIht6vcrJUV04xNQQ5OXystKcpAj7vN2M
mpuypyFX1Ev/wf6CmycVvv5njWbFOSj71blAmZI1oCCY0npbxGFl08iIHquqMKeQGjdNBdd/Z9jT
56bZRfw+U8N3O7B/8cwjsc3xgwILhMt3Rm+qee62IrmCyq5loFDWPVuSR5ip8GONcEq6qKIM0MFW
fwVIELQHOLVAATe/t+wueyNKtl6oOiVGH68nl3xiAn/w5r8z8EjFp2wVxGWNeW5LmgfY0v6EXUz3
hwQ2ujOzFefIxKpcXi1pSEx2y7WGMThFMo+NGSka9oKlkCjlUwBC7sEnNhOrYkg9Dwfs/Smr55s5
mN6JGph9ALx7uCW0SBZQ+WaWEInspXJpLL9ON4Sfx/v2yahWOQzWGfay24g59KHmFbXeL+FYDBIR
mrzrr+L2s0hIKUK5fyTq3UUe8Tf1uyzmaRd8/0AApsY2MganyUk62l8LV0WD/prQcAuJjhBq4fJA
XSoB+YoIw55l3erL2uwn9wFzA91qP1pdXupT7xgw8cGrbsaDgYAOrHnj+doo2eDGMohg8k+XLxmT
3CUswf/Qy3rldKfmt+EP70gVLT7auwykJ91g8mul9nvVv62pHRjqS2LC+RAlwdvTLKu6krC0aJlS
I2iq/7wfrug+5sIYYfxpE3dC6XVRcaoLHq1Bt9Zi9yNKOltQH+8u62SSnORwgoryThIoQQROHXcJ
p9hwcA5gTecgqY1SlkoCLDfCYWEJpypdAjAfmDyzNJplHMh67ewqYJQ155D6r91/2iHYEPt/16j1
XFo1+3+bTHQBJvp+tnd/F775hxlxEQDyeu/SkNGWgRJ0j0SBOIsl0llwEXdtCxU8Cp5L7vP4bavy
HDH0urWmXS6Tp+kNrDnwoqxsyoToNY9+nKOST6Wzkc+LQNqa2eXREKnldidk6v237y/GAlk33/6l
Eo96b3zeh4WcRdXLcrmNgb0V4iI8PhOneI4Ulk8kDMCLdW8RsblaV3Kqz1h1ePi4B0wJaa9Fpvsj
4XLgmuZK+EZx90r1aRyHfCOm6yzc9qhTo+i97GSVWRpEZk+B72FIRYlYQsADKoCH9iZod+0+tIuA
3F4GyO4pcBmuUhi0zlPLLl6773WmUzMBFKQlD809gdTVRaGGgdadiOvInDbSTXSukyBWkOg98bWP
MHGl1R3TU5g0Y70PSuSh7mZvllWMGBUZIza090sez2jWEsYyFOY5WgaI58+GZb9FV1hhfbXRzuT1
JXHuvsmrOP/ZPNKmcq4y3FhBlYAAtd06MYehJjOgsEkAwz/CbHrg02riaX+eWydSyJG8cnA1U+ir
BduViT7KoOgDyqCwLAFkGfGFWeOCjb1rHicEQKig/eu83vARCW8fElyTXHdcYBBLe9ov3kiAJTVY
Ego+CkRh1hWhk4ob3+8GNTc3NfFA2FmIEkpyPgFb/gT4eTIRsKjipffG7pEUiaAUu7uDEaMkSeXX
fye28PyQ5sDii6ibyVxfXgJromopylb6n99f0LSwGg01mheRzxBK9MMxeKGvvgm2J8hHp+hgS3pT
o2ylzDaPgzLw1Mh+oROiJ5JZ4dgQtPXSlBkpDzXd9w2CeUMb686Fir08L6SWqxFPcD15ibh1nAHW
sEYyzj5j+hcLvHYFDX/3KzIQkh9DDAh1erxS3p8dEnDvKBRrIRRFncC2o5/tjCTSglShcKCllWS4
pwyDvrduK10bzwJLbZaBNeaFi8HxHk6k9W3u/ywqXoIgP5DsavDsnyTDAC9x7C/aqxpfJ/lsOODw
VziGd5L56O9jGCxOrmsBarVspODX2/vL9gv9FyTyYR6pEc2bfFAjUhAcoV9ysHjFlgeeulO+zYW4
NB0HXIg9UdPnYrnN47b7AHAnLTYhehXB+WBj97kdtfBj8BtidP16x05cqstxhCdaUsmr6pygKOYQ
MbgCCdihQgpsvFu0BlGYPQslKq7reCVMueEFmUrW5iVgD9b5vEhDFZujmCPcG6SK8Gjsu4f755l2
LMZTYJ55CVidR7Qtv5FFyI7LB/zMcErWG3BETagFVaFQLzVK+VY76R1UEsqgJnODzLD2SvETqm6X
7dCF8NpIqq1NmF3nFgPDXqcLp5PC1+Fomg8TTlRr+t69YUk0JcGDVYrN3YFf9kxPPrCT6ndCCw7c
mlVNnZz/dBFxVx2hUzA3HZBHG6h/Nc5//yPdoYQNLu2pdCE3SvfFENn00eiOeBPfcyiv21D3EnU0
6XdDBgEsWzmT2KbqqYvxKdNtXRpovCkpw1FU/A/7t9FGD0yBZcWNqHpZdifVu+1MHaNHrIKJbJSC
cLp50MBTGSbCEmUQKJzz5Gdtdjsc3B43OcV/Qq2EgiMWVm66Ouvcdde5F94zp56kDQQtqCLVO7oZ
xfLwfAWmsNeHODEVqon/h7BELIFobTH6CkSlFaPGoIHkXz/8GgEjfHSrO6nVh78b/Asl43B+AfAL
h0SRT3wNKkp2CwFISmqidSgDR78B8Fy9l9e6Qx7hKMJqCY7LaDJ4kxWjHQxd6+XRyc1Y7leu/ESd
6rt9ZWQcXwMCTfKw8dQL5Ce6ggzqZbzYdN0bg1YdnTH8F2FQZPXOaVFT0l1dUZ/R9OkGRpacXPFv
gfAb+J0mXbX0cBDgwW0SFs14B/grmjDC4AvrogAMK+0asufcJFHkBcsyi0wWFi1IaC+n7dPPyIXW
SB+t9p1HnsboP8kfP1DTkxZUnNi5QfpZt3/qlf4MqxzVf+wH5KCy7S5uLlTub0agWtYvVZWAG7V1
wWPoVhuWsaKoZIJa4yhhOSJ5nABeoE7G5uHZbgAojsP4XTtx40fnRa9VEpw+74omBUOD9NrRHpdC
052qYON0+Pgv4LDdnZNYGxR5N9pJsZyN9cQYf6p7srVZZrSXMZ8Zu1HrznfBcJD5E70wBcjyw9WJ
Ir5AXn+na+MUFpS0ghBz9wHk5SIJ/4ZDuMISTm+nGI/vEpzIm4aDw8/cHNSYRjq5Mo3rVA4v/WLv
yDQZ3czBLFsxdIArL9OA3GaCTv8brDz7P226D2dS7j4u5wPfGIvSqEp4T9pB6AX5ZVvEFxzF9Hfr
iYQmIEeJKhOPGX2vU10oYbRl3eVyXANt/RABlg0JvMdweSubRksKzgq0LSrpQ3k9dMfR00HDBz4H
yy86qGCVxTA5W+OREHbFjazfXvjkUKYaNEFuPyWjdMuzvOW8N7Htgvwcj4gLwVpnr2J1yjdrq6nz
ViWlRrsVJWbQl1b+E7y1ddmr7/IIX66ZmrXcFXGv/TcEOy7go5N9mvZXXqCqDmUPylZOlWOu2oL6
jNc9BqBekXlsIhP2+E+1nnaasXeFAuD7PLfaz2vG2Qjrm2thPOgGQoZQ5mufXxdcvyitO9Nf/+XI
xzGTpYqAMrXdLiiAVEiS+zkk7IAAvSXjSqjqAbaEZBguM898RUjoEHEauVviO4sGudvq+/CEpjtk
zOFSJLVDaJaGpJtPdj0sz/LAspMLzpSuraQhb/GJiI+2frgYp3rl+EwQGJJQP5VfPx9Rx9PmkkGJ
tbflA4LPR8MesJdFmO50fnEXwF/CxykrXVk4MQxOjCb5AefqAig9E0BKHnmJDPFDs5qowSewW8Er
uHKKcvD2VB5FwkA43mhoe38xqfk9nyWOQIDr1HoSp6E4XUDDioegfXSyoUPb6Th38mtffOv6Y5Uy
y9kh+eH9XOtFMStx3aJ51xmBTQVKWURcrz208YlbWmIuvWlBuiBO/qa2aVwdZ063jF4EFJfKYe8X
aekB4rDhy3PoyjVQu15TJ2+baTrtAz8kXvVpOfigd3WaiOYDzp810kP6h75602HEpiVOXIgU6cuC
078yi53Sg72oIBsnJi8hMKOl6UYvTKwgwwlumFv8cc57DxTbQwA+mGxcFoE5VBx2cyalviu4AR3Q
mSiCQq1tvJgPdhoIJCU+NDVm9Olr82Y9bBfjBIuEECpmQEieGPe1kCP2RKBPUsfiur/JfDXkRdvZ
uhGmgTCqLNU+1/e+IxdekKjZfPUaQq2Z0LiH5II6WgaE1j1iYxVsgPPpcVXq0/PTtLSIyaPEKftG
UqbovkbndrTmiB0Cb1oSUyhC7VAOK4l2sa/bXVCdzMLELvAk2y6kHoFosav4ISEwa+Ib5M4dUhqk
5TB91bAriT8NZT5lBq4/c8tS3jMreEgN9WhgtUKolnwlUF1PBM6SUpMJ8cBcE+s8wErxqrJg/Gfp
aN2yOL0dVyAjV25wFwZ6xlGuGhwPkeevb8W4oIqCKalprA3r6v311Rozb8yRU8r3K0/ceDtzDqn2
NqvgBPPT3mZLPl7w8a24jXJfC0mC9DcHtlWUjvNNZlp63+Cg/jg+VryuUgVH0Pti8kAwjXQCxs+o
oPfyXF2uP7pP63jDiO91M5+adqfB3qutE1Catz09YY0MY+bZDsYX17MRwkJylndiLoG9Tptps7YR
k12QcZlbreLSKvfz/fdR2/aYUNk4mJC93lB1mkMs2ObTVbRRlLxPn23xf/dosaAC+k7smilXH9sO
XsZqq6pBSMkexuZloAbS4z5qn4OqD5E8v24UqjwBrxXC7Q+l7grp7jXMNzKhj1EEotS7isUdrQNq
h/0svmcshF2V98BkdrLKY5pwC/xSBMsvHRXOYiC35fRwNWim27dD6r2gkAr1CZcMzuPbGFvVg1kX
yXTqThTr/tzWtFEPiNh1aWNjvPUWiQW2bHR64UjkMBbydmwCX5/an+nwkdRFTExMvvzfCHY1d+nq
YWFNxN9jGyK7GwZ1FUhuX5ZglF9ZXPyXp+MQvbTQ/YEtUzqc6FzlMKUVOgxh+BDG4/jGieDteMmi
aiCzIRazmqVZ31Bnz+PqffpoUanEhuUyhgSJjxeZtPG8kHcqq6Ik7F79uI5syBovKDsTeUrV8uYO
7BxwpcRzy7BPe278HUjSEEt8KKjLA5mydjFB6l7yDt+YzXk7+Um6IBKKCWiRk6BLG15wsO15XT6d
8UMpmhcIqTqgaXJzbofMReSxVV71XR79FWvKCHRIQrEjlIMXZWC6WjbG4YirRBWEgHKoBnzHJv8M
3trQ8/Lfjhf/qWyoK7Wmlsf1xAjU4/EXIPloqQACX//WWNNKGTF102PKaRVq/NUlh5QiH+vH3MPz
JvURjLx9LL3YRre4gy7ihfqekhIiin8Cn4LJTltHYfzlBAixTDJlbC2DcrRFtTdnOqOOoGW21AUg
8J6rNc0cvZZoK+5jcosU7OaPW2xF5iRq40k5zp9AArfewLQQ9gCP1sMr6q6EaZRxDYLEQgXsA3TJ
MG6IZ8InoJ4AGuyfHV3wpdWeAun76fo+08yXuTHO203qil8Up0HkqhXOYlYeba62/kLEKQAgpub8
JFwznTDEX+Qql/mg3p3l4Z2NCI985Nd6GKy7H8as5NuL3OwXjdV5lFzEjHMajTr+9qWIu/RHqOq8
kUB1dLqxmK/32O2K4a6LOUmtPdaZdAURIoisafuC9bo/KafSfBonboROx4cH04spzNziYDIlG8e/
5KPPdcPg1eJIf6xKeqwyMS20Xy3ksFrXrkon3yngNSkcdCeHQKs0X+TrkTZINH1BJ+zZ0l3Uya+A
9xv8toDkj3nDSH0UHDHGmFdNP/Ov6X9D9A/+T3DpCEcbOycrst9PMTksIkIdyOEkK29p5jWeoc7U
fqU335CZVJFDlwsqRChD7ZHI5uRaO5wVkV5Q9beSHNFgwswxp/SEgQmL3rB68k1a2iU5zxZgASnd
ZVvubGkfTw06jcZUUEm2UPyBhFoy/xwUk3FDLOqw9ui96fGAkszmJiwJ/eNjAbjl8OycfQAtJbPo
laBKMcsJKjuSrz8eZUxYPBmdBJujPbOBydgUlpWvguzvJV9xlqlyWZjWa0ulfnyVbkl46wJ9VBEV
l/jmY9SZ64wBKzJc7bqc7ElSYDYDR7uMisSjs270hGsI/WaQI1tLNjoe0gOZmdirnPCLytse8zWf
HC6mTjqg9C3QWfRwJ6UdQtsE2LvNft+Ax8QN5GaXzqKECV1SpPdvFfKtv1u+8Qo23T/yoTLa6z2y
pvxQ9lzfwEqKVzyxQovS2DIFTThxB6Smn3T+HyGusn3Py5plt/f3OCWSKKBLJCTbAE2o55Pv3JKm
Qh00Ex+hmtSiAqXEhiH3YFx223nAOL0C2vTBi0Qi1HcoaxJOrTswPIa295xPYKTJBKHrXpiqoY+m
fC2+HNkTl6AsA3FOHdtVkQ7rQzAt/wJUq+dFoGN9pobcx8S1KON5rlD34NIoDKOeeAtYCRbP017V
8H3Z+ToJyT3UCTRcZen5IYFodTn1WtAjuPNK0OhaARGgm331XYG2sWW5KyvTlEwo2E7XaHoC+NDG
OKnFiokKkrrweYLr2di2IUW8V7D2uMnNtLjRdNQROwT1RqBcJ3DBmDQwGQf1WT435fAkHbIzBRvt
gbdQqDiTQJY4xSS6W5Itwlg5PQFNcj7yJfRF+oXVZabQXnY3TwWr+yHz2Rl0NKFGNfLWSvDachN1
JvF2tjvSYhue9vRWJwbDkuOGtP7323dQTcqqzJUAzD3iMiqXaMLevuZpCaSbq9xUdKRcgR2thPyY
OzgvjtaUIZ9cgEfrz8JlpACtddmlWGEIf0mVcjYmwg9OtFgR4m0cdgVLlkk/Jo5R4u8aoiR5RfUR
ENeVamx85tH9MoB6QlmV/1Ev1v+kQMRr6ff1dfYgC5IxBvYwJm1JBdLbym+Ox5iTkgK/TOkkws7A
cEy0Y1J+ba02N5GWL+0Ynq/Do4AJJeisXwtGiavhjRo+XcO8GqTdN87eG872RnX5kbrVwI11nPPi
nnhYTKAlpRhpmUfYQZ2ZjQqcO0USrgqBPv1VdNY+4Qa6ZVazxsoHCzyi62ythaAQCRhaT0h1CXe/
RmTgJxQ+vybG3qDl1qy0ADcfrdvSuu4BCqLll83ykoy8udKPFdBd5HAaT5vcn3k0wv22vwNtXz6z
WQE/ANXWd4Bo314UD+WDHdJTiZJSdzW54KBHV75lnuEr1fyuIRs5OZ9uQFoNA8jFPBm+yHu3+xt3
zY09Eao+yN6P+45kYm2e59oR5ilk4ABoSDD+2GEq3xpMTgnSlssRaq4cubXpXE1iOBgOdhdZfRDS
fmFI/NG+AJRM1Fo3npcUJgsV/2Hd40RienFxaO/FXH0+0Tv84J/fgMrFUobr7QjTcYz5JssEenBP
KSdVDOLTvQ9yaWZr7pQygVF8i6KtqVXUTu+Bp+Wjn9HZGJBtOOHa45jcXbdGMxFmc3FN8GONK03P
BkhF2p1mHktasZDDkJqoOAdAEcDPsnP87T/LY/HuRVa2aA9wDOb29LE0PE3cGG1es/rs2K4cj2Ca
hTase5K7F2ezux95HzwiFFkiB0W4+Zdnn4RSnAMnrveFamqx9hiZFvsy7f9GNTOpRA1qxnY9yijv
/l3uBWA43lRQm2u21eW3zoN8dM+PK5KO9jcijZJhwIjj3xOB37Nh6QnrgG3JmhsvVwJPaBLZUCzo
WBnpuhCCyxPqMSFrHM78GhQbdeeBGPmjbulDqRMQD/E2dBOxAScEE6UshUO8wNhlJ/ib8zmm8GKD
mNtVzZ7OvXXdctDxw2ax+gK01woFiOW74OHfYJr78CBYXNWcLBVaYAbIBKiQcU1Zy41iJI1KrcgI
xKubiGP+gm51IJq7rHUD6x0KBOlZCPbNUntWCiGiWt9ZJ+kuEwVK3q7qjOR4hkakRuZ0jxiBFK/s
cn954sa+xzYuBgEv8COpx9CYUYBpCuWl+XC7miCn6XpX1SwnbcZmlYTePTAqwshllk5FdSLYRiQb
5vJfgX+W0eBcWFkXHooTitDRDFpGinffCVzGjOCz1z5xv5b2OJZTc60GT/qdisKVS1wl8bzzeUXb
VqkrVk0Mtdljj7yiOwWjlYu4YgKX1NnMk4TgIZASnw3unJhsTp+ZtnwLi/UjG9NFozZBJbi66lWd
4mTxMxb+FNySLGOkaI1bda6o2mCvyvr5kv7g7W/dq7Xz3iHxWcswhMt2AoiJPqXVJStx+WSDAIi5
7jhKjqQlyZc/b2TmyEVXxJkPXL2E8QOEZc+6TkbsSB7B4x5gzHxUr7NYLs0UNr/bPlBZAo+V6jit
py3EtV4n2QYQmed5mYJaCyUQ83n/AYFTixwZAGQGiwL2G5c7SvR1EWJ30szoFCdFZ10Tt1jSf1Rg
XGWrykANzj9bdt5G+zEAhFOtDMXqCyuYGAxl5vaCYowKVjy2ykN3YEd9m/dM8VxbXoy8TeJoAXQY
3KEldhUOqKNLa5MkGp6rrbPEt4W5wH43VR+e047qn1stmTaYW4c/q5ccRkZUleqjrFWbE9+4XeT8
gBAWpUFl1lpDDBrbfDK+u/T0GkN0y24I4n/vg8z3r46CjHrgd4t1MmxGbmIXw4/aXri+RPqQd8uy
STi3L36slTXZlFntPzV/XjeiJeEuGv05hBEF4//JL1WbQ0v10ekJgXHKOk8z1HoROk9DfW8md4OS
K2blPK+82S6QpQ8+0OSkWFTNRQUJt31oNo5yeZshM4oyzkrKNct8tq+nYTj8IAqu7eSe7Uz1IBiQ
gH+CWtZlMN1Ll8RfFfG8wihMCDphKP40ei9QvfzDJZGDI8fetsSBhNhaxfgRkiaEnfCY2snVw7IW
z1WF5KIC0mlICxuBirxnwAO2KX7WZDnTOLSWMdxQLqOlkTw35VgtQPMWW6hjNSMfh+SYfPF71/qU
Oth9FlwHIfaZmaoSKLqkuKIQFxQ8kZ9NiG8EXd4EO6SQUR3dyFealESyQ+rAR9SNfovHCLtQDmuV
IawUlRBgr1WvreYJqkLqhWRWn6ws/WIeIVUU8vJjuFPmZXdHxqDsE0Ov6eEjTLfFqW9+SBEnE63j
P703mDTPtqX4XHWL9XqPrKCRBL9dVPT3idQvuipMvUNJOqmopHU1hMdL4JYW87tGstedkn6du2DD
dif07LQnYfnUm6lQQIN8mHMTjziWSKCj+acg1A/DOpTVEWJK2U9NgYJHDpLCJH8xOtjWnWMKfMdm
yIQaj1Y3QzPpb5ja3iuij4TiQ7DjNuLMohF9Dw+O3cStmE9fxFChRXhLdILXZX/3SiDBUXid5l6i
m6CEa0ZPExdgiiWL+XypIh6AW5OsYw3/B2NZo3vd9v3aJ3AUPuyHxzsA1hvW6REVpWotBV6kJsFq
LosA4+nSKn7g6fHXt3Iutt33WYL4aD1Qxjkdf8M55uvXFYljM/v1JSvX7AdzI2YL/N/8ItZ8DikN
/odzkNhyu9g5pAZN/FNcyMpl6gcdqwfBIGiE9osTxEpzTM0Aj3mEhTfSIqhLmxc4sP8upemgIyee
0wAJqww9I3SiCnaqr4ENC7dn/Gw52VVLFjqZmQr+CrjXMYEokenCbkIKbo9EcNtPDoseyDzSeRz7
faNC04YpJCID+AaQFPM4t7CmuQRXXFvQ0ZR2G6xkmjhG5HcrYFx1McXRdqm6HqLmlsCd7UiyJHMA
fypLcoQkGZf4m5OrTYs4bKaBUk10KWsJLYxwqMVPknm1E/UyIRnS1jviRMIX21xMdV2KunwdfR8v
xwOmWVwBy0ZnTO0q2csE+IVac4V+cFKUhsfGDQyCz52tS3JkNZyUZzIl/RFyKXyDWdHmiwnviC24
vWLUETdgiL4I8v9h+5N0TcEKkbZn9UGVB50yk0zb8+Vf9SXFWBOcCgzITpElzRe4jjguGhHfdpJI
DznD6GL0dY9lxQZ80Gn/PaNQhYMjL6JKA03mwmAqUNJLmJBL7fZF+S3vF9LmcULZxX+RPXY2/erS
4TxM/nTIzdBRigr9hIdaHLesp/WR1IVjjWki+x63jN2qJEjne8lHk6mnDlacbj83Dl3A5ZyQsvNC
ysp6a542LHw03f1ncsY2cQvc2foOIoXf7Ot3fjbDr0v5yOT2K+dPI3WfK1mXtZJYzGx43f8taOo7
XApp4/Rnla7hboAdwTEDFqUupfGbheIMQE44MaLYPHrhwtTOq2Dpo2IBqFitUyHqMEM7OuXLohwW
egLePgeWwFeV5fVhkj3EyeDevKPaWXjoVmSfHALSqMXtwfGewIZCOQj1OIb3kgcIqb4Ql6lk2+wN
+tEjAoAZZjrMJhcNdiD6PmCDGGyqiIspud2pAGkDPrHc8N+nqz6FixajCgy9YcIC5g4jsZc8Eycs
oDFpTSj8XxzlYODhMkr8sIKJUrk+pL1dOJfgT47tFIb1c8EJfzD1CAkN4o/ewb4/yqDD5KfxX+2g
DvXsJtuFaOja7L0jAxKF0iLREpZJGTgW31PeS17x+ktVtCu4og67gsmQWtCZoa+/yQgZ2Ch/XkwO
bnFhi4dL3G+PqN4xcekS+uFKMTG2QTds/LANq7Ac2v5D3iOO3K9PVCTeERa7GLdv7ZICHRf72hNB
xYpmI3Z/Hl8m1u7+LuYbkE8CGtN/SfZsOfi7y8miSJqlj/04iC6GWIc1rrne+IMZOrP+tzm1IGMG
xkjmIN56ekCOjV5GIKNLuVL4pijFomJFQFzm1cA7VcFhvkBdo6BB5i+aktTi57Uv1m+8pBQi2T4+
v+jc62kIfcGG444H4kThl6Wpfaz3VptJf/VZuA7VG3ahdtuHxiP3og2UDa6OT6b83bl9CgRrL1Yb
1m91w8k/u4AAR5HsOsYulhz//gEXEnQSXLnLTp9jQ8BLo3UPWwHE4DV9Lm/LkD8eEvbe2mj4ps6P
rwv/RKY7kAbav6+qkPwqobAl0UnQ8zZey2LEJ4zK9q1eytmSYznTHg4vZHj/zkyqVFHAglmNuFeb
hqGWW3ihL0Ytw9cy7luWprp6gWXeaVwpUGsCXc2pKmAtOvUG9xf+z/u2RLy7OXnN21fCtc/lMB9M
MElYnhOqCQnd3LhfN1YcVNhZzWDpl8Aq9ebW62Jbvg+IaPwgIn4hHooN1opzEnrorNpyy0c+0IxX
cNIOgStQm6wrD2umXlAqllKWBfAOYG0HX5qkVi3RIJF0YsFLncdoJr7aERXNS0JBVYHqv9xtWy9z
oS1KqALbWzkO3rBiZwYOpvQXWtRNqJ5BDwo6cpDwihPUsb2u5RhqdBq7+hzgpAkCfGm2XVwUduFO
tRCY2w5t64KFCtR2Y8agrgyLcTS+ZpMGejPo6i/HXNq0nYnc4FeeA8XmpyuqYXq5+oNb6WP2AZuR
h+Xltov0ePbywG1SwXGjrI9NJZiWvAwJsjXlR7nVV2B/l2ucfbquLF+kbD4RefOtVc3KUjJYLpP7
+iB2ztcWYT9U3MBG29BIgPBSjTcnmw6J/E4S5vkOC9n+J0gE2ecpgQIvT82A4jOpwW0H+0plG84u
YGiPZzEcJJwjSSuQnjE9CNJvQEW+KDQlxYJfqWdBWOaLJZCCTRNtSbT5pbGoniXX5/Ut+Jtnox14
GhQXqoY5HjlHqN7LnzwlRlnJOhf/9tiV3/1pn/J9OeOt1lSJ9LXGOaCtIjR8VX0Zv7/sq40SHmKN
18/AFusJIQ1lEYM6jgq3aBzAkTd0d/uC0SRUtNk2Et/B3QBnsCKydk9+Yje0UNVE774lHzV9mF0a
dCP2U7wSGgkG9bVnBYgvVyDWRh7XOu4xYbc+FSLAXjykGQ5POhYkRlWUgnP6OkaBmLbh0XrmDJ5v
LmIm497T2yYpHp2dxbcFtZoaBx5Hl9ftYi8tZEVtURtLz/G8CXdm7cUgekxGGHtL3iBhUA/8wou4
PM9zdGdKmrDQZnxlJqU5JxLQ4mcyq+8RJdVrl6GKcue6n2obweCpY7oEHJz8ENzRDDVBqew6767y
/p/hN5YwcwZU7ev9pMPIROknfcnGGE6R/DUZuSTR9P6Y1tw8/oh9zaFLkAjF/Zs6i9cFksv62K6Y
R/w3GgT5LhHA/FA/007ug6kqiHdCeK3qaTGOrr8E5wEfdD9uOeaNy/miVr9uaNB6BPSY3Ah3Yt3m
S7PD9DPDXM4Qf+lXKyy7WxPZRwJ1zY8dfP4kWxN97oxkXwPNllHLYrD1YiFsb0Tl6Wl0U8p9zqTP
pirQ+VKJjruvsamoglMIFsq8s0M6ODwvy6vph0cvNjFLJY/LtyMUe/QZdwoBCyUhqtV3pwriHO0S
T85dCndtgThGggUf+kSmXTxsmdPFs/0m+cvdOuE7q89+hiobsei+CLICvdizc+Y1BgJmXoSKV01K
A/0FxlBnq8hLE58bzMa89TLC3CLlF71Thx4XueQboskqANaZQooI57Px4r+pQ57BJGxC40n1L3d3
SxWzWC0hAxx3//yu7nZaFwca5N4CVUJNrYCq3eel+YYak0hJdlDC1aiXgnd3rv3OTTigMheLQOqx
ThqbOBz3PiI4H7Bb037F00S+yEyfckpuJ8dOWI2H7nbC4U7+VN4JpK0EDXPxMbRG/9XB7IY4AF8a
RPIGKfq0CFaVMRxqoz0GqwWqKZkaSlbolM/0o51DTnjHGWTdxAsY6mqDpKKEE5SH29FNBq5DvQ/p
Fq9Nws6+AcsOtBbPCQpIwPQT7J46f14FBkm7aETc32SWJKd2oesdpi7jjpBLZHM0JBESopEmE0xY
FgxyK4Sa7MlbJvyxK3delPkJBSw4VlDstc1zWEg/MIZsNfbXmFJUDQbgpMbzVP5K+Vsw7yZ7cbPO
gDhPrCAXEKsBRTUvwoO2wsWj+sYPrgbiCM8fNaRXxXjCDybzSMx02ASMYO/kqZibgMFY6yluoNUH
y9TV5JP8lx3ocm9PxMrTuTggRnWa795TGPCSJnvfk0pGNgQLcivGdF9qKM53a4ziEfX1ewxqt2fK
6/X+ut0q/wTRnX35hNXexgqMyOjUJTd+JVyJiTrISdnRHeMsjFUzgMAcomZCB9v1qH1M2r7BR+Nl
7/5aLtBtsr+V4q2DQtl6z61lKRqQcFziNnKxPLtwq1G79VjBpvujTthzt8OjLc8Be8Zqktojtc/D
xkipZzEvnlP7hA3SmkFc4BiMuzUi5sUEhN2DpP/0pZip/3VKVd4lsvB5ZBHNztMz2GSI4dfuJoJc
0z+FBeF3w84JU70TjWpWulxopDzuj1TJbFU3d7mDbWoal9osPrVdUvmsSynEaGAHvvaLBe95AOOV
6Q5icOklFC/njnU4TB1p+X3g0qrh00xXdd/Yz5lF1pxgDD+ehBoKovSJ86UjI9uVSLU6UgFyFpC0
nW0KNy4a7QjfvNZCWqzepRFHQZOgAQzlQpeFSHqo1srhx4Oy2iWWEilEUF0dOGvgCgMpV5dagHKZ
7CR0++Asu4ZxklwC9bdGLVoGw+nm3LW2k60rCx95FnqhDF8Lr5/FgavFemoKM9O6JmE2MxaUv/LZ
DG81FdSPtAA+u/Ala6seClgBHO7z1HPeBax9Y5ngJBWVa397OOnR/Zrmxw+kUOflBLZSV8MMPzIC
XsjRXIKf9vUioXqNSxI9Thdn1qyKwKUCAKlexqWXLjH7uL/r1r5tBjMMyn9ftHcapq4QCpCyI9gm
97z3X4/jsVbweWWh5epYxktrjGDKnBzfLFGvq0yOlg2XILSj43+XYwZP9WBEICAKBKqOysRJXsvR
tlKaP5Jx1JyLnCFyPe9RK98Isu5/moPnVfs99NACIcDj7y/z9o9QdFoFAesL8mxIsJMqTJZkAkJZ
k6MtjlPCeRt71UaoTtlE4zijtU/Afey10u7MnkH3kzZUEGYaoHee3OEq4GNu7oiPvYTrjV7YW5Bh
ASY6G6SeUf0JQ2wkbzu+tgCvRQ6cHBJ8vnUBiWyaydt/zpgywJ2yqWB1kLnF4iUD0RW7zZVVJrdS
vK4DcsWm2EyeSV5DWf8HD4Sk8FQ70nzfRlcpmot+yjIF9XFTKOAQc4S3RuvLDrFFE7BTweTImaAt
pC0KqIys3MlSNmG5hoHCbXGW/E0xbiCfwbzisquLRZggxOxuj0/Fl0VAHf4uReZbzLPeRRnxzLdV
SRyjDWkA0eAPOXdGlBcfdx68kqckVrMvE5WD6U0uXcj7KuJWhsOuaBcT7aiV+OGKqMcTB1g2cGqG
CKDGJeNnqmsrLUTCFCuYvYLUyfY228wdhybrFka3oqJeQS6dKDVTHGMfsIy/rEHH6vbXTwnVXNZs
Ka/Mzl/o+Vx3kyN4WUkfAt9YeeauiUgCVjKTOzuZlS5ufM98Zb3Gn8WpVSBx9Fiaige9bMATjlu3
PQpzMCplweByRKu73iCiJ1W4dIbMA2MGGCHNuRRAaPtmgVtGxhAioKunMz6g1Deh9piz61fRVWAH
2jAnKQILT3KEB0dY1RF9ULLAEyWzKKaQ8cjKWSiJrAGnglJJIhi3jT5xYqods1bk71z45xZITwre
AmqrI8t8utrthtc5qSUv2VfdCzl5JvIaeF2zw9H3W2UyD3u49NXr83olBY4b4mOFzgFE9+aqc2SO
qv1CZ2mK9sq1SnfD05Nc8epj/sZv+7VTKqeTbNQtcs9LFVrqsUeuKGzUvps5T/PX4HFgGLmetR2s
NYFEgrYIUFIUrbaqpew0EXTl9qsxJo57MfMGH6NI3YO1Ax4RhLFITTiRwrY/Ai3QOW2BmjQjzwVh
xfFIUpPkPKexpRA02snItXTu1FJgQKjdQ2im7qj1+OZ14JnxUyBmhd4pD8NdonHWC9sf4ZYtd7qA
L41jSQs4e5hlBubXvmIZ6iXH32lG0itq7OubzIhAOWfJBnGRly70nC89NW/fqcsTV4qwOB3M2eSS
Gvo25G05d8bMwTdy7r4PAVP0+YciiccgTIPAd2sNFgNAVOsN68dPaI7rqQVVMveO6wubswhamOOy
QrD6FWZDU6J7hDd+RMgsW61GyBW6WsFsUoppp4VqSFOEQZw4v1lvKOhAcU377QN40lZf6Sh+KRiB
sJNZ+lZzlhvkodanK14h3TJHGcnMfW+DGdElvYAAjh1r4axuNbXSgVOiDMkfXl6eFHOQH0R8GL7V
gxvae1OoF5jdjnFvYI/1I33S3ABNS6ip2u/SX2dgdshtPl0Q06yiQYxcSKU4eSahnTiUOYE65MOC
/LQJk4hTnHmtIMBwKJvo+CMSRWdanpUK8sMqBIkAmmrwuVWL9cPqRVAsn5jHGHZq3oJSAbf5mXbr
eVbZED2pnsDF8QDm41vC0+1ChYxYo+ec41uqWt7Oat4Qd8Kc+RcL9BTaXD7YZzWBSijjR9p4tm3o
SQuxl4tbLOEkhigqlsYa3ORxANQcM9SsOqNmvKzCaUAtOoSpfxCKA8bwaEOBSsu3S7SZByI1sKd/
SNGKSnT9V2M1eflQqJJZqvWp5N46JuZLTwXLWa8ckLn33Pf41SQsOucQVpKDmMZk8Vk3zjdXAPgp
bfhkm1CfpLe68CPmxSbfg2bUJyMKLvVIF8iBlMmfVDn0yDFQaohTiz+xC/BraCQC8POkXmzMD6wv
CJu3ToHJpqojPiUZ0G2T8nA8g4AhfdoHlbwNA8Yn5g6HeEUfR4wecrco2nDDEr3e0B4QxVRqUhA3
6IEHYv09fETRnzG98TjYd9b3nYWAwU+oR1mSbT9dAC6Q4a8RpWMy9P8vt9cs8f/SH3WVh8WJoWg3
dwA85rr15gloipiC5wv02K8b6WdXvbyUJWmYiCdURKJ54W/F21a6yEhH4UIFfQZlRnlchIJBjmdO
pHHDuI2PprZ7e8fAquCOQgz2CPeePWNgrF3NzOGkbgQojU4Vru8CDPKvHvoVOMzeHswDErClX/2G
q1LAYJxYyqypuSPjo+al/OIux7nZ28OE8skHm3GbLm5BYvYi6LIY+hXMjo3rk5ie0vpq95VN1W3I
jLCpqUlCbLAbv0shvDeCO188gv9sf15zpP8SKEemV4iKECdiVO8I6OinCGJgSHnGemkwq5pwG8Nn
uBYip6DkySHc5lhh19IXS0AznzaZZRLrmv7xMljKGllpYz2WXTfpmPSdHFZA+1T7ZFrSrw3HwK/e
3enCU/rVinSP+lW8iUL0WhR0iB3HFbA/ymYLsDSd0vjLzFJSwQDdOmdGGoZE9TUVO002+UBSkqqQ
UfH2w/yyUMWTINlS4LREHofFOuMDBuRG6SGGoeOYJeF9S/0x6Ybpk7xJxB1k3arL1Cy1426gnGpE
+h8iVMvOOfeekUVydZ3Jkci91Yko4oNiGL+D8lQJny+OM7GoxdoXabk8UTnqTAPuz7GC5CROmlTt
Zt+ssKQ3pIDAP6H1NcTsebv5KYiKNa+hJaAt4l/SS8BnnG66+6BipztnHY3oGY8uFBsQZmZyHk1D
Ta79YMn5t3pamw9+2/g2AfskjSfKqfw0Ov1EkYrUL8w/Xf0TH+YHJhiphN6sHh9nARg7hUlWD5fa
ybHJrPjefu1E3KJszYr5MylWLu8F2EmVNwJRenWTaohoP5at6F3Uo2fLeBvhcUDkYQ6b1mG4h4eo
9k2nz5rnMIXOzWyoFrQLiyggiuKdJsBE7f7gMzspLoe3tQCGQEufIsTuSagm9bTIbJDTZHE3KQK2
W6P1rElM8Tya1BBlIrPgCxeMUR8mqOi8RLDTacrxQ5eMx9yHwtoj/S8XEvj7cSIjAOehQPugeSYX
9pNLjev9SyWDW0TZTLxFb6q9GNkBWfie4UNrng4EkjrvwhYUnmPBEiFbE3EEuue+CWhD+u1uGKhz
hrtO/o5+BjcGDRZRRY2EEglfqhIoGXyOE99bqp0Wx2oJhuohvsqJbbyv2j9wU0ygBnl0V8yfC6aI
+p328Qnkl919WlSgsXX1WZCG5uAk0yfNYryYVW+15xkQ98cmEFvJWnHi6c1o1AEG8cr9e85HEOhO
0JDSXyDwCvSHGJjJ9eBEYC0b1BCtuBMXgIEAoGVKSNUWlSWeMonV9UYcj793UZAf4D3sgSPjMZs5
dTHPowcW7H9lRmsHfrQOLmwGlqvqlwmEagPJgxwRy77eNYAhkJ4/9Eq9FQCCH1cWIdzQiXqQrwed
OfoluMkyAY9u0q86SGV2s9rfygOKpNCtv3oNSYdngvJnN8E7567ZhMahzM40oQoHIHJY+RS8HMiz
tw/+lmwtbUbmu5xLwWS/cyKimvZ2F19V62F2NpfGxLofMTML55O7FSFLSzhj5Sl6H8WoK5kmnIZu
J7qsec+Jg/uFz2gO5JgL1AK72Zv5JyhcdJX0ewlGjVaOMVcJkdZ9de6eNKwy5LIdQaHDg0q1BGpG
UTA5pIt3zWRqn5erkApvF/JyYljaB7h7mZeTAckMFGbBo4Dzwysn2WZrWx8MF28HErVhf2Wur+32
nZjWdMJSB0b6iHOAjYtxnSbHi/BuGT0z1YgSezu6mGZ/HtZEPxc/zX5AAPjHVFFZHwZgxnnUp9O5
0+vROVZUtzTZjfPFSfqbVBzndY6BW/70A+t6Z8QTCB+0msHy98EOo7DUWzN6jct1dc5LWxWtGX2Z
BEUXZiVtjKM2SW2lfnDAej6e6GfR2364v5VrJsxWwOsDUTIDSbXFIRZWNpqbsGZtYy1KIgqlutsS
Tc2x69sU5OrFY1WT3wL/rMy7ZTRx1cDLcGgOfUw4zSzrapWEBGlSBhcF77xhXWx4hOGSqEJPj/YL
Tim/ckgr3L3okYtLOJ1l9eHMTkm6+VjyC2udoJXieV7/klsiIsfastLTlAIH/03ERjhHHhp3U7Ec
h8gHp831SOlKMjlT1Zazu332DqwVehF2kPwe9z1oHYDRRaf8XH53kdqLGnfR3gv0W4PMW41NmwEV
FQRyAd5OUUrwSAkXncfxYmkirUGVZG6l1PxW65omfEqCjytdXuaSRrhNcrvYlCcYH/8yoN206skG
zKrBZ3Z62o0WQt1kk9kCLgm4qBZ/7Q5N3NpMEu4zMQMTJTs7gWB7zeM5ZVc6F867VQZypEZ4+MNC
IPU8laKO7csN6IqczIe8rEIJDunNpo98qrO6PSmDOhRvM3KBKtxlxWjaEl4K2lqjDzJNSSD5DPVF
RlRzvuuyoxHBBBVsVAUKFZIsFyJt5K+vjFMkwoE/EydkWvxAiNWSVq4BrJi7k3PUqUgmvjCQQ2AT
9OnhStivu6H7XNecgCCl/vcaLOhuJ6xU4ZPdeevhyAruw3GIBPddwIOoZxemnsY003sIOQKWTKzS
s5btHcMGp8KFzi+BbGEvb2eNOFLW8VePFEMNPV9J1Rjl6EXMQMjtYmaOtM0ajj5sB7bGxCSTK8y2
M353GIZ1vS+vRgMsneSqcJEiJzYxSbUaRzTut5BFS7L7lpO9N+GuhadTl3odIk+irmX6FB6efaF6
t/a28lmp05vjeN3bOxIZTEgG777WEgkUUKLoX6rDETkIUFkOY3kyD+hffxPnKxb292JuiOMrv4Q8
HNxBG+BjkYAeTLUeNxR5YcS/kVSEL29gUrEPA9pFNmuO2RcGCNz7p/KSn86z6nEfMxrJP34FHcAd
4aV3cdzH9veKsvfAv0Oc2THry4A8CmGHYa8SPvBG+7rWExKU2n/yzIj5GK4O6ujsFtThnrnEw3Yw
hWW7QQAS0fNTfNBboKJu40LyWUemMZ/D/s6j8J2jWsBHkoJFOliOdAbLnWwBonCOoJvmkTE1Db9O
GSNN8I2EEUvaMAsvyJNepE+Er5tp3oPEQ6Ly6Nhegp3aqjexTFd1r0546SimjWw+yIOl1wA03J5d
HcCyyM3alESXR+z7fsX2nGByGy02EoqfsmLbYesSYorzp0kgVkzNovd6NkvITlQ0vaKa0iyE0DEa
OXse/CsbPwwXb0w0cOqouu47ZA+zTUkyK7kYSYgw3teYtfUannZI6dlbqjTNXMhk2EkzL3Jj6x9e
uEcRM/oBTHZvV8J9xIN93Hin+dXtdu+ugT2x1qmI/tq/Y+ABebqmF0a3SBlDPit0/+iE22/WDkXi
xfi7sTTmXoRroOn5evSLL+AI0vjwvWMIuRmJLpDSfQmJw+J1A6b4xSTJ0NVDbwNVYm9ka4uYAvPb
yNLXwyol/1/6ZyHykBO/EqdayZNsiojj7RPS9oCygZNofDEAn5pRVbVhnQ05mQrKUyTi4/kJ7XZo
aKQmWOCwR6XFK3a2KYevrSmTBbbCABXMdEjVRfYCjx+i89r33fZt7b+w7njsR5QTgedfbjoPefRt
MwSjIjQ6fZV5dvr1zhrVw86W40TkGUQT4A71gCFY5QJK48SwWIML7Pjg0eDJnBEa/xTIIgDiPAn+
OUPudbUPA8Zwxk+//vWXOml/7SakhPjNPXIc7dpqXluoztaUx8DKEPHnct9P60ki/MI+6nPFR9DV
Gpf9nLhA5w334f6w/89hk5DARl2Gtor1q6asvXjxWrL1TsGBmdT4lm7L1JhZA5eesWEEbbiWJzLR
EyDUlEAu/J+m8KgjqN4/tzDbhgfyKg0+rfuUwXhnvAec5/1Mg/CjVJYrIrUlv3GPQGPlQXAHFYGp
PuJUqVtAoOoJG/ddAdBQBbIhtioDVfL64uf6azaG2csqw2FimfdMQPyxJzAUDDT2t2gtzsLVivK6
6l+gjGeT2LJd3p8AkDPKU7OmjHZcSXX3uVAwH5efWjuh2suCGT/UlkT1fZuydCP3Wi81bWBrQ7j6
a8M7ESgT53b63U2d3dSCPLl1fpK56DCFiYQo46QVzLo0g7FCN/YQ1Y4IM2vskdNjNzvDAlv3jA8F
lptwAkoAwJstD81dTGNiJIWjuF8CkhabapYexLtJ9c684008snQ8jKK2A89eBmi5MTNkhWynD3c6
AGtmni4+zaE5EHpptqUz0enhPZIkh/Wh9Kz78By9HOG2uSqfQfJbo7LOZKw7rNGHa2zPjFAua1HE
u2ejNMecZUkrAbjd4hU4n/q/VCLwgGX72KQJR+FCGcBMY7wcHbLZZKElSWgmTfhvdFVQZSryJyBc
LdEvebrWUTEYMeY9Eu/m9b/W3WkNryCRbWNih3yYsyQWjJNh5NfajP1wjCYMMvv5cH1a3ZOgclxN
zgDNu3nPrVnZLosvmmJxF12blXOEhcBqqIjiH7eg2O+ZdvLG4/UGA91v5fXDU+NHK6D6dwcGUNFg
UW0H2P8HvU1d/G5Ke+W7bko9bKmZpPxFDrSr45tZ3iWs9D4XCnfFgTRepuu7NC7lkC0j6HwDQSba
+1jTPoOCixOb8suQBYZXDAZ0yw38g4XLVlyzjpUy2+pbd3gW2Uoo9hfJk++iD5+srnGlLXINQEVf
Yxww9EVDTTKdrQk7saAlWK85tisDEOM/TQc/ckxBJYAAR9xBlbVT9X4iLI1+bioOYTcqDi9BQ/mr
8QpqNJZBUFgo+AgJTB2UMQxklTH1zP+IgBB4nlDgRMOur3y/QEnfaH5hOc1cq0u0P1MutXeb04BT
GYMoeu3UIyrnfhfd0jantjL59w9lvnKfxYtWGH4PngZQmbQZD8qMK0lGPmYgpuotxQf5kuWBnZNn
wiqZJEsG5SoLEhokC/wtGY5Y4wvjTMRKLPPLI420OyXyodh3wvoSUDdz6GQO05PdJHUrcJkinTUH
irW4yMuy/Yum/KdVYRDAiddKfUYP+bBZQoH/5ka5u/5TPxsL8MvMEXfVm6AZUKAnmU2zo9jECqcx
LYoI0SwpsH5skEdayd/JMhFJFuJqK1VdpS9WpTBkP9R1/c+ebtWCc97rHiP6+0gGaXcU3fvWD1r8
jNJEgQrA+5QBUv9sxJaDaofPOMEb7yR2ON88fOAst59FG6WX04PCjKBokOrUL5jpabj66j2r48S7
9ad00QOCVHcpUhVhLDhVQrK4lP8pKFoOiLdR/n+LqyO6VOOERKjqAEPuL6lz5GzxA1wx77daJDBN
QnNwBjjOLlORQyAmFhOcVkppnf8gQnVEieIQ19/Yy2gtOIjoA+OCtrFPhqklHWPyVxrMItKx4J3v
ETDFMtkuBY5Q9K5xeUHfebr4uOqYjCdKbGOq2N1HK4RKf73fkXA+cPv+ToKkCSpoIE7P/s+tS8E6
YtNybV4OxxGPeo2Uwkv5IhPn3R4zrIyzSkhKuumd8vr5k7ab/cjiKr+LuMBdV/gC3EteNGzx4EI4
Nro9qzPMMHAnnZIuHWXiYo4MLoZMsitgcRo4FpPSBxIueqoSPY3pbKVtEX0nvMCH8PH/4uDSDKcS
/S0pYQev13YRWy+RZUaawBib5B0RXAqbGp04SBgHVngUTsFrmqFO5JnW4r5DAN4/NZfe7ZEQTUyH
dYYto1847yc/mun79viS9z/X4qbOnwhW6ED1xylcPqZWnmU51Xar9tpM/ZpZZPfP/5+cKrA/beeo
FvbF15SbwBUbACv86ItbqU2X2XijxtgJYmeXwrfbua7XDsA6dP0XoXfxmHUO+gJr7vr+vgrbX06g
JqvXIw4DEGM5LulvPZzN+NAKye8FruKttYp+CcrvndfikpGplcOL39pbx4/MDZzddsxFBuYx0NMA
1E/mn3DSrCUQGSthJTgzJ+7fqPbZiE2c3ANz2Cw10Jkb3HViyTztbgJN0ahlJ5GTeoFN+SKl6E47
osVR1eGFQMjw0qGcMx+M2EBXvN1+Zo/sqlOvv68BGBGAnl7q5mz4DEJObzcOSl5k7o/OJNoU0Sel
Dd5NIfBDK6cwYbxbAPFbyx6Bd7ZJbZRKf/LZor2fwk3bepF7NGTPy53dFE/gLyae5JsfmG6aNeg/
phoIT/5Iz02FxrhAn/XOvOwybREKykROgKv/hP/G3IFCfZA14+OhpYfmdL3j6EUaZGIGWWEDakaU
qDPNvpofY8VdHDFuSev44JsDANzFqBY3MpR2ugAMz9zU0IBjBVx05M17mbNd0FAn3fv2T+LJFPqj
sMdvJrdvpr4g+01Y0xCpykcWZaSs8r/a98lNbCDXwJDkhcSwQE9LRs/iuLB4WaYmEW51hWeVq9Rc
IGqaQxZ3kXY5Os5O82JXgDONho41Jf7EFDvyDVsiXtSnEz2rP8fz7aLhi/xYr/HlHRwjDfY6Tq67
f5CEfwJWbQG5Tal0IkwRFytXGQv+1zK/aaHZIywgU9yFcrYlfkx2rTJOM3b0P/jmTaNRV4yR88RR
3Kf5kK3IBZm7hnpB42ZjLnYDyWqPrk4jyfXHssdkY2qvODs54c/T84uyZh0W+gToNGuuEAKOGtf9
ShRN6a8MoV6Xrc3qkNY81qly7RAdGq2D7RO5V6bX5263biGz3GC30nnX7s6mInSfuaKxzOhx8PB8
DneYAoC8pc0Aa7Er3CiIIsaBA4pBq4oNQeMe4/lUIGGmJ4ltY0jvQoaxtbFMbw5o8T36PCZYv88R
cnP+fW0aB3jPKodSPhsmpBrI375IIrh+nRxhiPKf5tvick6bam4Ut1DUbyKL9lBTYfBoeoD7e1Hu
/KSN+jgL0F3T+8j0+h4LjscnfItWGEE9TpuhoEs7e/eOQ01wTacomhrdqGQt1tVuM4LUAO4YrMOX
1BmqR95DD2I4+yT8qu5C7YJm6h+R2m3FGUSFr5I9DTvGrF+RF5VhJITX9w41onwP2/zvnHVINI4G
GzP0hwhO9mpVoDHAdvoJ6DrfbZwBSBpkucNOXQ5xgDS4pyrjXf5N4owezFPZDFoUSlWOQtwbkwzH
ljz1a01Kb6O7k/jV+78Y4b9ycRsv6HgXoj4yFIdsIiSQKKrq+UcC5oYUZKhcb83Bul5Zf5oQTlbj
59uzpzQQ0TaHMP2JIunAZqAZxjBREvg6EYvtuPN+zBen1ycp6Nej4uwQerGkfEWfH1WXRSomlUpM
gdaBu+FNJqfQPrNiD4S0aIUmEK82v7LrUDNc2iS5WAbt8ExQ7iKc59cNPDOvbUs2Wxb9FGGRyIk+
ZXwPMobgclrPlnvfYadT5WegPz2MhIj/HeDtUBXFEPcEtGy8TeuABMiNHx/8Eh1QDzeRLHEvwnAW
pWBUvcuxlKxpo/meKIiKfd0dU2nD9b1wDmSeY3OgdevqjisZhsfrwGSw4Y04BGo7CbTep1IXOFGZ
UWlpcfZbmYJ2s9zztoPKMGHciAgqDib3Ujc79yudwo2wTsISPsGuH04ivU5mA/mr0sOuIhVqbZ1h
2QcT/7+Enu+47vu79zMsUwJpOCDeL176eYDTK2A6gjoi8GHVP6eoM8VM9dkbG55zFvbk9p0coddh
FvR4YHaRcKsf7NlbloZ/TBvGy20y2vnyEgDo9ocTUSkVaClFZydAxRiD/PZl/ExvmV9KlICyh5iS
HvZIyeVD/QaeGTpKtyk5Iaeu6AdND9NCIgbtjSFG3PPewzdqvmLJjS+lG7KXsaz94WeGgWoFJJZP
3/gCN6UL0VH/SlmR9JMvautt6w07q16GCQfFirqwNEwYod3kzoNaPraYLo9R1KAVUdxmwksFK/cX
q5coUY+jrSGFgTguo3YKt+Lm5VgIWV7VbdnLDR+DjVhzRBefoHdzA5kzmiwPj0DKvADTaXpir35/
e1gkqi+oOEuC74JM3uYx+mqbCWKIarNauGNeSaLsyl1O6Dahm2/bkn2FELxc2UmBNrUMmvxKDhgh
Hj2+r68APj8H0ANovseGPB5dnLvVu+fobQnCw3i2xHj4E8WTC5fPZADt7HuFc6SeeHZ4bf2WYonz
YCoUpoaG2U4ak3jlFqfm2ukOwFFlN3BZC0WcS7KafCuRFa7pumlMixLCYmsSpoZ+dvltIQ0IRUpd
ddoNZ+0uzZtno3PuxuhqsyQ2wOTSZCH9hS94UD1Df6VvzrfHQcoaNUX2ZZoO2BV44nNcdE/B4N12
lfwzlZ++Itt01M/WOJ/etPlT6m8gA5HMZENjsio5O/XfWrEKMTY1ybCMbfEZbBgNvJvl5db3dOfM
ydD+goJPWlJ0WNDKCYcjgPYOIo63aLYEnQu0yYeRCOhZMvwMjMlVoYwNFbDAFeAEgUqze6iYO0Z5
fMTrYf07PFqpGmgU7vqG0o41FaWmCd+FCT/XdFEnpu3yRtGC5JAdxUP0WL39k3oBBnbUhgc09gD/
fDSsoSZusrNG5uUMPFVH+tSjdEDbagyinfzJt47SUBlN7oPV2IubVrbPs8ydn4DaXtaNxr11Mluv
oLIMVzi0MuwmMFFQQhCt4IKJMb8zvDCVk5qmu2EoIOJq2ywTZajB4hXR8qqUNXUrFfB6X+k5yXvg
r1K9OmXgtwOjgt5St8VjaCTLI4ReSc/tmAjN920dFjX+pd7+WALWS/wWR21kaDquhWkYHzPgvYZS
UUvyYo2oAAa98P6dfnP+YalPv3jeBDeaBY0DWoswAE8ZbKhe5Fxb8Ement+5GbGzqrEWp4Q7I3kT
kJ+7QtHTocNxf1SdY5ilZt8Rd6lgigpo7LcU5flsLEBDnJAmHeUQM+dGs6SA+qBz81i79eG/YeQy
mWR5f5YHbFZ6h3po6I7pu4bELDjTdar++peEvqsOv4U5Pf2Rg0D7QFdSuaX5qnXkimFuSVy/+y83
Q2QOBrG4/+K/Jsndljfy0x8Vdj1ifr1heKYjytzwDkdu8yrWH8ld99w70zsJ7vgld/D+toRwZMh/
28jM8K0NnQZGlS9s6a59/86jEHKle+ABQVqBchc5CrkJi9tO4sUi3gcldvOMTwCMIYUzPEXEU1pw
r5LlJe3/Xj9iMw0C1lg8v0yuYrzwZ+FuZvGBvLoOUopUPKEoEmh4JuUsYSSYPZqwGj/vOzPtuFPY
7n0WOAMjib2dvFeRBzUE7fehBWclVQL5krwiza8ws241snIMagvaBaGjQ/44QlzC1mIwhyJtlLkx
6rTr3iLJv5ooKtgxJTpC8Zd70gShc18ozhLpSk/aYIAr4ET+WUPuPHo4wMJ9bScegz1URFc5NPSk
giFEi6DocOtbFJIfPT+UPUTkhEBXK+P7jgeSLaot282RUXuUZUtiU7fqQKwBoHRAD0DjkatVWGTZ
JlSvLlBsfpD0FXwjuL3hhPQrNa+VVRdFUbrrLugdsznJOwkiiR5wbsSGDAwZgwV8Ycs/npN1tHY9
L2iVj/trNu7THn43vLz5aXKeXKiH6Kf+G4EmnhbJ1FgnbNU58QWfQ10I6/bDBsy0THGMu8KDos5z
zKbdk7sBOMrLQc8oXEMMK4otMtLbipnJFgt9Mkhu4kOeLjzZQpi2Oq6dfQdMYwEzx+SVWHhVQDw8
03R5T+5MppYX/zgTwE4M8DCbzVoDBNoSYJamcjEjpVvVxA7VM6tMrQnCAVxZK/vDqrJh8UzKTxVS
cAT7Ohl6O0XinxFRd1+p5k/lhn24JFlGuymTFY5pLQmL5SrGjp1rA7bfoZkg7Rn5KVxyrCp1+2W/
jBc2q5EbK3R2CCu0o49+nDTepX9l6N6UdNVRr4QEFqBgaT27GXmQLLOcqnRsq+Z5tNqn8PoB09qO
BjmC3Sk5I8gVfO+y1F/AJcv3u1ZGmed5skyYwiGt3fldemkLsBi1FMon+yivDNwbcot6Q4wpLNz0
gjUEZIUQFTy92ydkMDe2jr75xc+Nce+F8l1CQEXnJH3KJHHb4SECQWc3IyiXLMXpWO0U9YPZubdJ
r01wQ/icyggUmqqU8vHfolyvBWkv7W7uInC/JAsC1+5tPwcfjz1FMDdBMNA8tjS71/ulvbqNyiM2
XwWAsi8pxmpSkbgYEz2woydMIpJ2iKaecDrX15WKmOxNKXxSVSWlifz8jgN+lEVrc+nZe7r6rUur
dfXaRI3dVh5x9CRpcurmyKZscnvSE/D9YiSpY46RWeOC77AcrbW2pTSLFWiNJzHK1liv4dmtWM1F
Z76K4SR1oNhC13LdNK40+bX2xw2NoUfcSwn21VTjGSj9KsU4h3gCANaSkT2f7mMDS0iaPDasL+wb
TPjJpgKJq2gTF+shPWwQPyMmlVDIzUHZibAJcJlO4a6VSXA83YbeJq4ORxTGWqkpWN7dOZjxmJve
iKS3yE+dwhIoIlEQEDA69in42GkP383LTBRoxl07o7rOtC4PE7x4/si6wCYPQKkM0+poakPgr3Pz
u+CtCzcnYpWWmt4E0rRZKEmqmwj8AxwNGyi3GnoS3xKgTnavNZiJtUQSrD8LTycS1IYJjWCuuHJT
/HwSKODnrMPEmgyEZI/dBvjZK2JtG7uWr4P5+Dh9QHka5kItotr9jEWoOS706Ze/m+o/g2UJ4SEZ
Stb4Hsj+QYjErkxyVrm+YhHi9tVIrvHKs8TfJzRclSb6oZCamfXVGte+s5tGGCEfZo9cEMMeZG4v
MREX+q8EV+Qetyk8VUqE3ldVA0qdVXSmAhgWdIMabj2EzWgTZYT00Qk34pP5JGxbxWTeHYZErbX6
LeOk1RR93kzmNMYz0OBLrLp6oxiHVvxf33IemrQqn8BO3VytXCTDj+xtoNe6/L/ZjuEKUnHlZQtS
q0aydkNG869rBOXBk8wfrt6Ndhoi0DL36i1xaVShYhhaLHj72Z7qJnn9xymfu0S4oVzr77NJsJdP
ilX/zzxPw/dfdrKnZLrqcM8/61SEoo6WsOHqMr1q9DsjCE1KRPfdjrNmrreHtaR9RMoyvKIaqT1P
HBB1gm20ncxxHZrrI54eDYLP6cZdMy8Gedtx680Dy0nJvqKHOQLOoX/KHYACxs0jPUtLLFzW7V8G
7y4vFafgzZzn5wAtzi5+Cm4T/SuKkzX4C94wOlTuxiTbmPVZYYFUz7tqtzIyrnLol915XzIilGfl
beucOdDMGrWwC2ZKSyNogcGSXvyw6wFZBGeSjVQchfOoFX+UMbJDlJI1UzzlQ1F2BeVcZuncNXwk
eJ5fr7ZXVCiQlhXoinRmvs2XO7lncyje1NSIx7iJ5IgaGMY8Yp5SlofMX9p4Du2WMY3B89maQD6o
hRipB6gSA1PHnq+bVZ2PLID8ozf2wsWrHhq/04hfqjJvoduIBT5QKWxzO8R/iSaRNc32cjyFAftN
a0CJKZD5t+wD9MutukjbyorSnZa+UTWdoYoU9MRl4YyXHTEJsB0MrhzFXQd5FVWFuNZMZl167EbF
4W2I9L5+x9Q9s1HRxa6ByJ101bc2SggFyA3BJaSSOLL6W/+zIxNYV4IEXXcqefQMk9pXBgqS/kCd
pdK5B0oVHnTV2Atuj5Uu8S16RI58SNEtRhn52H8O8/+xpguEI6Lv8/InJ2HKVMau4+m614cD5rXN
Ux1LYcuUuP0T2w+Z+anTsimPwDQ4k2J+8KiqVbXHrbYu5raVfvpZ4DnvLRAYuy7H3Ie6sxgyp0u3
Y3khQjeRpSDRX34tBCnFPmk5Ga6kt/PcPm1VdGYOtnZ+FuDrWI9kps3cXXUo0ZlhYiFv5xcKPQ+D
hdvv1V9BLZ/j8Qdu9LU/7a/SdsPeVAjJ+JgOwH1o2FcesAFn5lu3BvAlvswXV9QFJvmC/+GewDEb
zC9SPy9qOEfBuLgoYUpG2CEs+G74xMFflZpGSp0+PdQ8efmxB+1QTDUoekicLkXc7E+dIdy3WsuA
mTr6ayelpq5SQqVRtOUqQTwJMcaR73wT/LW9ircunrj1lcSf+dR+yZkiMi5GP2yzYgc7eKbjSeFn
9YP4oBOkkFBLXrqkbbPrSKnmyNdp+9t6P7DMv26kLmD54RrfBMHhOXyA7EI+mDB2pPLrWFRozw3z
beSbMF0SskyS4+fX/sOIz4V5DsW7xHASaCUuQjNSjciVQZkBujr9bGL/s/ixCJViWaxSyCZ+ZjSY
PUdp+K3fAcqxCfWLq6wZlVbrLZkaNdYR6IF2yNywL3TVUTIl/pWJZgth0hLRmKUXt/hfqB7y4KTR
bO9pfIjiZKUbLcrodQRVU5KQMw7L81uSDlp5pwGMJCu1AxIhNknwbKBWNsl+nNCWJBvSIXfk91o1
Szjqf80N9u9V+oOCpNac5CyfQmBncakE9TMyt9QDQ2k6rQhVEMJu/BTo/EnPIvE1ss4h9FEhnCUx
xJByxNmaDpFnVReVUCZUKwdYJFUNUGmILTF7Bt8nIt1fB3+1PlsjziwDLVSKoVIidvhfpg9J2d5o
TkmJ6mC5/gSLEtTwRWa8ytHCbZODQnbrs15Ifd4bQrXIdQANMKgD9KwjIAINWiugZxz+0d0wcaeJ
Zc7XbUVjovS9lRRUpY6tA9APfk66N/+NyUsyn0aDucwPr680wJrKDyHtjpRb+QMgVew0q601ORnJ
qMh59pHY3QsgN4fbePpYDwakvvJIO344bxvK8iMyHyPy935BIV1I3B/QO1Ec279/oiJlY6TkiOC+
YRXEdALrryEPIEGfXe85BwhUnbOwcxJq3uTuHlsEEORX5b0K7zjjjeMWyX300Jc3DDNXl/ythF+s
Q9is3bY8pdXwBX2vlfcPvNkx+lBECAXepq0W6BHqadWe3wh2XPNw5onvdtESP250v5ldzlzzFNCN
SDYF8Kkntkizi1KfD8pqZWuUxC797MoIJ4e1cDnnaKXVW4Fs1E24g5Se0qWMbFKK83Kh/AmQRT1A
u7Dos20QyP4U4Nlu9AjvJ1qt+i7z0Z5Pwy9QCdtFv8EvtcrJ8WtqZRXgNVTABn/3MLNhrmlYJ5j4
ja+OSuPwuLb3lrU5vYwFAPt7wRCRrRMH2qWMWh6C9a9ljH4Ybj4EJo13KIEwFwzCi3XsqKQIs9h6
Hok4cDXTAjPORli0AX/CnfCanclX8TTJBgdmN1KuwL+AWJcBdKyMFWIo7cZRN1DyOF3Ls+uBol6s
1fAVlTkO9PKQeMO1hL9qVLndtwmrxNB9gMjpIa/aVZIOqAds0gbxH8M+5YhYLjr19Bq6j2hUVodU
BcK66wdiP3ce7rjG0aaj/0UgDib5E91mt3okwJQWEImEQiHVD0q3NlPk1EOkZUXeJ1+l8snLmdQQ
efrFbdQpo2h3HITf9O5DbuIYHLP5FTwZ07TiphnfrXAJlfyY4EZHtba7hSsDLyODAgE8pFFEYBI3
yzT9/Eo3U2U0X2YslaEkvvGB8XyoQDAqR7YVw3bG4EEkiJ96apMNuu2VfJKQvcRlPO8XQpbooecM
fJjfD+J6qMhXNM812GjkcLtdNwRfCngkovPvsgHJwPmGFztoOSEQ+vH1gghfJd5LDuA9suf4UHu+
I+FF9Hwpg8uud6irmqWBEZmHM+RklMs20VlPw+FFxt9gRBQp585kZQP99Ii0W9sk3ziWz1ws5mWL
rx47fwOJ/te7LOFKnMVTGQoinE7zW84PoKyvsqdc3sVdwQ6FAOnqJ82Gv0rIVpKa8baV7APIrBR9
qFm3Mbw2QHABLb3EUxcUzhdMt9Eh1xqFrILZaA15kXp+wOIUqwsPjthKU5aEQP9+uyoRy28x4fUj
gXOUiltYJ8my3kfv1tazpULN7ZmEXcCN4z3qJwEHLmjq44RbiWRPcaOngdWhrJ0Xk2+nCoeX207i
2FfSDZDG4wmPtnAPu4a6b+Jp56/xw8alJBBuwkKNqQkxsD4fqYCB4iYgrZO9YJUIrQKkrp1N0cE5
3MyaBssKfG+jCeVr6bnGbVwVGzvFOiBuqt5Yxd21DPbTkj6HTshmuycYAQYduk0qDdSLwge2nQmT
TJ7xCHHZxGqGHvjcY5hVrQA/Ta9TmYReWEvSxjr2q8NEOYZKUWIdnDabtoqCAKa88zr9KA7OpGFr
1VA+uYEkFP+w3NtoXjvhv147yOSVQLNpTxKeVZcRLHzyr2X0HnMQAEFGSHaAliqf3KBNJ1IRMn8G
qADlF9U2K03ZcXteSsUG38sWmOZfs//UMYXYOkG7oDBak+YhNqFE5axrgWNAwNBvaQY38wTbRxIl
oYq7uUaeck/H3rrR2ojVBQo3lrHSkMrPCLIYyUyB5cmiMWo5SC66ZCP279kBp86bDynRTZECMv1t
o1l0QHMyetM2omB04aO26wjD6ywXa7UhJ53SX4ta9YzSD+gJ8ZfoHb3m3LMOxfEBdoDhBuj1F6iR
9NEolRWRGTVe83+BUcmtfkUmwMAPXDuqeeVZf87MS8bqomDY4e5fke7aJ6tmJv1uRFFOPkTqvmsU
w57+xTTQ6PnyDd7w1DXz6Ip3GICEm81Ij/0jFtGaJ9xPMU/ZhELY02gZ4VYIrswD6BMQx7dKbxEy
yZBXSfMosLh91L5niki/gKrGo8dwNtG7w6ZA3P8uNlwZdQUv/+Sm8esE3/eUCmXqzW+W3nulQ6EJ
62UVpmRb2GDBYBdagohegJUHqH4855trcUFyLnftAU5mQ4c3FedRek6hI0ghY4JSS9lCbnGHuVHp
u2A8oVkbS6uBUmaLI4fpnrNmJvhS3TzrKtefM84m4bskkm5ephTnq9qxTRKqwyWydJW9b7ZNBuJ5
LSPeusv0UxzFy76CaRcEZDNZq6j98/WqZWPPDvtVT7AadV3vtucQVTjfTUjzHUN34JzHQstWD885
Zo0ApLc4Hiih4M2+WVDQDdxZyNUZH2xQb1sZRsuZ6p46ExfArGUJldaB6Vd1UIa360Mw4ZnPLi21
6ElJ8chwY0B83uFlQX0XLz6DWiVCKFN0XySn93Ohb5+J6TcG5I7c2itVZNCjr7lFHZsPqL+SxBVw
bJ3H05E6nQ+yGs9w/klU7wQpYJeiDlMFvhZACr3e0hzqRc/C+687uvamr9pqqxVHz/bjJBBtFXu9
v9BrB4iVOwIZR9C7tTH9ecNLkTKOPnMEiLZWoeqY+eoklhQMn60pJLkGCo7euJsNuygiL0ZyDUcg
ejM/YDeO4zTLlANXjea7N9nc/Vq+Jy1Boo6TA3PK+SdA4siEOPaP3Sfw+4v2Cl4tkB9M4QbNM2HD
f/Bro5d3Vt3YI9EsW3L+UFK1f1Lf7rK13kCJx0tApG6LPUVjKdwG3zq/AFK7C+Wk5RsGQ0NjN8yY
yqv95HwWP5umpTcvTyh0Xc4g2bXxhOGs4CClV6dMajXip7MQb61iIuSO8iVUmddUgYwKkuw7DQJa
DaJK+3sc3WaWYoTJCohtkgL9mwel1bWttXkSmu4EE+guL47OwUMz4liNBc4nEPnB9YcIvUgrtund
Fmku13hpjr02X/xMl0F2Rqpd5mAYu7+AZbtjkP37Q7cINBvQxxSe3r+XNZe/C7o5fQVfpUgEi6Bc
XpC+eBAiezD/einKnzIk0+BfaVBehrqijhuVPcwUXY0nvDK2oPXmYg62LOi6diE5B/kQaId8VnhQ
KdsjuZ3nh/NmyuWIIvEFI0zegBhiqHaT0AxOoKIVA9IRg9KBfLHnTnZltjGgxV0eUlOO7l4ufvCC
S9m3D+ivzzCgN/iLs3iwr0EqtjJX0fOXsp+rBwkguV2EsHD5AnDzzJD1Hzdzy9lfKXSXFNd+O9CP
YMvWjofFyxNrSqiRR2Ongg/miucfI2sJBCmSrQva7f9vVqJdwn37rJIZldMEXfAJzBmLxNyBMlhC
TZLFqv7Qjrj9E5MWj3wDKrJbfa46kaykM0qYZRJggMv0ppIQJUFDjw401ijRPST9smIkLE1+Wuuz
r3PQJeJ2Jd9pV+94v1w3vpu8kMMf+XStJeL7r5WfVJlOKs4l4aHgZdBGTNjaY79xhSi7IVdEJsqp
Yvs+5pG17peZXXGZHJ5r3DgB8fAWxIpV0BXPik9I5glXqhoZoYBoTPsEtYh+E4U4bQHGFISlrybO
PxDi4RaBlGaOVHibaywfNxsE8z2AfXqFaC528DzbmOW1+6jj2jrLaYLXHDAjepRUd9Ls7tvcpM0J
OpWY146Ej7uK1503ueVAu1sZDWNp/hBpEb3CKrQ82gFyDYfyozgvHLiWM2sxIoemfPyj6v8VTmJk
Ru6buFHOHX1XU7aPbvV11ma5DH9V2ORlVot9wprEBlRemHCoE52ITTE6ahtcALxvIB2dVKeG42Ia
VgaEC7Q6cgrQg99+U36bMaLZZR9YUgSoey4Z1LTAiEoGG5LVkPPvnBFc1gDgy9cGgLB2GqRkaZp6
AK8v9O5WmNQ2orOQ2+BaVpFZcqX7oWoxfGoUJdCBxaGSHQIc3qw+FZhdF+Gsq6Dilq76a8m6ujyQ
SujiTPtGlpjWK7S2gFpveB9MakCpjIBcQ1cs1c1PCj/d898HQa8o3jwJ9arPTOVzCefR7f1K4OtS
RQScBu0T2oPbCvqV7/3VW64/Lomx312vJkYZibvFH2n+6e/NOAR4j5fRziZFrLBaOHMa/U3WfjuH
pJup76rvdm6Vg16EM7bnq938M4YXIb2pKsF5FhH2wssgTml1kkh+QIvcovhipxeLBecf6SGgjNda
Qj3zsO27o9cKnbyjU4dLJAP0SjpOe6LypG9Ym9c1sMXA72zgbUP4hR4A1+0gInq/v2L56PdZe6z8
YLLH2UiZOoWUHQ0SY5I/WA2iFNLo7h+pTjlefdh5jFImI0gkNxPVOWgvVh9MNusfO0PDlzpeOOp8
DkpEWuT5ClmMsJlZjSPEFhav2eNBGapQDavU/hhZogpbp2HIC+Wv6FEPm0yPviiQM0QNQZP/FaTq
2ZtfkDj1UwBbN3nhVUJl/yWDaYJE0GhUbtKgRFEFB/s7FSdFOHMzFx63b6ZnQ3s3bG0jWa3XOQ+T
GS+/VfZQmKUOuJi/PawNyeYjaQdDtvzctgy3ZYuoatPUHYRF+QHjZVxj6OEV76ILGCYqoO7qz/y8
hu50rbenYDu+SLBJPwVkW5Z7P34yn0Ad2k4xBNzCtqzoTF16gWfOEJza/zsA2T347YXe8q11r+fG
Az70CxSjYNIX1F59dK99F5epkxA+NZ21RB1TK4icQ7BjVWVnveqCWXjUbcXmkWvN7mEtuxdEgrxs
ilPKUw3/IOTi9Z7dr33apEqU2WjMeHCqSUdI8GyL8c4yEtM/8iOiUN1TUdESqQHe9ezfBLcNHANG
v9ogmvR0wQq95suZKry8/RDC9R0WGjMiyF3SmGY0a5fqRt2qSYIfPPDjzc38+qRrY1RDK/H/3HUD
VJFQP+ZBohfDtdH9U7f4l3tzBGk4kg0py+j7RY3bIiTwn66p9nzv415AwD4YxMJVB/1aIXO24Wxy
bW3PKH6DITgZhp9wak4M8HCArnYFQ4nwbMugWhtlgtf+0tkC3QoCTRlfR9U9uhg2lDk3PTb6Uylc
MCyfEHiDFUu/8XEucK+dLBzNtr9MeqOOc0SWngXG6AZ8nMybLeBuDkgczXxNuEMUxoPzqaNMMkMQ
mRp6HulO3JPIo020OMGiXbYMROFBKvYg14Ho5z/fYsfh6yUWRtpDCjrHtGH0yVTQj5KV/lWGj57i
GorjbTJn9q5H1N9q8AYXHOUwRqibCx+l35N6DCzFG9H+HlMU8qsahu5dyFVCQ/65ks/J2Vn2X0RT
zxP+ATI4mNsDDp1afcFx7r7MaR07CVTMBz6cv3IJWH58T3jHvxgGfLh3InWUmnz5sFPF9DdnJeDQ
S45bvI1stO3uXaKaHCaYz9zcJShIg9Fhp4yd56jlinkzlR9IfNzziAe3+i22Lba8gNaVHtbEAN6a
gEAzGN72t9YjagRJRdOf0Y0BGkFsbzYnqEd55YC5YQoRAnH8ofhPqxQX8IAUXBHmNZBYhjF2OvAK
ySv2KoeUOv2iK1lS2AHNsragquhaN+kz306SHcmHvRAP9ElfwamsFnlIVFItUKl70jKF5POfFmEq
JuvU+D3KiZMvH4rXq7uRwnAEQJH9rIkHYWl+o4tqj4FBNdNCN8ha9C1OdcCISw37Nor7m6UwuvDB
h19fW1mxoiMPxFSR62EbIzLvxUtvFkfvZrpSHvWcAXUfHptSQI4kA5ovAgRQ9tfTyBPUAb/yc1f0
z6TxZTIVhN3mElxjwgukQljXXVdaJn9R5WZxzpTWRn66apnEfqfRziP0wIhtRivJtUpRrCvK8i82
iFmuBaca44QG8tWawyeEdJHGYxIZ1SyKVl+vSJuQesZAlcX2EIFA6R47TmYHM2bMKZ84s2j7u/N6
vMXh3qrdvaV4hB1siBzCWKupLtqjsALifETN9BdP6CYDlRlYSX+P6hpJdb6e9oqWH6BfxNUMw5Pq
xnDyc+eQsLxD3TZLvMevLAg6UOK7DYmv9JIrHsZo65tH/0f0/SFQhWjf7VOCn4xBEDjhuCbozXQt
rjpR6Buhpo0Pr5CA7NxGdaJpEVTGdhcdNCaU/b5i837kLd8LQYFGmrJVpJp+48XBTlyqfm6csqsm
NxymbjIkDDP0YSBYVKgcMZwja91YNvqlZwlM1wZbUnWpe4mYGAavS/9riEUlIdBwzV+k7UbhVFm3
3k70Q/szOv9w6TnxR2RIKcON3ZunLstWhNUY4lJvvukdH+6NrA5IWENSuK9qo6J/0LSJA7pqqcRT
9IyeT4CxDKKGllJJJBlOjyilLwO9IRqn3+RYBDvjEnLLSD4/Uo0OZwR4beALjYYFFn2BIfqnX5/9
elS4jdA0iqli59xDHPgZsRszfcU6lS6sV8r4ht7cZTlleu3S057O2afnkJr+WTY/qLvZCQ67pE4Z
0VI+2fWGJhOBKc8ymgzj8DxNb6iokTc2E1anOGKppCASWLWnbwHWWjEAQluGKdn7b9dyHNHAcji/
+FrLGSC8V9W2GnLuDpVnMV9HuqF5yk7+6lKEZSHlVGXIpuNuHOcMnpxi+pU9Jnsw6hKU1N9w1b0s
QlSXGafY/FpjCOwZg5KaF8zX/LUSbFmtGeCjD2+TNWNPisKMYCh4ZZjX5vkRRQ4ThubFBtdydmm/
DYYFHKK/jTCV4HqnNcMlttLyXq22DSuDZ0+txTpKDvue0420jDVwqCnIkRDzOg9CAkmZTfE5tAv7
7kUlYPbSJfPFtX0pCdmGVA/txLmRV8G4sa7a68x3bnwhM+tcSGuWf0Xmx5nya8z/v3LGL/hbJwa+
EsnQvjmVvg1jeb7z92xDnHdAMjvVmyu3sJvNLkB5qgS2nxz/y7O02RSiR42MyHe1GBjUNwYlPJIC
2t8ynLEoO5LVHlV28Lg/TGZF3jFOqTUGSiYmutn0ijP7QXhooMfmUi//ULLHQwuTGT/fVQglPlU4
8TvyQlWBouBUDr0l50pS6WU/m1RoJy/3StCv4ufK5tqfOy4aEtglIHTcP1R7ai79y/D3qzkZa+Es
1MWQjgJQ/5LDQviQU+tQmWLWBqUMeAr1JXfNtCSX7To2y5SdXbOfFitjPh2OL56A7K3PTrwEi08N
+tRyk/eIrx2kVvz5jHkxUFpMGBlgIPADXBMScwRCOAhs9muXDdmYZ4aFLrdYVKCMOFpWwyE91KOp
CrSKoVdK/VxjDGjGKndlYojMJl2Mi8OySUEMCC+DBgv1EQ9cK2ZZIHMIALFmPrAjZy27NrBnjuWc
LLorkHOFQUmuozI6qT7C41F+lbkHKlzxP871agNZSrQxuUvl864Jb/GDL6EFXK6eVa8DDragQ43u
AQqUxMgc4/BGY2ZTJHGBW/WDKjjg45zsLr7vKxc01fjm9pUGSmD025SWGcMfZ97oQWyTshbvPcyO
e0OHD3bjs7xXlq0yd+LQz71pngVZU4A43QuOIuZMTAqHCOgwUl8W6+c2qatTDyjUILZGq1qp9FGO
8AXDIHMF+zjDGlvL4Rq5yJUHwaZg3cQBuAtSs25TyOBh57IP5mzasuaecJKrpoSxSeMH4lpTfSYy
iI99ZqjXqPRW0sLNYMiHWcmIrEicIsAbo2a3Mx5OIzyWngk9H2QuREaCYB7enQg5TUxuXQiLddbZ
Uc+At6vMWSYMAaqRSL65OxJ6buA0vJpno7xv1kIGcWOr8Uplcc78Oqfv8Wlp4LWyd4jg0+yPtW3i
pVmZ9IUyNGdBPmoImw7mjScK5eqJ5+hedK+4m1N7Tg3ZruL9js+uXWiobrBl7lfcJe+vAuCB85AI
oLOMYWILJXh1nx9D2E/ggEtQ3jSB4AfzxDUrkxkRXxsthfWV9MMqlyIpsRgOQth73CVrccoVsVjF
3S74mpi1KRClSZyErv0pguFwFnk6+YxIoQecbOJGuAeEJkZQLKHWjNUw7FMnjv52tZERXurvS4nU
AjAnk/typjd1Un6C34h8IEbATeU2YIHo/6uTfq/gH9LXZrdQx+JjkYqu3h1X16lv7Mz0R2ZJSV5w
MLD90DJ7F+pb8/7FoZ0WSd+Fe8Vu80+HiSR39DUyFTTaP/fH7wXX3pl0CCtYdT5tvFauZnFgxYmw
WoujlylCtsimiB4kRYQlM0v3KP2rpWgX5JYB0wMA28Xhvfk6rzZ2jGTdefYUiKMceAFjYYwwhcnE
mWTqRxIT9SupU4ZvMqn08xuhWnIAhpY15zab0FoXFW0u4FO+N0b+eGxs4TH+/m6pIUuBi4XSBQj5
tObJ/0wdyzwr9nzW07abNVdFR+W7pV/gt9Yw4BfjRtKdlqNnHMfYqB7qhY8sWJQ61KN8IviskpNk
V27POAEElcHiRULRQ7nTyPnOYzDP/P8Y9h1F9DuOQ0z+OoDmfHnglcoFxelVajaiwf83+LI7FPHn
e3+tUloL8+CZSkl2WZ7ozyTopLypG0HT8fvV3PVT0k0Z5Wq28WEmoH1OeRRtIgz2LJL8RUa4wjTN
oRWYy4spVcV3SPmPRJY1ZOYynTff1jalm2m/E+JyJsdic5qVVEGOg+KhSTeTovjE5i2fGnxpUVmN
vDNxGm+yqzYYo8/TTsDnwmF62O66mO1ypN+wl0oORLNYg4moXEXcLHo9mWy8Et4b5YU9vfMyoYcK
VJ7zv/Eu2m5ugTJBcpWO74rwu1Pa9965KD4UUBJrEvlLjMiyNPFMUkmXW41AFB4fYiY63QivKMAf
Mq4qRYV6AlRTML/+YTCY07v8dLsdZxYh/cST2wKcEikVnTYbO4a3P3XZxdxqHEgN96bsPE2/KkNb
PyzdJrvfSsgfAcZJCRBIUHhhEYrqFElB6zZgEeMZArvwCrkrZrDMW3U5rHTUOoV6rJBRHoveFPOF
GHboL7/xC5xklJi6aM1MAtPlry4W4JeoIl0q/CmrEWbRUI1FgCT4xZMGe6cAjf4ObkedqUbs+2pN
oPz2RTuDS4495i6XHhePot5z4NVifyparcc81eyjCZoaQ2xup7p8+IWOr0tA4zlDOknY4vhEh9Y9
AKvUcmQRDBywjch6KKoccrSnwpUDbTlZ9zsnc3m1gVqpdOLKvoPMlM4q0Y495ULDAfRsvRHtQCZK
+ZjU8aSE5xmjH1LeM341OXvhQk+r/9yRnD0ST61A3R+k2Q+mnEbggIFE6BmcYZyy3eygefmEWHQb
bjDqtpIgo0Az/T/wfBIOwjqjTqRV6eJHfLrRGMSP+3/Ct8pDrQULMtI5yEngEXU0NtC+gCO2VFb0
Fe/DLj6HmwGJ8gN5C/Kndx1fMn+Ee9Nw+MVFfdTJtvXzlt7N16dccfcTMe3z3PAZAoaNJbOWeidy
4oCcqVymNend0WQ675DVcH3SPcme9rTXwYwOOg8CDY3Io7ER4+9Ymf1/f+Zj4MhySUUMda3Yj/Uu
tOWZuDTMn4hSlcqy/1drspUpn5Y/hJTAHMsjTpbtdP9Wrr1GGuAX+JVy0sVfHv84GDxFuxZAlT5G
6sKtmwtBRIrv90ti21Nx2qVBxD/E11ms01AF253gB+A+1JzWln5tLXWf2rHb1yzgqTbGo4PVMbfO
EnD3xfPvpnrZA59c+Nzl9majtoC6CTPxGvzNJfuYGuNJZkzQVcpN8jtiOrl+1ZvFGHIrXRDon+I6
SUhYv5MC9hpCHsjGsERsQ51YsQJfbrKWpcFVzsHax4HjhDA85K7srw/4eICLvRJYqscJ32YFTyZh
y6Z56+3hOYT8w/XNUYToIpuv8VBflMhdrC59erpN/JDCdgjk11Mli0DgRkBCrQZyh5HGqaugitQZ
+/5D8u+QSxYiI3z7q0c1KTD/U2cJb0YYW3voqHRfbaGagmvegG4yxOs8ho9DKG3dGUXU//vyAPFd
0wGIBvvHpfVjFZp9XaDmGnoCecxcv7eTzIXEZhSnw7CwHW99sNmFBP53wND5iOeBgdasVSBBuCur
zK6aiStgNTncWWs04ndnhw1aO4el8j1hYYKa4q7x6UZHds9nxitIEg9Kqqm2iDBACereV7+bqrwc
iAFSuR20Wyec5YogN8Fl9wdVg7uYNBeSxJnU3a2eDp/ayC1Hl+fYqUd1V+x3oSShNyS/1vuqUSE7
Jh28fCCmDc8t6GYHDbRerGjI15stXaNUiQ/LYJEKn4BlTTnrMMljUwabzoJqq4utdxzKmuv3DN6N
V9fFdO7qpHLvJPdhU/E7qrVILSfCq8CIjvSkM0PKmtpCIhyBWHAjWayBafMWjKD/iEsQw9EAx6zn
2ymuZVwE2cyQTpEByVWOyfLARRL6oHND13QQplrpy4NUduREtihYaLtA1aOd4y+7CEF6vgDKnLJj
gj/ECssbNmQudFHkQxZuN52Irtcg/9TUquz8WbiZUz+c7CyPlKItBZJ1f+ZdJ4+Z97aCbaUo2Omi
ZhD7GT7Ge9VVvpxBUs7JYkp8OG/fQWTMTvuxuG98bHQnii4MrnoVJBi2VPt+yHdb0mYlAwuYkiKn
DQp8/njjOpngT8f+8eaWT6S7+HpRTUfoiYTTu0c/hAEa99ihgSi0PXuNrJL+Dk7t+FX69eX7024r
wqB55PReYZ7UIADq5+A5/7HmKbhN9yyF2G4UHxLwp6tAJliSs1n/etqoPWAZAO4XEIja3aaR4924
iNfc/HdQeuf/OSf7isuzVFbB9VLmaLlhO+vjbxWO4/jDeX3kQ/2yVl0WgC+CHbtG348UTVirkPe5
qBYSh0OMYh7pfGkuymhVnjQ4hQFVbTN2r7H+ea+oPKiVDazCkXKhLt3jbF21f6AU9WjwZZxJObZY
9jTy8ARAWiLCnLYJTmWyk3350m2g6/lW9wddrC7TDQUPrdL/YImpdvuZkl2zdklkKvv8U+nTUKgM
ev+npt9HjYuHSihnbj3Ow/yIJ+7p4DXDX0BY1NaFmPFxi0nrEDxGaIrcDbXuCcK8vmPL+7uci/3B
CAVoVzFjeZHcGuobKMH9fE67TP3OJVPiPcc+bN+h8o4y9vf0123I5qA/4MW9M5fg7vqDs7VSm+N4
fH7tCpU1OIWUTti/vpedwCusAMschu6s4xbLBz4+6xGJKR1gQ7aRQkNX6xfeCYpn5NaPmBHE3oX4
WmgRTdw5oj/6k4dZ3RfYeX46hBYcB+OA/cXsDWia9GP7lahPnl8kAinAD43Eyq59hHRKt2SBZF+K
R/6OYsT7MMJ8liRaI+jTcUTnRtpGgsx1FtrENHqI2kNw53Ev5K5J6pdi4tcAsFer3xt9wR6APlca
HRSSMQSshZV1aG9v7NPD7l74wdTDuLx+TVOFxQ199U7ZGTHwRVO6+lxfN3WfIF9qqd4BQZYQgk8j
kDrjP7GAgYQmCK+FZkqJvuJMTOjhheXEZiKxzgiwYN3LWqxQM8lRN9NGu48HZqurGiXgmHZiv2eF
nEwR4aosoAEBkrPj0tOperBStu53pNIeptIrd9imWOsrpolBLY1+56qDS1dkssFoAf0WBhhncBF7
xjiHp/VgeGmCAfYB5dyFJStEu+eZB8JLaJoF7aJ0b746jCiP2AqCsH4tmrE5UW8Z/dVqBOMnoBds
MaGj6H0qNJSsPOGG3g3JqTb86NuyR+QKdUNehprbnZa2qW9phDA5H5oA/SCdzY/DRoysYChCc4Qx
XDrJ+8QQc9nHGVpihMKNZ4KlCQRWU1IPlA+8g+NyFxxQQjLUOCxRcvu4qOcVj5XfzA2sesbSecDq
5PoUYfPMDr2YG66TWar5vP9gz/WhauBLAjKfzf4wSW+XgK76EUAVi+FrKIYeKKMeWuyeVcA/WPju
ElLvkCzWFWDsKCxdViFY0zPukvSYcplRCznY9KhgjCxCXxcdTBUF5aJ0od+RMVv5+R5vDTXYrlv/
2WaqapWhOZKEeCa86fs3u4UrR312/joZ/7Goiwy5wluk1XNmtTIDFXXRUXy4eZqd3fiUJH/nHACg
7RFeNbBs89l4tVkuutbBx2oER6mVtRvL64xAWyNzedxk4Q4c7WN+lO7W/Lk4d7Gq3EY2eh3LfghM
/Qu6P03yRYIpZIUT7AFa1gMAL8eHdpclMo7Kef3tmHAE5aN5+1f1pYJTcLW3GYRNBK05oXjzjpNw
WxrC/+oGxXLH6CSUWBnuXI1HkX52I6krQVWpkkm721jp4dAFcFIH9+3Mh7xfLHRYxbjS1OVB0yIo
yY+HK8G/YU8oBWYvHQf6Xanay2wG5bpcL+fl+FebDpZKTaY437KNxaNajGkq/nxsumc5Q/4kh6AO
zJcHOUv7co0awxx30ECms7cVkvCJqXg90R8Sg5E48DhqW11fdCX67BlrHzpvOwe4vI2BZsd2O1sa
iNeSm2ItCBFoTrwrtQ/+HM7+ZUGx1z20Bf47h6V7cExHu1b9j8/ljsEM7BTjh+Nps4EYTGcbMl8v
VbYfSNezyjTOOk/rO/LfDjqxt3mxcxVJpnH87AWHafQkZqtHMxkoFwQi3oZYD+1+Tne8IOLE3UnG
FTNH92wLHLG8n0DZrFdUWP0A2NYmiCFlkOsK7q4s2DsD0aBB89WxmHHbFcYui4JQmR+k0GctjcGW
pFBbis/qUNwWEUIluo2n+LdIbLY/lj0VmJQK3RldDaEuQPISuqQRDHycft4HmuSfK5RB0BebHbUU
Y4dZVC073D8DYd4+cuoUvuDV5jZugDVcJBa7J3+f+jo77NflpAxTuP5gpQNEyVl2RE0s33BnAF+U
4eb2CdOhNruYyVQkE2xHQyLhT3ob54CKxpBM4LQ7cDXAGLxA9Uj01uIgEBCB4H1ceo4Qma/gniiy
HX8D+oJxkj5rUrIfDn2vaMO/W2lbC5a2ooyHVKS/SANx1/7v50ir9fG3xU808539MEqDcJgcQXIZ
e1fY3+xJcrapWfz49dqul/BWISPomimK/kwDyg6w034GapelE6Pog5P3guioTmsDoS8DcFmLdGSt
cqjLAdFaIqhmQNC2ttJLhUikTXjBE49IBD7ulVDuDsX7CHYUzNk8qXmbBc2DlcMD798W3u0sGoUb
ZB300fVr0rdXH9zwtD9eS4NNYJlnHOtSy2fouc+f+XG2W9m/x9WWNEDIZSnA3Qa4VYcfQcE91MQt
ZeF2IrVwRgYdFp/GfzAH2uOMN1/ns/tzs1ZGLMZiaNF59RJlrOD9pgh5C8tsiZlN7YXUzZUwEKF3
j1n5MGF18QvFDdpS0JBM7QbLRmXdBgMnKfBzM0ml7Q5ZQ5Q1RCleAaxKeiqwzPmsEsT6Ah4jBuDK
LNMjFF2WGj2IRzWCicmjfeHzKd2Rkfc8ucLpnzJUAVfkkEcd+6Fsp+fCxyKK/MkgBiV/Rdm+hslo
Ar4YnGGwZatfWXw2uDC/A/FfmRQbjDicHgEVTkEqMjG9FfHKhFq6zsIeKc9PVBrI4BsDrOgLXnzk
q/vg7hq5e6k2r9oVf8ZkPQNsN6uTlbRGHwimj1JkrHE8ktiPhucRYN1wrqZOEG/A7hjO20TOJ0jO
pSRQfYNCnsawSk3cW2yB8xExhw7iBWOznfSJ6Au5Gp4NqvjDq3oG4VULeA7pe4ri+FiEmupP9kmd
+GZG6uO8dzo7rZw3fro3ylSxNy12w/W7a9cDjMGVjQVS49WHVyvXDFMtjv7xuPPwrrlOAdHG9hJF
GK7t1tsveXFJG1hluVGuztIy5LzsVf78HaXzfomZsQ2oIfRKbxCZmxDXPhT7lPAPAcN0nsUnwjXn
FzqAEESZULdLVo69wL+zQXB6QYSTSaXHNygT+FPgfTUevXHH4jh0QIXwD3h7Gn9frtPD3UYygwFB
Kz4IixcMWv9IHlBqo2o+SnZomh3UctxVZE4KZWkfrRM5L8mtJPdFX8Dp+wn6S25oCyeRoiZqpFto
y7CBgS1SMn9aaeHPTEMThQPjP5qCfNcbT5gVi5EPRvvdY9YgmUJMFLOUSwl2aNt1y1GLv/FlYA0q
KJU8Jc7Ceae5wYYm6Cuq6ZVxXRdYbs0/etpLL94+1isAhNl+ATihDFnUM6gPhWIPfuj79lxIon4z
a+0z0cdyNTdgRK6xV2V0/seY8neAICI7GdjKkHJe0LXXH8nbcXYFaJX0YDiYdcR/BOVbSPdAnD8H
dVAveGn/4XyCPSh/NahLPs2NR6dQfBMBF/QdkjrNQ2UXZNV/IS+AlfcjiKktyjAnus3DvUVOLDze
esjN5BGQw2hRJCm33vzQbgVaW0DC9blVekJs2mqk6SuibnJQpJt9rjznkcEqqytlgdmVQCmCMW1H
gqj6u+QsAb0cyBl6INVCp9GobonYIju4n56rHGOGkBGQCWWjJGRyPnVNy73CHDiUU/5V2GcTnSio
esk9hH8AMTfRxNP32fCTs7EidIqposQlx05vrdoGQNnd8rxlXyRbcmytG9S93Q+Qo7AGnhjoxsU1
KXUfNBP+wWC792kvMV7azks8BA89HhhFowZ6HUpUXajiqLzkiJzRIF8e3tiWNl1iwJJQXy52cmDu
pUgbSM5YDfuvUe0RHf/9xhiWwcE+n3NIHccLJzJgroVBe0Eu8cmHCIC7VozEpKBPKA03ej8nHtY3
x8VTnXuuBzA1E0ECV9izXjccpi2EPFQ35QHVw9dVo9sH4A44Gw00Asfx37TFUNir6RZq8I5PUdmA
br8SMQtF5o8BzMo5fkwGxXLWynBl8ObcwrJoXP5B6fNlKTQgz/Ge6Ww7QqmCf7uH5dN4arkBcDtL
wwuqoO8rXkizRMUZ89Z8Zssn45wR5FPHUFblUF5PPwdSvjjnFXVjIfCZtASZCSdt91lq90dJoECz
BXLNF2QGRHgx5R37z4zzjjRB/dLbSHWwt7UuDvGnvRGKvzAaJg+n8Hi6ED4Pbi1YqQiIMusIwp7T
R+N4LqvbLLB/vBvXHCcQfX8nmOSg8z1xWnYO/sN5zIAVBkX5r6dUbRqmMILbElnaGIsXNgL1J+1L
X7Hs3gGPRhcQTh8gTriWhQzoVkwFzrs2AWK+gy6cXKUHZqgVTPoS5xAdfTw7Fj2hbuA7FZnp/SmA
cS92MZm81G8LTyfU2f+3TnhIIZnzltbbCguLqGQNtCmEo8IEUeJBomzczsQtENdHDCLm3tiqInc5
qqUSAerjrV+wssAk4672/NT1rDNMny2aQh/GDmXSg+/jABNeUtNcwNLqNLB8sS3b0wqY1Cvo87KG
TjDsLtWa/W/AE7Bsnc2jlUSLkO5PnfA+06DU6MU3mrRc3lUrsIWQmdxZ6kL4ECWe/1l3Warnd9XH
0TvakMtsxm5mBi/O25CpksD96lhsWY/CLMz0WixVMQQrnG94d0YtQ+YHKXaFf5e7+CstdixQSMV1
ABAe3757j21o+Ppqh/Xaca1ZlFDdw5Z2v4CMAMeWPdl73Rd4iVY3AsGzOTifSkKZlel5sgRxSNZO
00ZJHEsbtVUhRoE3ohLcuZvLvKRA5X7N1kOLNtFefLpJyyMffqSo8ukiE3QnhIVgOq9ifMEd+Qe1
PkeDh3rorz23xGPqSRhb9nBCXsuuPRZnX+/F9aTqQwz8nJ5wNmIQRZCfgJmUX3wGxT1RzXMpiGZ/
HTOocyhnuQN4f5csxw4erJVN1BphVaMpvsISfSBhrGYKkrwVbgFulcN1ya2yRBQQtmlKVKbYuwTj
bemPLj0xMpESTehMRPZVgbcYukyly8zJZaj4E+1le9uSm/5a3AnaUtsnIFReBYlywnbnxO+hfmht
OJCm+DQ+b0KRPwMkbAWrZfCJ+Tw4XkNsUQHqJAOItlorB+P9S/owpzqa/MfxgIhkomlfRWBtqSYE
DyJb0RJY7mH+WAU9YWGDlwX9jTg2w7i2I0UxT9qFt/FVIbqSrYrxQPz7Wzj+E93Bc479U+fldaC+
AN7ngT6B3dIS7zoBiuPX115B1SlB1XlsRPpmYeMlTGKKfttV4uWSfHzdxJujpx5PEtbEY9UxeaR0
IjY5JvKpMnRzh2DQjFEIPm4kJDxblXG3C19Rhwy7iiDXwBvRR+aLCdoTHNd2S4+QHWKDF9pHDCH/
c3N1/Ge9cvg7K46at97U732aftZPO83jv1fwFC+BbH5ox9JDhlrbvbskg11wfp79+QOly6/WIeUQ
ZU7Dlg4j9rwbOgF9Je/LDbQvVGqMYfMyKxpFxvDfdlaXPcKYnOgRrPxLIsqYnpE5e/Hrrnu/g+b2
GnopgMY/O6Tkq8OBasRcWp4pTBM9u+ox+2fY1s+XvFceb04z4sei6zmv8yecBh9QMMCG6hwFu6+p
2Z+q8BqIycUmdFsmqb0nBupHReRfmYf1XJxdUEe9ml1hUomEFu1ykZ0jRy2b/xFooGPrHlps+cQK
7uKVCrWpAXLS+J856e4LCLQ2KILO8JodsTizXSV2mH3Vo3JC62PLg8CEv7AgK49MCh5ajkAUaplj
UN40YHPIFzV323WYg1y5qK1vmSZkeKXhxlGWgTrxqz+ZFdAeIbXoZBuni0gU0e3HfgSska07frLQ
aHp7yJPZw3qxg4zIIPl416LELAV5/cyXT63zklu9eriamyiG+ymt8TanAGPcv6IepfiI3o69O0yh
8mAVGPayiyBqtVlyHDo0eXMcgeomedndaq/h9jwz9Uv+azutH9f769fnEfUBDCuPbAHGUjU/HXft
GGXY0UbDPVhnjuY4vcIZHljDgovZWBpwIJQ5LQyA0F7V2m/7iYNZNBtbkuisqnuOpLFHiIeVlEgu
uq83rC5RN2TTUqJNNID9MVkAvKE3YST4xn5B6fu4IsW7IMJEKXMEWS6vgBt0Z39HJiY0mOxq5FZE
kxWDANmdRzsO2plrZnaSpNK2hvGkF8Aqz+YKOFqePCJ/Y1E9xfoUlgFFCGkvwQv9tOaflbWZJzPN
N5isMOcFV4Xd5VC8li3I/4FmaXHJ3MWqir8jeCvAxpXKwphgJ/CcsJHkOyqbyvxHSwJO8QUd2xbQ
BuLVc2zK9RkDQVoE6egspvr73UsjPmxYsXHOjh9dcyKX9XywHJxd0f8iLWJ+TPktL/177wRawMIR
roIh6WDmUdHcstu9MueaOqPhr4PsQ7t5EAUX7BqS3rVRh/A58jHQOI2drLJb/mD3pUCCcuGxJtwV
lpUO6IWVhZAwau9bf3knfsD9dSy2Zbnot1c1jbOxWTfkgiW8Lu4JA9IKAh1oB2jprjMgpE79UnqJ
aK+IMP7w2WBDbeb9/yRrd+CKrDNBV3f3pK0EtZhgHA4uTqMk9uvp01CzO7IfugADcsvb4C/I5Jnv
N7iKOID1pb/fXEome2XCwQ7jeLqQTuks5AXARl/9BKiQONeLrLaI9kPpjBSplZKJTVftlkccKwhA
0ms9BB8voWE5Jml8WVNA3KFC/y7id379KWYl0IbDwo3lRM/mtDg0Tg3Fo2DhKcFD/47mbmWU3Ugj
FAAgnbJ1WpwaY439OBJLN5nnw2x7aKKw5D6amUl8IFWb8cjqF+rXkPVubGKLWQBStt2n+2AMUWKT
TnUhd+ORn7RhbENcD/gNvot6ZOCfX3J3x7IocGPJ2gHRz9Lg70ZlKkNEJ+ufFgIDR32JSg6Y2+EL
NWo9W1QwV4VpboY1ZgDWGPnz0mrPuJrXcpe3ii4Yg8rzWg/xCXFMq0ikjzeH+Hg4dVAx1tErpeG6
LJWs0eyDhpQuXTsNshWP7BUHmu7zFo37NEt/anSOMr8ymJ98KZTIHHH49AcbT4LHQm/C9HKQ34UJ
mDqVWiEznMHzWfnW6F169Dv6KgMB9vfrGFqvxVMIT/87puabQYrwC1PLo1ELGAKtPLN5brT3tjz8
A4/k34NSOfEQF3vNU2EybEtmPkimH3W8BojHFv77x9lTSy7stYmOSa6E7gwlhRv2juoHAe3rhcnW
Zro1FZDQbwi97v0iJsfcVVdis9Eycel1d6bIhXOYnNgi0Cpu/rh6NCVxJBXU/7d/nZlv5cMSxufw
/Sh2rQ2EY0mg30ihw6/20FUR+2BkVZvUgcyZehu+fC4E2Wt0BHNM/X5dJLd3+lWJmXl2kC1Ul15j
vRDseZAp7UTtQqWFW7XBe0GjNZTrAHPBEfSrObwhElfvZ6f9NAUxCSO+N5z2DQWjymHwLOZtFyhp
VX9chORy4n1z86rxKFf1fKqyDUPXs+4F1h0p+A3PzyPo+87tdZnNt3yCPPLWP5Uexpvw/5Zof6Ij
Tzznav8cs7WGgVX/HcRjmbSjHRpmevEJ1vgIL5KZPhQrT10SspNerfXHq0yZS0GCH8TBmUn7aL+P
qhGJ0JFOTVzAJ11GmJmRB37pcyYj7EF3QR7FnS/67wXT5ZisqwOncaF5zuf6mOD307hkbQQmmMg4
PBk0Y/06YHj3Jo13cvmA9u6NWcfT89LaWCAvcGXtiCYdnKoXtwhY4xGQf09nu6h2r7nOhEOqr9oJ
x4zmz1mKy4uOR84NxlGT3RR53UH8xggErmoevbFK+1LBMFePpzXhbg6Q36YBL4KuvU2zZRhEjLJC
7IbboOQ4wxOj+U3kJ37Vz18GRpnJZc16SrcfrPGPGV7JJjLzDqwKORMbCu0MF3/s9Ud49wnCX4cp
OXqFkRynB6bMHvGIYrTZUN2KG+qtsExaXlMdFQCq2d06wYaOCq4KjEz8r+5FFtfG1/gzu81+PZKn
KO6Y9TioNdyby/W5+m1kbBU3NMssF5odXPEfN1QYWtqRv1JsMmCo9Sf8Q6c7p8DE67hnvaA2Hhae
KkNg+jkO/MhrrqJ6xcL3ZD8WQrWGQNbbajIcZT5IhqUejPGYtw9mVTgv4fPKWOTwNQuxbcEAImh6
BbQgAuTx4fUPgFkaAhiviJUy8mQrtg/Mp+UH7YArOGiIDz4iArVSqItqxTudWFwZiddzMnIf0e/O
FG1z4xeqdgIuZRc17PgezuyEHOv3b9RFR//CtFwDOJMUKxHGWoacUZ81hJc+AJmeilB06D7Yr1YM
L0OJkfsMtLRqldGuN7bGqwJqka8HdR8GbaW4dZFpesJ64N4uZJ0AQK1l/T+m6zs4IHcUFMNpdvJY
0p0UkdzEkt4J3EeB9xnV7G3JtHlj9bNWO4XKBy2zidlCcEKYp5nZqh61ZgS7KiPQIki6PnH88447
G9IIoeF+TFV3IUbZvIa8/aI62FqYq+COr27x0CzCDAi6gmKpo2YP+fpXBYmEGuSSnyKStFN+e/P9
tGJUE+ENMljLauMsjo3SddjhpJUOEwXEZ1tofqbCHcTkLjGDJe2pFWqCjwguf0+Q9eY798vy9znU
3TbIkbfHMdAV5ZG8ToYACCU0d93k+GuzMpynCOfTzn4jSS6ao8/cD7xuhaO50uz98q3a1dnWtb12
kZl/yJajeshhwrAvpTwJzk45Vhc1NVDZH2DGYsY/6cOv2S+UoYemRn3FJW22YORIrB4DJnPKcthm
61TNo5d9S1QAWu5Ri267qrmAPPV6NR6MQT8ifUeI9kek6W6Uaj4V8xHQC0t6W0cQpKvmqhRatscE
ww71Fs80tL+i+hN7JVq7PEPJL9ZYtmfhd+L3Wa6+r/uOMfoUv4BWDyxmOm9HY95trU1EOswYTiBv
RLSr3ZL4EJJ39f85hqlLReoO+V51a8o0w5ZuIYfoOQw2AQimng3uswSYBBXq/mu3OPEpZ2x4W8wM
2QCp7OwM+oO79oMy0uI+PVJYFVUGRFgrcCcLL22mrZYC7aefW57nXxpc/udzbyQLWoXA+RjIlN28
oGXBuYlcVnjfwCJGkeRD2nf9m44yunNhCWeJGXHTxwdQue9lrMFJkb0sP3vSpV31gy1l9Ahr+0ie
EpCa/qOfzGK5mmzvgae7aUrccg5eth5ADtU4BWd1srkP9KrsDNX6aX+4CjEB/BHgODL28dUzconY
AM+6EfRKTEkXO2r6mUQN3G8Sf3+oDPT5KwlV05Of9ZKWfcQSZOR9bsMmL1XO/sMo7k1TTvLZcVo/
Q/W+BvDKQq29/HeDxJ4ycbaIEHqlmqDm2XSU2EBKlaPdO0XeQHDM1imRJrdqzEXQgpNtT7VtmUj9
wa0UOPfoprxTHrTg601ZI1jwAKladbjI4Vj9e8ShimToENgJkVS7XcUFoW7/WLHamtbTo1JObJdf
CoMeQNBOvJ9wDaY9Kb0Cwn9NK7hPu9cUBe8WZmpicklnLOdiI7LnT78EB6VO4eEmBHgbQUvJb214
hhk07+6c1IjwRl8IV7bRGFN+G/28d3ZUFk2lve27TWlFyFq7Ts+aqxHZOTgewTICZ/dwWIZK0Oa8
DCY+zydL7zQGIY5EmMT0nCCazqVsUWS6ULRDdm5tWbnnCP6Vtgy9HInHXxMJ+fhSM6yFD4ME5ZzM
LymaNDP5RSfSHQlp3mZBSwJ6BeOyxTpdW8KDADnGLcQto1vI9abulisWtNTbmkJS2smGyFOrhnJH
H5CAPWHu2HSM4ygMCf+SbP4On+5+MGcOhFkKyIv3F4rclvtGHjghV56Jipr77KwfWp00PXY0AeM7
lFPXhFiBDaKM+y/UJ+RIfqmyHpzIB+cESsMFm130LsvxnhYUEY9+RC5bvBKKjFjRqz+GaTftpmux
M0ajzYqTKRfX6qXOGx/O4mAcy/OsQ2JYZIg8BEauvMQIT0ZhFXOiZEbT1WwCtjDX+69HF24XBpVw
vaEd7951WJYwlXTnNAKlVaZoeuOa87Zq/xgopr0odBXVb31qUmF0bTqd6Ff9g9htUG7dCAVeWZ+S
gobA0CC+Z/pPC2GKmKlswuslfYyjceL/uVsAvquU1jmf7hFpVW68hGBdOZfjUmEimFB+m2/XloT/
6PaDHKVelGxCCWykxbpf2kfA0bL1u7aB2Q6LjxTpI6IwvYF5b788W7FcOGASX7ZGhMB3mx6grMF/
oU7QxvEzi3eZNroRDVpkzHRa5yTDFhlGZwEwCTVD5UKblgvB3/E7E6GvupktOhoKZwNJfHYZCljM
cn9QZU71wZyiQlNb995973hmGXLUwMA+hVUHDGtZv2gp4yQK6OmiRwW3UuaeGvi2Ex1mln47UGZF
2LV8zmCvhBkfwde5i/sgZ6XWZPNbc16USnSk8BsO213417QNJzcKBqjMSe26iltLcZ0Cq7dMHEop
ZpDrSsQo+z9N/DCyX1eE8NbThslltVocWzZ2F6v4mNfow54tFbtheFDDZ7WelBSKFjnn/LSeA87t
mUiuqP74GRvFiTFsr9KlR1Syto9KzCr22rTrAVeU1qZmtq38vebMpBDiUj2LAjaEAaexPwG+0W6t
9sDsT6bCnT0LBcIp58b0OkMJkGx7wN39h+kzBiNcTRshE1yAVeskHMXT2C09U/0mCMFcM5ss2L33
B9D22MwaE2XBThgCQSEX25t1zZKphBA8ErWAvOFLUbuXWe5TAkjO4FSTdAXKNaGWi28ZbmcgLmiY
7+ZPywDghtM0ojtVhi+bvgjKJVmAkdWkq+K43WKzCCLs85hvwpK8ycUBL5wOKL5Vfy4S6SfcZZWr
P9sW3F18B1BkLxDJJzGR0p0Dj+/QpWtejsRXHwNirCPs/Oc84nwlzCC2qCmLpbldxqPfhCRuZJHb
VALIiV9UPyfCPfQ1Q9n7yGq3JlP6fCLcIMvI9l6aolGtMu3BOcMmD86ltPpZIibsUSocAGQdOmx4
PTnoE9prFR8mhyqjH1zTMGZUFJfz0l0GCa0puQNGWO2+GF9sb2AV4NIOXpUHp1YhTRCdYTxHOen3
mGCfQX0ssbgFm9AyAh5TalTYPu6it72NFHrOhSRvbiBQffldv6ahmV0TlvXqjeB6WWUT2F2uyy7a
ZvyG/RN8yKKHQtzMIHybO0cN4+Wmq4mpmOpWM9lAW8Cc3nIzYGacRvic7uFyX+Xs5Yrf0YS3MrvH
WRjgJotYD6Xd0kHLVVFTSz4WsFBWhM0y7B+8wLGs3jfwGXLL3AQoJVOcKGpyit5yleVpnFE3d6TE
Qr3o1RnfGxC2vXObFPSLxvQQaqC0tenvUnv+Jq2RBCorpHP/33T0FM3b06hfXjlhlaPu26I3/flP
cWwItq71/eSdTP2tjxt9iBUAIwCEVgViFzA+MNyYtRN7kXB9E2PbhTfOhYndTi4j0g9ivW3w9vZB
A7y2wfc6sU50R4skqCbABnPCrrm8889NPT731vfW9jIIxkUvrpA97K/ck+d3LNeutAmirF8XXCPI
CnYuk1weuG6vveDSQG6PFdvbPhb0VLMIBG59T+2bq0Hx8xWZiIrZRh2Q0GbRVcd/ZnaXMxh6THuT
ybY+AjpXj54MYed6e5bXrGyTmT4vS2niIijvMFcUZF79kGROgW1rOFYDY3gIk/6m46MzSnTvYPpk
OkiL7H1GNrkQIOt+ApAujtfesbgJAeEUlbEPLmRUH627zYY1sUY4WWX54dM8uE7hWJOr9bWS4xZC
Z9yZa52QaDlLUVnxfUPdJRDEJZfqEYDL1HLtsGfGWdxmOfVIBqkIM8jfmNbIP54q1qUVI9yZTGGW
otTmv20ruggdqY2JiyuLswS3VstZezTbU06Dc8Dci+qm0e9YLj4OdJmxRUJlYmDnOsJglnFaPg1Q
mKMDxCoGE3R+3T4TIml6JcsCDCG3CdxD/a4yh8BXfIym50rjXKQK0bHpztyQ9KpONECylz1zEsix
02ABZ+GVDdnxFVyzh1I0L2fWIbGYg44gRDkPg4uPSUaeKAUWgkMo+rLEopAI12f7JwfJ1e7Fwof4
leDjC1B1woJJY3MIFvtIicwKdl8yH5bGcFMsXe5t7TeevGEIT5cmrl1vQRjMUTMbEqVB0NcNGT7n
a/I9+Xl9DxrDJgDMhClmHW2TlLpzUIksgK2iK0uVxwyFI7hxeAKvzLjfuYWLru3P8abEpYSl1r8T
U2oUE8qJFr2/GDeoEaemadGD7Xk0Y3p2xbL8pOTwcgECohZAVXs531zpAeJ4kWR3edSo4GACL8/7
bxudLUI9vQwQQWcNZr/3kUtfQdflSPTt+OcrTCAmw8KkAV9BjaIaRVfyzqeSuJCwCewYeN/EJ68k
mp9o6djoIQSvQZXw5Ol1T2yHLEBdFRF1D8HME2WXs/9nJdBNse3asMSOomd6IA8O0vRlLkM5DIbW
fzJ/5BUCuMLULv0NieaYqMUrUbJDw3a3JW795jLYRjdtpRMzvMLDjiePj24ZNPTkUOa4jnP/EDD4
S8gAfUC6A395S8eu5YDFtzbQaDWUkeU7GOiqo6dTgBOO/Xgl19r1ztigiaS9n3ZLVKY0X3ZGawyf
eYQEyuk1lEsWlGktYKYecpRk5O4grBiQln8RDtsyaYmX4InpICLfWQCrLv3uEjAE4ScZIOqWgM+y
+LLl2oSNM+BMUem+rwyvbjrWKIeGVxq2fPSVO+lCcYqm9VAivIHQgp7o+cL/sir2YsXhEqWO/pnv
J6/yX0WgQBvHRdZMv9vsOthd8/5b0cduhDZ0sYz/WElGm78BkFbVnJvFW1mxR0lu+wpc1r89+Ume
yjZhloDuN3rcupuXWCNcTX2NMc33SbuFOKpgrNdXOb+ip31VIck0Vs3VgdtS1kDTBSgJmJriO8nx
8YmToz7x6oAf6PgJmQZYkWL4k9sCSzuBBFdWbyKAO82oCaawDbJL8MZPsU7Fb8nxFPHoVQq2jZsE
LvktFZmTws+mkbEY5HGkVkUpZAIFnLY2kOjvyQDZCLTWglDYBHnyyGIctzflnougxL2VKBwIPhHS
ZD9LusVOjz0xL5DhzG6lASDSW6Nd0TkBnFZ8XHVaoV8T/QIgHbt9udolght2e9O0r7O8gaVLiW31
h5vIwrWS5LhF6XbPy0YfzS85b6Kt3O2QgSXAkq9BqKtuU4ttMfTK08rqBG8GR0DuIOti5qOCdA+z
zsH9754pfYeAR+5BCFDz08rmNrp5keM99SgjrZ5MruSwXQixeb4GQa7MUsiOf9/33raWcSHeUsts
e0jCd0grPBC6g7twoaccRIP2NooFravyEd0iEkROiYR2BnoOseBOWYUkivp10UMhX6C5jopiMSUc
Yfm800JSmEyn0CflCBNcXAXKPsihpILvAS+GTMFCZYIQdCpmiQwbWE9Zd6A+nQPTYcNOclPNeHTv
9sKWoTvXTm/4HmdZJjG8HVOJUZbQnXXJ2B5cx8yk5qoSoGPBYdTt6q98K4W+stDQNBvH2LJazbHe
o7e4krIsRdxWy9u7QNYNM+zEYpXnWZTRAA0pX9YO5tXSVv1VYKSSdoSfXu0I9VbEYWwrOmKMM3of
lm8i3yOOUm4EZRLT5INUxfNF/LFBeVo1YCz5oIwnn7h9GkCaISF7xIWVKYW1a2l9fwPLjn9vGSfL
Af2rUoUVjiMRukIaW1XfIXKHNa8gUC6Y6u5yCPmQrtge53ggmfB6CsGvChiyvNBxOsbnoDOju6hi
k4cDrx7VLHvkpuwONw/SY8SBc9gwGbSbMjQwkOicki6x4z8qqzZlWbBgj0eXYWR8NSUhwk1xmYQG
SVmFlzZ8lrQWUKQ2JYMqWaHimmeXwYuLRvUSvLp8cAzX8gndkGbSoKeilPJmmxz7Kg4LZXsADnV7
wYa+HL8ReQ0cVN7QVAUJB8QN/nsqRuhCnAxcTJyROTPhAhuNroIj1bRVQ1kKG9bB0x1HHwtpZqi2
BCsLuiNXw3qAUh+t7qdes0Wgd5XdQov0d7hGnugoLTKbroyt8/s4aG2irbdXEmrvocaSkqVsqTKo
yw1V7YC3pwcRFwrIYCuAXgBnQ1hIOyZ0aTodNXeHbLAeafR6XgHV0peS11pZXpwQy33yS7ovz8zC
4Ff8KPIjBft2LbIpfO2tvdNxKI8NQFt7v0V4ZktY74cuO8P38zcO7YY21RUgl1MO0SocFZOULPzS
fwUWjTy4wXgBlZe/GlmtwwuFcLIBDc7Q6Yi5dqZQdA2Adb+7BQP8vX+DLC4GsqlpkU1HqpQ1h9oB
tMRoDR1I4gafkvYrEXYAFiWlw3mWdQOVQKqLaMp2rNMYmUNd4lsxFUdDfbebgJQOdunDp3iKAwNA
7mxsgpcEbe7Jhb9YCiCb326H0Dmy6Xkys4fMV5xy/AHGCIjFfE2d758pu6cedsPo3ekoHZKs5K6S
fFWs7J+NRa0yMff5+2CK1YcuvzCeJxMSSaXHpyi/P1Z3P39yS6adwuf92QrKn0NmCtrkWKd7evRq
KsVjGAGUtxCSl4Ayw8ZEuNWO7u9TuVa+wiQTNHxbT+AfDUo5O2Ay2XH6T453kb4aUKybgQwG+VEz
3FZ9ziWetc7d9scPmVK8w0L+5+USSKHlVQ64M1JrGhIA7+4vpko+TCR9IoB7yTUufmbDZjIfdArv
CZjnBSijf2jWZ2wgUN6lVmheqNxNtejmuyc6OZ2EK6b9/1ahIUBW/C9wdn7UK8dLyKdK3m51cw7+
uIMTXHsaMKamqapdXsYDmYkGYuPMuFZE21PvRnPjYARCLIVwqkwVFcFs47aDaoEXSsHc+8LgPtih
JVkY2AmpR+4/u1UE5sESbYRWaIYwkXI6eKOX16jkgvJoix9Q2K2hJWmGcp26p8q/Mzk5/xxImtGQ
1gbSqcNXOznPBun8NLWa+iSQdl7gTzLV5hHmTXTQy3iD8iRgZQOHGXYFu+dSu9bfRC8fQItAF5zx
3Em+h5PTu0m+zd1UDqa87aFwNO/9tmtrZ8o/QGTUyS/bSLBd75RvBaa7pYV8RI+vcX5R1Gntkaaj
7UXsUNRJmgZN5qqJEf6ceKdc0s37/E+tSAZPQ9ThccphvWigLVUT8shGzCkU0K8sKg3T3bJtZ1qT
JlTzEmHu/qoafk45hV8xwLWNMdcrxrEMRb9TQtVElHCewhgZzboe+C4JDZUMXARpgWkG5h30muRe
yZnWTiuWq7mLlksWoaNpqWRIlDi3p1Kcp/44IYZ8SsFiXMKvoLKX1h+VWZdJ+7zK1TOH0ZPJ+tiG
8zrfmdR7u2uOQ9M2w1yum4P5oqQVHjVL9gdI86ksBRCGbWeFGWmBCgRms7JIJQ7rZ1dfP+2fv9SK
RBWfzjYLTQ1d2eYJIaPWYuHywcEw6a1WOaf1vx4Toy266Qh5hOJa9zL6Y7zwxp/iaZicA3/5zrpx
2vmIp++wPEvSB08feyLcCkJ5sgU4pNH9OJm9wK/IVpqyrVl+Jf7ImmrHBKim/LHuOuNVtKQ4O6eK
BxjUoClNccPqhN2kJRsDlWkgkIe73nRB/JpGdUDy1RmADshLCog/IsR+eLtH4gMQZGRYrLcS6h2L
f++N7AoLjGbEuhvRIBqPU48hA4xzzBCkKZmWmqJrVCqeXdlYWJgWvp31BjksQg3tSMRCEo9hYaMT
dc2nXsedP0Y3io5ahQi+nJRsLa26iFHc7O7DLz/QCYkcZN1MXuWHv5xQ30BboR0xgvHrEd+t1ryh
bAZSFaP5ez1Ghu6oPiJyZUAVsGglQE/Z6i8YZkwWqX73RYJbua7WhNuA2P39dAz3psmfh97plZvA
kggskk7dKBZF8TpEMeA7nI+K7XuI0JOohfxruZm2PsbDcJ0AfErKZZ5/Bt2ARs81mCnSODiK+e+M
tgUqzj0+sFqDz780uODQqBoJgy5e7pjAx/wT/ETG9XHAYdMEs4Tlqdwqa9hfUFI3mGEP8C0RDSRq
Xui6h1Jbgwq6ApGGCR/5UYD61dMK8tAJbEbzZlyXbNjS0qiUkjNLIa/KBnwyVE+3zrfY7Dqnlm9O
h+BrGIOG5afLoAF0NrqZRIVqDVMcH1d71aEumDrul9H8a4Q5a38ZEZPEt1xogK61Mskv0LlseSpl
D8yX9ZtOLWkOseTsqhaU/CxpiyyzLwNv1+1qqzJ+ASVxNwdsvzbyc1Nuqcv7uOkUDMQ1SIS4Jf1Y
BK4yozI3m0c/RLFEt4LCZ4zDVZWQkwQGu/P2xMGWD8kHrH7mwzNWOj6CZew/aenr5zqyRv/G2i+c
zQnhOa9kcOb1/q8gNWgUr4KdXut7DeB0tUeI8AOqiP1fPoRvF7TO8dvxRhEovxyazgsKJNkXtKJw
WUu7dVUcRRuUEcrOnrikl20xjduLwobLeKTcjF+g7R3vxAyoQmYYg6Q4u0H6jhKpRa6tIKzqTxDn
mkRr/HUHRO9KYb93zu+D8rS7R9Ozuvb8JNRNunMdc2YdJ6SyT3fz/xxTtU9CoFdmGK7qi/8gnOy2
SBMoqGNuMxG8BFaaT+UPtZT6k5EEdTbZKsKtlq2cBT3PQ/1X3pwX6fyE3zceWInOEKS/k35ErVxh
zm/qTCAahho/hMtQ4+grU0x+mQH3QOq38ZXgXm116VQ7bIy+2RoLy/BAm1QK6PIBGHGcSt4/2DQl
Afob4NfOy0gTKmkoUSihBd69L3S6muDj1Osmvc9hcFCa/LetzSBz/Q4ZQBrutgLtubKaGqdndFfi
5ueAT+X+39BmVltEHK3/FZlYRByy/Brzg6KXmrbDykEbRW+5MYIRmHKSw0sYZwOoEkPOZqyHQfmR
oDLGCpBlSl5KMNXvkC2Q1fbNeRlQiNRdMtdjzedHqngKfTl/RUS6MIvE5QqWzOW+Yx5pVWC40s4s
Dyn0mkFddvYO31NlIOif7OEPbqDAIFfU/cqpV+2nx0Lggx615+CiAZK91C9QT2K+NuiTb+1Vc3cc
C118hJp2IFpyfhnJ5W4/LN3M2jdy+a9gvtzxZAgjkQKnV1LMN3m+ZIxvxB0iHKqvS2VE4gc6itAm
MpiDrCZpUzheWJ2p6GGnZ2ic+737dMd8H/lUknBhn/pwOaMN9AVMsGdWJqQLlI0KOEeiA7mxPJwJ
4G0xI7hn9ImESgguUXfNuSOL2Euo+5lnKD5Cwz9sVuJzIXuShNTfiGE05IP0on/V/RLS4f3qzQca
6ECZS+TfxfqKW9E8CG3YEvArvSCmsbsNXgHFuRUqxplDMY6wXt1Pe7DhHLpnR7DCxbgeXoBVMheK
XCraTSnZFbAvtRXpxiEXrn4xtddd7u5VLB/Ej4NumABvUAoDGCIKm4Bslvq4nkTbNCLcD1MlIHca
bNFkLk7SZJRXj83lVrLAQxTIT002kygICasEWUAT1IsE3KCYtf/BKFn3xpBiR0Mu+fRWJ/FFSbfj
GAlCa9OQY9fE+730tO/CerrQyJrUbEJC1k9HeFf8pWZ3lQLPRoIr0aO9A2iNbhIGh8ZtnArvLF3g
UhsjflRrimcb//HzsleHXqo0IyJfIvALkmvGL868NCNIKuQOaxjbY6ei8hR9Pnef86oZQYXS0xpB
jabPoBd/mBLHZHRTpKGdLobxRL1BbZJ1LlxkaSfds6RC4NsAr7ur3Jzs09RXy2OQJgTvzkxkolaZ
v0VijAyxqjbeboLRwtGAvUXYb2rezT6+VGNxmfMqJbXFsOGcHsIGRy95j+BMMr4BTlVOn3vjYP1w
HsCfCUBypM+Rc73InxAsJvGt60PsdzQB65ZPcsWXOwET1V0Kf0FhqyiDBp+1pHJGIqzAgYBSg7Hs
WkPsIkNbrDHFODnhoXtRwYCNAndYF8qbexgUUFOALYFr7SzU+9B6djHljzei0Qcsletj4BQ3NgyY
9FVSYQCbyQofRk60ZsCKJMW4T7W2wP+R6iST24iWYU7ofArldahQIeyagYO6rKY3MqyVZOJi+DmE
B/dsiRhUOSZ4q09alzvFU8SrY/ftM/mtJ4FZb6L7Kb5rbOKMzSfsdo/cRYjUMEHAigEteLq0dmJq
D878/z81wucrpEGk5crrjWg4yKFMHRKZsNHeiwIV8mU7/hHcpHFamdXlKD25K/HmqDv/Of917aEp
wnJqWP5zosa4/JaetzYOepDnVhGJYdgPVQcUBdQ0Lfn8zGiBtks7ssDMWdzyXkor9y0FcAjW/HCF
IOCy8RWqI0mo1yLQGBDywvgsG300trPQWEeoWr2mnKozc06aIFCJtPazVdXvuGgrJSPn7/HHlZYT
LTSvo87o4gk26TPdFv2uKTfw7mvdmFjQvKx4QCXtLzs9OViEw07gX3thgj7/Yoeby1ICUGON4pPJ
VJVZXTLUpCzxeRvfBIAacklvctZiGlVfkdu8rH6dPe4yfZGDAjW0AZWG8M2D+8TOYO25XQkEiqAN
7R+U1SasnIR8fLiq7V6n9R60mgVTAvS7o6AjIIrBZXv86Ww4NBNi1EUQgApQCBQHevq3ki/5LACT
6On7IkwrPXAEYHI3ZYuEZQ1np7Qra1R/jvVXgysBGX0GHAgp+ek057atB23eQCFLKfGcVURAaYcq
1lPKtfWTGWQxqwOkc/whvtt2A1ZNo7djBOLaZyVjP7+Q8YtqGCh4YpcgA94dRpPwmCzJ1p/37N4V
CG6bBg5ClFAgjEbOo/JAZjM3A0PLhB7RGdD0ZSJDTQOz4NoVo1x/r/51cKSbof6HLwjHrz5fcQnt
KrRibaW+qKcjdDFq9zzcx74tUXQsQmOVJ1w2lH31Kam8OWw1mcK+g2e333NqSzf9CTuZP4OPPwqo
quVnaWQ95WsUYjRZmrlYXsVXNBUo+KF/MidNuTVKaaN4+DoIQV1J9GT0r5ii+PdXcnYQXJx2FlT+
DA6pUkN7+UR9Dk8GxQ8YN57JEOighccNmyA/rtsm3uNIUj6VcQujKwJe2UUqXztjmm01IxvtqKHU
PgDt2ddfd2vpQ7yR6KKl1I54ZigNhMTohmoXc6Ci3b+m5CW7HOxSpRsj/oT0uXxupn1FBEzJZo3s
ejt+R2ZoQSJlQSU+th2jxwphS/yly0TEnm0YQU2tH1GIJv0F2NV9F9IaOVApy24eRSGzloNaPkS7
ddkx6aaok9QV/DGY5Msuo4pydCvjb6NmH9Qaq9M7FZE+UwXRyoxphk9FeIMkw+0UD8WP0cMiOEGm
FhF8hQFKHtQdsUg0jBMQkBlhuyDQWdeUwp/MvD4EtsZt4XJbGGwhcZn/OkDibIFNvh39fMArGvPT
Jz/DRg2zsKo62VV6iLJv9xAGYrhnfLsJ8wPil3vptLY7Ta0iTu7hbXoRLt8rNOE6dQH+9Nbd87XB
DFxXVxKA8FsCd96fyz32Q4UNSfRZmb45my+LmV722j6hZ3/6L6Tey3joEZpkWMavxcWxEEQEfbkO
kQKLfdaBin8VZLT32ExRyo8QUnXIAHdlCBUtIwWTCQWpH+0sIWysoYk1pzI7sjn4zFzHGftiZV5E
4lpieHGtqQ8XuioqieRUwWgKdtvJTONa0XrPpMwJKGxh6wa5BWGEUoP1aaPQBtANS5YSLmwbJqKg
EK/HllFZ/ku8sY/w6++vMV7n+6hcKapM41dvJ1k3lgFaqrsunVzCF3sS1lcebZA+DncFlNRGbDTD
mgUVo06r86Lu+Ih95PkRGwRez5n9hb52PdbTS+y68FXnPwtg+8eWuSfy7oA8S/i4p78/oQEGU8Un
p2IhW9naWlwgErC3GYMa1BU2/HbJ9XyNtAbiWxvgT1vBvZdwZcQhctJvlDSpx3umlQ8iHWuHowMK
BlxqWdcw805XiuK7Oblu3OePZ3hNK6b3kARIyVs6nvblE0QNOVgzYm7e6WQx0Tng5iQu0jTJV3MY
rRQ6V5lE0pLAZF+wVHb2EaCjXGRmbGDhyvZRwS8bTqHQEja7KiCs0Ye6cYaIriz0YHLf27BlotxC
pzZKQKs/YEaF1kAsuQVnpmwTBVGprmSguxDZsMdLdw62rZuzJVtitPG1vzzKqlTQ6AIUSpvwD+1Z
nUM4JhKeUgEg+ft+hWlfkyA1x25guCgQNPbWN65yVTOb3J/vo97N/d2EuatgbIJUxpLsgbaHPgWw
nMylH5OcL3Ivww7xHI8dyWI7HVjsLQy6ydeTqmZwXCAaDSUZl5Eqb2pRwFSX5xC/msDbEKXqKCu7
VI2Wb1SazCJiHpqc1Gd4xIkLQ5ty3YJSgXKLTBPcClUZMazGV68SYsRenbgHW7aqLw+KL4e/ewE5
P3pFB+vWzmdKyoXXH4g9nwYgvQMSZaOEht+8jvM4oMIG4w1xnUISadrKlw9FM7iQK294u26WEyx9
xaZ75WU+1pdDLZFUq+30Q6xHOJQF/Pbn5beVMyGcn1GWxA/oxLu+1mIyRDD9T14CyJkwBHDLAo2f
q5Qhiv1A2KJPsulKS2bplGPxOFNk5mEy8RAXDU5RxktHRbJKRLh+bR4DsISZ70QoLBH3w1MCPPVT
B0IOT6JNdTDeVXJPCIKd3f7T5ZSCH/1fjySQoqobH81bkK4yd2FvUKMIT9BbF/OgB+eQqVx/dtCj
UgfEKINdeiCUTVQnlthHl01ic5HR5Qp6jj1aCM4Dlp7ogkPMuAHyJQEBruWKCvy5EX/DeFQBzmX0
NNB8KZiMKp+3cYq5gf04tzW+VBql8te7k5GFRSvnBVrueAS4rOlXiP1YseRg6KoTGdtFd3R7RFl7
iDk81M/ikSwNkToSh3T/1cLhWMHsmH40Bp0fdob0BtDHdfmKvmGnj9sH3NdIkWsSV6VCzNeWiAJj
8gNOoiqbORz3EBe1QRHdT9VUcmkGeOM+sVPpUsFcGSZSXb1XGpXobemM5c9OfwLicCvzaoCF/wFF
fCWoQVXQG+WsRiaN0z03dVZX7zXWCjV2h8lOUzbBXz507y4kb3g6pyKXSOjWWmrvuOf7dZ1PA0eh
P1aA+/9RIvUomiS0Ug0dqAz5CRCgVFLCTmDT478HRGhQ90px454eEVCfBK1fec+IHmn9Nxm+gijK
x51+S+0PVQ97+WfmUgEeMdSQE5kbYc4mF5GrdHBrSIpoWk4mVGBr4FPeFTf+mAvQPdNOsc27LFe1
QqL+2dBtgEboUXCJwC8o8qeniTW/gCLGgTWlD3UWmjJ9ef+VarJv99AR5E6BveG04kpGTjymhdGB
a5bNwONIopjbImx+pxU0vnzMyzpd947f5lsK6qQJJIkTInkOGGZUXs8nZMwnlTk/KJEzVE2MTlDU
dYd8vORpGJPoyC3dSPmMCWVHTf98YYO2N1psmZBxi/SRH1z8ADlhQ/slBrjwEt243JCcw14d8v6u
LFW/rHRshoxs84rINCFVbLYp5A/hUUaO0d2CShCh9KAPlJl1sSuPn2ge06VkFg3D1r08F8grx8Zx
UMa78D76DBZDK1TmzwFjuMBqj8OhdFidMS+Brufm3/fU4SDMUOK1tOT0nh3nB2O/5ITTrvP5mEZp
YSWM2w6uuInmf1AK9fF/cF4MxeIHG3XfQYEdlYaXlbi2vvmg6jZAkXVsFsFKoRMSIND1dcEfONVy
cfh4/HZVPJ4rjUKY6VNBVGfJUfkKsFxvf0GFQTImxU9OnA16RLlVApgeA6odCQe+BXUXirmDVGBW
H21V8wG+LsHhnt6g29F/k0XG6TSy5UwvzYqWwHfde028Cn3Gk5O0mciumxwVa8wiLN/ifk8inU5W
WjMxcjNNMxuzBlQxfFiDcX8zeCcht8b+wTv56vKEatUzcuR4UDfics17Y8Rz5Fr0ESidptqpxCs+
LvYyyVXet56r2+gdhPt0QL8gFo/FDFr5acFN4ysZy7MRhEP6pTq2W5npm0J1vnJEZOqq6KOStXm4
WAOrIZ9eOkYpDxbvLBUEhE4uR/cSfIjDZknVQM4gK9uprgodSpRWJeIP7R06tWNe+1a05Rzs4h+D
1C1j+T6guFjU1nUjkv/Vg4SloQfz4cELD+1I4o9u6v/OEkc4kALsdrynCuhUwQIRAC03nVKC4Hor
BdPvHY3D0hl4hWlCfRqdyRpDIbFE2DhtHiTjSee1WPZn36RQzTRmLgbWMF9aZmBEBskLl/IiDes5
xaDK1Chp5bDMpibtvesYfGLTu2h+Pqnwp73ELQFpsIOYknw13kR3lpfX1jZHlMrDIlIT/vb+wLU+
wkJ4Paue/2UdEM9DSv3VOlmUwAOtxXrRSd8u+Wtv+3yl/IvVuW9/pRMHneYBO3vrF/6E0H9czY3V
NGexs2o8WBEhb/8uMtXhpoTeVoOROFN0Dopv1xpnOGUzVL5tmJcuQKqkK7l2tSl/PZlpXDba+t7t
/KVaP5XQKZ7xqDfJAAvWS4zU9IWBaTAvc31Xhs3518wtSalEeMylPcKg7drqgJ2jScFI9Ad5ZnZL
PzrzoWeFsztvGnBY76YcrpQEVesFcDHIsfiGBrAe/3CvEh8naQsnYtpY9anU0NQXnmkBDlxXEVHM
SCfMJTDM6SjIQm2k+J7Ud+sYhwLrxB8Urh1d7DDlf6Y+EqVSiW2q6Qvo+MX6IuaL+POC1vZmZMR+
jBT3SYKGD4ZR/XR75Y+kKdvsUdrqQ5qjiL8Bi+/+XdSibnKh1Mevl1YfLE5jwUZTdW62RBDkPd3G
pWbl+3aKp9sotwdWNyMk/uEdL92vCYc2CrSXDKIdFF+chQR5sSCr9D/2yo4iOSC38kIKq6CgPQM3
hlt9vnGUOvvf+HKGj4g85dN6I7OMWu1vg/A9wvYc0LAh3LYql4sBYtc1bCAWIeMNAewgroCiaBR6
Qf+mS4+ivXojK9w6uPEMTQOmIwsv4OISgeVRY5JxaiLfgB5r86I/GwmXSDs9WWYCwwgunXs3F6VH
X2/F4SgKPUFhFol9+1j8LyiHIZOP3kYSRsfn5BPMfZv9ILeUN9458HP3TnIBcqjN5IPhhp5woL99
l0vyrtwK70G2fuPqQuSlAy2AE7O0HNSAv4ECrD50UMWdFa5WTEp6N1pTpo0sLp7hJtFbCgBtrkx3
KDhoQnwbuhnNpXbrpWrKDNCNOAIDgz5a8AbPNsQKV7nvKucUJc9TgAzFVb5+zvbpSPJTIV7HC7N5
ou//k4DUqQUDmdUvYcYq3V7KlBKBWL6MYfQTmTMKhEItcNZxtCinOKrdtOnNJUVA26ZdyXxFEec1
ZTszPAPLITn2i8upDpiP1PxzWfDEXnY2DEU5fd3sXfOCicF9ofD545zCFeWHsSM60jBba2op4Xtz
jDNKC2QjPbDOjsZ3RLP4I2j2DqTWauYKKLpcDp9NOe26Rju6pShVl7FfkT5+g3ROsb/Ex/lS5eiO
5bhfuRVySxXLGi7OQqsLqngrjsi2W8i74MwFoXPlaQNsBqC7R0vh7JCwPRhxL6bWxqwSfnzDXtf6
lRkJRd2Nn4d+vjuOcBlfYQ43JUKb7sOIk6ermax4V7A6EQal5yOLK17ni2AR/V/34D3FxZLNNDPU
DWW9ojkZwPmztSMvkdZNHGqx2AoVkEmEGDV0/2OOQFNpFAmFNk3hCF8JKlBwEDKZNBJyCAcd6Iie
BEeLv2CC9JBseBILJZE4fDLUL4SWiXIPQqRdmXuiefkcgC7Slw/PrXPkt6oSk5WXPYzpP34YfZ2z
KvKzBETgEPeeEcfcwF1G/wickVD50HRTAdXoCmvpqyRFXcB7hjxDYD5B67qtaMAU6oz0QkwfI6kw
Cv0y3lfUGDayn2B87D9ozmFPJVoImp8Xo17Dy5E+fBu8njAm0NKB2cE1Z4JphjsNKu7QxqAflPDc
WhYWsDS43igZRZU5MTpzNXSmwaXhVdHqIyeNkGfaLLT7qvv3Knt2EFdS2GUoLZUku6HDW/MGhaAV
aJOCdODEnoxhySufjKFYidvUftH2ApgGKf/+SBoLR7bb61fWA/x0RHqBbW79bJeEDwuTt+i4dmuL
V9rbKUwUz1Y85dcya+TUI3lVG7qhuYGsAjLcUXcJh+zEniPtijEsTiPwL7IdU9jG4rrSnIFnZGIk
D4OdIg5BXT4XX5OtwkFHGytL6or+KtF53XnEgHGv97UChTZIw8SoeeZXiDV10I0Xf3GRw03QbNFa
eW2UgYBfvkZRDJX3TcryT88v3MFAqDiFgawrbinVvL+OZW+HgY3CKpXlvL59NjLalvcGpjVK8qKS
9iu5rEudxvZQzIb8zL8m36GSTo8WdtQ6bYBIt5ZGor9v0kR9RmbfcYfP084rTEIRke2Srb9BJOu9
BtouSLZ9ty7FLQo5XdiC9lCASyKEkVpTOUq75LvbeTS05jEzpU9jYrm+KV4vhCHGX/RKwYolA4G6
/sDy4SpzQei70S7MiG1pvE+S7AjEGRR2iP3o15X6ctnepoq8alIx+hlZENJWV0OlwLNBjeGgjK9I
Jzscph5I6lTfjcpYIlNLGS7B2mNsS1jC7pL02PPKiS1tjn4fsIyG75awIfVSJNxnyykt01li+C1T
rniFPZNir1D1MO30ZTOyDLygE4/0VSHAYCMsQetDbltlCoEl0NKi68FR1jv9eKq9OeQz60uy+lGD
jzl38Z/ir/esxb4aqe7wvwnhYM+SHMw5pxmjUMdAQOB/nAjPKMCyI5EKX1YQmOwZejhNzVjvRPrj
y6B0MzMQJjwbhbHjdMxA2xw7fthPzB0TvCD91zW6IilxMMm0OvG302bGT721hovxvFjTVlYMsFOP
9184xJL0JprcnesVqYBfWf+FomuFTzo0js7+srOMptE3JShZo+QjutFQ2N7E2lAri778CQOLcKcK
wXEFR0pNEDCkzNA9pv0x5wVPCV7A5pspkDuT/YtCOyKeIVcAWz5q57O+uBTSW0gwvhkJ8tOOirhN
Yfv5D/kjbt9R9J5b1OQmfDow1q4XNdCR1lRpWSo0U8ReLzdFroKYNVVWV6JaRKj/LZX1cJbdOLKW
7yM5hybPdK5toTSRQR8JJDc+AzyEH6ErW/UYGvk/hhfInzm4hkYoban6+uxPF2vZGiVx4t0JdP7o
ZhNpzqwDYp41BbAJ4ZOUX6WjgT8pDNAaDZ0mvPJXhooxLti/LaUEttRjUyCNdE0vwndr0kEFGaYT
AFNWQ/TbbB7+qxAn2ruRmZplIbKxo/nGYGxmJ4A3LJ6vBUVxMJi86fVoV/7zCkkEUTci8AHO6ruB
kzawwu7WFMzR4feURk/0kuOh1KZANTR8Mfrp6i9HzhhIXHzleGQ21f8f3V6WwGCIwAa8SARLqgOB
BjToHSFOVDdVvcYz8iL3tH6wYoNJUA5HsgPmfUAbwnxMtvnnInbtLtHEUbYDJ3knW8uxyhJQCkNK
OiwcxLr6ouxwyNQXerkYLwuzGnd96EoUZ2X2Ug4lKf71TVpCDfwcXl1CHWz+zisKP5FMQtz8KWtC
8nuokB3s3fVBnS+qrgcBsGGjfKkaQ5cepXewtLIPiRFBGWVsdpTEw0SfJftepyRaXlVytH7x+D9S
sC2MMTVuBK1HGZ271W96+HBp4GzbS98mTKTwFZWGrphCKMGiesr3tJC+9/sIA5HbOQ+4Vb+aHDjC
dzdfTHgqC8TwfIpnkWW+rjXt2iqGqbAb8PJvV/36P4NVEeYhgAMqfjauPrp8Jvgs4oycu0el3/n7
6V0J1Dqfx49GE8swJd3ZnElWsumFwtgfO/PQMk7oZ3fiqAxZ2r0o1YkTdf32JYfFAohGbs9dQi9b
9qi5m8Tn9PR4NV6FHIZ6nAIfIlSQm4ArTRrCzwXwK0Qpkp5d46V7vwtSOV2gqldhovE3ikWE19N1
O2CPeWfX5Ssekrpx3qh4U+PJSGvpFfo17JxegnWHgDCPkJbaVGtiuTQX6ZAbpu55+P3Vg511AvVd
0LAyANuynLs2FeclAGHeNCjEg4KfIuKEF56H2eC1tYUOHotERFH8U6wQkOauA9jMdepyUSE2k8L8
xpBlXH2wYY2Ftz9rh//GvPEhsZX/5BcxzQg1n55cfReUlj4jDnPz6yEZ7CGMNmxCG8NaTqLnHwHB
CFLDpwEb6zc5xt8WVjBNi8XSo5OJWSWkLiQFzvhC+N9sEpUkMByxaH0XBI1RkowTjs0tMyjQUdmM
ruDV4DhJkzBz11EpZfkKDDSY0Pz2ly8L3xGX+LE0TZjfoNsuEmQrr6/Tt0xRFTOyF4udbOnMVksU
A15ef+8/DUA8NMz+81I+0fPfb8vgsvxrSnHpDicawuD72y+3QGkkzdZnkvZ7Hl5hhKmpWUeDE0jk
FjbeTuslbdBKuZ+5SKEMHphCuXF/tkrZesgI0k0WeTIYnB3JWwxPYLj/5OM2DaehB5zEEpY45TAa
8vo5/vNXi2tGYrO9KPRYMZnI1+L5Cn3MkMxhQceokRZ3I2S1/G/fGn3A3GmFecrtAthSJFoxRre+
iSEIIHHlwip1JndBLsoeFS5QzmQG8XZ8AG4xYkszDw1t356NDTK9NHyQL4BdATFTVQb3kWpU1Ock
L1ZWfaIN1A79T9NzmpcKUuzXn9yxz6uPLujamMuTzbFbO2eyPwK15V16T+6uVp1bvOmtss/pARWM
MAFOl3ux1RjfeY5TrcwueGS5frVPbEbzMk+UpWy66Al5gicfpWRF9ZWJ8rH4TdusjWEA2/T4UjGG
ShoaWly27hltS1HbPMA7oUZ2a+dbZvP1RGbL784qKJ6yPYBxH0jBuf9om99zyPZJckyWuFmsQWX0
JP1OfxaQCZGg/tEacMMyf343J2+K236tg4GQXx1KYJQUTLrUwnUIL8Hqxb6b7nxh2+H8caylrFxt
cXn0AVWnKWvCtQqXxMHi8AOKWUIc9kgfnMFG978g8Px34GkgmT1J8bzay+RJa03e57KIaYioCa7g
0s4mokwH7Uc1hRhk2r+fPsmaMn6KxfLkmH/Nzyg10nikLxrzMhNwLEEnOdKxKxifxe2suh53BwM6
89QpNNzJXMWLLg+mwQYX8tafJV/p5WaFb/nSjpMKlTE1RAW+crdebIwcVwHs90rZ9kzRH9Bgxmiz
bJOyeruOrTCU/xsLSe1PiqpJN/FTqIaWMeIXKkdTaxzN/9oh5gTCwtQ5hyff0V5FLkhd/fg0xy5r
2cy/CtKX/4KUMj5DbeoNX5CwoVniKMbTlQlQB8j74JcdD6UGIE9Y4UvLw2QeB4dVHTdph2InQOWx
dnFE3ywZopi1vuGXDXSYbPlhrxJh9ho+tMsT3v5BvMVTwnX5pQVK2PrE+K2v8UliizO8qTSMkC1x
5JbaF1HLd89aWES8OkYtYDZpkLE6mHXOatVi3yC37temY8jDrvVFX4/s2K4I1ri8OQNylujV0Mge
X14QEYQNfRa7y8+RpCc8Ipy/HrqrGmMjZ8+JDrCsKg5p0KRQx0CjrVJDBR75+ISkYQ+vK+mpRVOH
0eFyVGOm2KBAhuYfSXG0lL6AvK1nOPeABuqLt0f8BosLfd+LYvJgFVEZ6TcLf2Uy12xpXe9mgqZ7
mDSrK2W2KyLramepqDK03yPBfyTpT0HSDHlwS9U/iaMCP4Qa/5UP6s3YNP1ZU8+TEhJVQqGmGPE7
GpdOB9JH0E8y3yO5Rq+X1KKz1HGb7QmWC0IANasro2JAyFl5oxt9LJDsEPtnqkR3Sptgs3K0K6BS
/wmuY/AWJBbzogm5s66RDhxOeC64VQHrtKDJWGt3yZwf6R3d0GiEoxOBnIcqnExhKINhg2CI4Moy
3vvIEISdFoC4moJKVrWC6fHHZ9AJcxKwtY9idPR7vrIB2/Yer6RR76DoL/Co8aoKIo4aKOO8kTAU
Hn33a54iDnzl7i/8HW3J3rUDe1uf8J+sIGbqBMRkGrYMTqS0AVvFx6MQ3ejQWuUHr/imN91P88xV
W1ybecCABtRajWp13VwMt6GTFdsP1GodzGi7IRO9Hvx+oyiO4kBs7WJlqZB+vnBSVZwjA7tx0UEl
uj8/WQjMF3qjYodMOuWRTkPHKRZ6eW95iGwBnnSwv4n/nWAanSMU4m7ewDzhCccpno0YnNNZx+ad
f8gJ0LvOQW12f+LT2NGITLru3P7J4V9V9UZqefSy/Blpd+K9jG1k+4IlXMI1cFma8sSEsllZV9iK
7M7dsLZWKOoJq5hD0sDlig/UFlXUg1mQZJWGxA0DHiWpIHAx4bnS6k/2MAfXp9+bYP1597YU26w4
O1wgx+PPUxwuyYKndMktn0ECcxEF2ggydMSeiLEuUNO5ZiRO0L2Ky1IJCdD8yLDo8ezPynCoWrtk
OAqbkBQaqIVgS2ehN/SZH9seymuH9UhsHHn6BOcis7LmMDMzRK5ummFLgcBNhrpkTZ3zjL2YPE2Q
zO3QICsVyUNxuZunzgOxifvvWGFggxMSINPMoonhnORbOdpSaTSD15HCgKPQnywRm18NbeBUlvmz
FmudL045r9z/a4W/CfDD1Lp6Q/xGfuMZNY7qo3LRwXS51BwF/4jvknqo2HB79MytDLnghF1hhC0H
vVXiURrqMHP/zO/oPwWsLLh9pkwUfnW4BD1IN0b/5nET7NX8B0JEDqqKKWNp8KFRwAs1MXx16jjt
j0eXC43vaSGy3Tn+swlU9TmV7YfSH4fYijwbv/BRbNKYTLFRnXJf7HAS8pA8aFQdXd80Vg+RttEn
OlMTepYjRw6IrTGUIB1XQXYEGa6kmKSpgnww6SM5KcXAdndtPVZd4BavEQMOVOO0AvPJK1WZGdvD
1w7zvYiYPwrSZCZx3bGiwJRiN//wW+aWkI+iVJGPc3UDVlp9QV3UvgXw28bNCj/BFhDeafBkl/zM
CmjWp+t+LRFSS+r2TVZW2H3wuKjI7NKkHpy/a/2N6CUyTNunD/oF4Z1KOLbBrPtKFvTRH8T0jUhy
vWWt8aXfgAIZjA5I38Ky/1sPYN7XvUhM9sNlrpaYThY8qAcIz4SEA28vo2D0v7ZDZX5HILT/NO2I
x8ThMitoGJqsoW6VMYWYwwyHWE+CuCCvEafxaq+RtslDi45XrbAC4/7hzmvZMTNAwQBHYGyya5tQ
l8JqRrzlkNJM2aKsH7Od5fKg4qACqsMiIlMymao4eDgF9wfXWtspZpfXf81cvtkTWpUOtl/PUZcf
llo2yuRZP1iyzxi/0RnAYGXDBg693S9AkB4v2TSsVH1pBS4DCVCWJw658fGRF/jcJlsSqJ5CXYwu
u7D/jZIBF7ezSExtoCvQV/IUGnKAXnTuhRMdmah8QhtZ0f2rfOKFuXIixKgMJsOZ/2sOrX56SUMs
7C1xEwXGLpDIU/0JKS7fCJIbEE+sHkIapa+s/SGzjKv2qPVrrcUIskG5W2XZEp7IxNHkuNK0MrE0
IeBIjiATLc46yP3tFh7gxwRzyOKPshnHwZaKfNVbKdiic37Qu8JEPyXEdeQMCIVDmKrC2xZQp5E9
wavpXGbgam2T70njRr4GN7yNyJUk8vgEkxkz1BeMVvSlfLdV6VyCiFRxtGO/7Egp/iXtMFo11HFH
RbodW5pLnm82OMNMZ+99a8wiMEX8jcGiBCdM65ubHE+0hpKKqT4GdZhBUPPfXI1FsJSCQrScxyZh
QDq/WkTNinb39h2Wi8Kwlb5zdfSvNuNlX6dIOhQFwvJjqWk4D04WCw3QBXLG4cHGjlVzaHUM9G1F
U7GvYWGW5GoJkxex/c4GpdKD1K5xWFAt0dewhOgfnCtc4apzS5/SspWTgPBri9E7Wqa6wi0cQlhN
3KUE5ipC3BdFPjWvfSZPR0cQgbS64yr6bHWQ6Z7O5pujGaFLwoS+/hUctGUIb2W00fGfL8zUP1QY
/dCfpUNGqinAPObf53nvqtO3ML1gfO1pv/EvO3JfcmBzqR7kKjQCLOEh5uLYb54Bs2A5q+iYN6uy
b7a/xG/vh5d9SglNbbKe9I3F/sUAxkVMBmWLVHgaVvbsqIf/Nu3H8rJqHoraeEC6eHNfZeN7amXq
3dvpgP6QmSD+0IWc5HyrOvBJdXrIkcjR1BNbqDB4ylkvelw07p6kXRDdNKi196n5i7CZAA2s+2ZE
36d8OjpE3MTfEkuvfDs2SdMSzpj5srxVcnorWBIKfSgNAMTV8f9vo5x/jNwdwv3GQMzwtn3Dvu0X
OOj0e1Ict8Zcb8ZEHXXBwvZrWuy0WNqenZiRYIyPNd7LIwM14DgOHcc12gbeakGkRn2Rl0XnqoqA
lBh+5Ast9KuMSOSH8oluQgcxeHQ7w158T9IJOLioELReUynH3TfkVxLXqBhugWcQGhZsa/+tYp7U
e4bIftXQt3lDufVkiVYPKHxo5WflQMbxA5v8vLcNZ/H2xeHxipe8rUlamF0GNSQcQsJhm+9+QVJh
mmW91UxnpBVLnbt9gf+xlNyI4Iq/T1EPBTbR5zgSS7np0d7J/ZXPMYKBStZY6Si5eF9zZKMh+GtE
U4sjbKhgLF/uvQTZ5G17NtI0zyIKKcrKPe2d9Nsw0TXCH7Q7Kx+Vr3HMucbrdV5tsNkHJcL8UWn4
iGFgNIJ1g7vYgiVx1/AnVIcBSSQIfDjtCzECf1B0XXDVXFF3URgp/y4ZMhwHOIxKh/cHRVgWu8J1
r/LDI9iILV+dfaaedFaVuUHqBO8dXOYg38kwnvHP/bjU7/uGXRrj4cUfK0Wg/XmZrgKBamG+72Dd
/Ny2Msl+oI+XwxQnvGkpWrzkZen1P2MgbQuYEWpd1rZonUpaiEBx7BWrSP6DC33DEyMEQRHk9O/I
RrHHkXXk/w7wq08IEaX1kTJ6bVhmZHNlClnu3rpg14AB7XzkHHoQbCFVwpohKoSGa5TjT2nDaDzE
cS+y7vOHc/ipxHWBHNyjgoU8RZo5QXlJXktkWDtraQyKxBxMVJWtGjIek9owT3dW9JN3G8DS4bgB
EEOhuK3aQ/b9GWxahh6ocYI6gEhI1L/Z/40uU/W6+Tc6g9yULqW19PMLX/CcsO+yiI4wjWG5oKoT
3xgEF7HgEjPu+4eRweyNRicRsysEIcLJOISGi1M7iLOnvRbL/ZX4KL5PRbSDs1pyZePW4Dvc9AuA
+DSkoxr4+UZGL8KWQZiNML4UcbPoqhUrXhzQdbT/oP+yO/odQszsb6XPBwUvYDjoGcVsKy+qLDdr
qOTGTpmKrx/uPmeY7vZEcy1mfMeSVFD6LmtcPaHd2uY0urvyuuteR22rWzOIWsZKxHDOwjdHROfR
FM3WH+a/oe4LEQrf1fDOkB46tHznFHVaJ8vQQYnlSlEY63/U3yHh22eOo8V4r3CfCTXt+KwWyt1q
ZEgjT/5hKYbb3d88GBOGAeqti3EEVyFh240EB47+WO5Omu2+uqY86iw5Nr2h0XAKYT5gNhSKmEEQ
qDYpA2wLT4ggmidzHlI8woqum6x+2imafgKJdhKnmTnpS2ScLBU0vIlqTDjFD58FJRv/TCSlh/Hj
C7hb4JsI9HBGdobhECbxq+QVaTtU5Myz64CAeGBCGtfM6qZcsDwbOqKCAqTPOb8tEk+BcxOtmIED
iWKVir0uADqirX6lnKLGMlKgEfQVplfiISLmVHJ1SiEIHHEkSdkCoVStr9RU7PaVLB4wyzmdFTXI
AfyMSsGLMkFoLVsSLyiZZR6zo2JVxEUjmrMdBt1n/iuhSq3XoHZVQ1f0L0oRvFD3NsjKcaUQDA6V
A/AUuQHxlhljMfcIVhFg0rNCXysTYfxNzsEdSqgEp0g/UwrvU90xjpSnLXedGBbhWaMYlDTnlDFZ
txLPkX46ohI5d86s/VIGS/EZqBBXmvMJGfDO6r35YiimJpV0cKVA6d8C3moixZcMGExxRstdE+m0
ti0Zh9OnOq1B/27YN77Hrr0keUzlh+R8NxgjkHoI1NJvYbYkWfDoVX1TkqGomu8ABa1aMh+glzzi
4EIVDaYSl1uDpdB759a0m7Q9Nxzcan7uVRKQr2dDqyzKXuVDUHorsgZtbbrqbdrb5RYNvxqAOaIX
2VIHUgpu9Lm0yvBGxoVCqcHP7gIgijaUclcj3inDMUPs8DqpkV0UTG+BbjltWAqrvKzVk2HeR143
jCo4HT+8HQT21xMXrByDwJyJonvPK0sAM2f+0y8SiqNCok7K/z093xqeNTh0FC5l/DiUSMp6KD7X
5d+FwiuI6cgxJuwyjwMHt/VGz2f1U+S3O4qXGY1WCMxdpYF/B6wf/51tmCH5sc9o6CySbcQfqFoA
JL1ml+P/vlANuQvAXccMX3gcBLb/6jsAt2dBIEqXpQYdrm+EzNUFWgWdvArNC9gDl1DcpIeYpWev
xEywNc4kwOek3D9Br4qO550t+/qYEVbX0tSlD+pQlNGK8KQfF4GWSazRL9yEgxYrfvXsLny+X+La
bT9sqazCt/TSj3L0NEcvXi7ntgv1mKuc8MUHfyvWXpu/3ixF2d/N6IudEsYk4udcAUkkNjQypZfs
5ZLhN+8uOKamVCDC8GFPBzhXgbwQSYNl+xHXIgPeLasfgt0zE7pDWGVE2DmRk6dPUqjqm1fMJN3W
vYvF4J/xJljUQnnUAPhTSoUWVqCEQAKlp+GMPea60A6KhbHI8OjkYQl+S5RWAlIwNlr2l9rYHpVQ
PGhdh90m+X9kTLYxteY7AzFgD5Tl8sYlR8bAfI/yltdrqJIaeGKffRrrWrJCTP201iqjXFk2zkXD
tIk3vNeNmimMINRKz7AIdi6ddEEslfLaPDuAQVqMLF87z4g6+3U/0mgTzY9BO0WjVo2MF3b67HiE
VvToXtyaGkfQ+qNgVSkBrBJD306WAGp8bHhbHD1sgJmQjOhxcaETy/zoyYBujIohqvGzjnfo3Tvn
guNFOzMOFBIQRao10mZKn3vWAH5iIjavkDyP6eSMlOeLY2/Y67wKv+FRJprlo/K0tPjjGr4lRB/0
SXDvWVjMY4sxbe1VbszbUWNTwPVlySvhYD6C7ESrdfxy4eIs/2F1ZLTAZo2qnhOsbE2/EQlRXlt8
FBM9OCcGBvvlq5V2Nb5GteN8WnNLN/F4nAQ3bEtAY6fiuu6KR9PsPXHW0toD8RIdtHvUoMH+uVWu
XvxTf+sTOn7AaaYvYIjCGR9p9S0WD19azSRNXYL7dYCa2fMIgnbX+GGAsQZj5ii9cvBQ8JpTNS17
/iCvy0H1S1T63XhQQsTWnT9ruBJegnLXht9A5eyDJcau0dfTRWFPbqc///4GpWd9mDoIBMPcRX7+
RzyVOEnBccDiPwdXppuFaduSBR5oaTp8aqQbMub+gyjvjuRMVbmhFU48MuErc85d8p9Z+EneaZcQ
rGA4ifTQHJdPnDKhBaym4SMkHUa9YyoaUBEbCAbjU+S7SgKD/z+LPbwc6X7h9NgVFuePfChmW0r1
X1OMiCLgZRgQIQE8+KNOJwp1dd+OF3mr0X/pQxC4Xk/ucnoj9noUW0rlE0wl6rk7+A7R+KvtZd3Y
kdh0I4a9Tea18985KFTy/R0izniUt6eXKUUD1MpyDIofzXCKgx23p/CNVI/cOGr+HldJRLn/ajYY
aX5cgVlPLYgb2WENv77HRCVSGQ+iY9Hge2vfvb4yVpLCe+xmJa/gxdreG97aBgKwRltQDQedwFrH
2bDjc5ON8pLtUZZOQ+97UiF0W3MMmPkGn4B34VtKRsoENmTGadHKXrPv7/xvTCfvIsnp8AO/nQrl
nEzQutuG+FDJ695WqDh8rOVun/u66IfE9HgSkY07njmp+WCLz/uIN5BtBX2eAEvJRzGzadX3F8Ii
d5Y83EhGu276l3pY8umH5fWXtbvzILmFL3nYk2C7NYBhmyGE7TfMAVrhSbkoJTK/3ghmLklUeHuu
zuL+jdOlchJtzqxGZ+Maa7TVZquVKjKK8mFbPcSSjXBUaMFYTZTrp1wOrIQemDRUmFA5TwZEg7oF
HT7BdVAMyKDjrjJKYbIS98mYq5qdMGUsH1IA7ma2KF92UdXAh4thB6INfYeFEqLfDtBoeQmTTH2P
2EDD8DYrBuLXMopiCNKy8dXGiO+uMTDv6HLyD0bbh4G0fBYUR85ZG38dsvTcKV2dzfJVAto7Iwsy
udDPU2xfmflHn9qle2yRv01Y5xyGN7jdSG5Z2EqmfVlc1C70tXXs2yuIt4jAyvBqgJDvLwLfLOz4
lcETo9nEyHcdqUZzlWDf9wWt5vAlIYBwRvfvMODMmEyRpFlycrSPQ4G44CICz2lG8TOB6wrOI4j9
0dTNQi23pY+Y37N+YZc4y3a3Hrdc70U59k2eo/tAFIsrpKyP7570MVcW6nnnmhsBEtV4MN6c81yE
ocyMSXAAuXdTmkOXQ0S825dGi5cfmBT7rJjSLb2F8SX3aIRa8VE9n8qP4BwIxmJ9+hZOxdDndr2w
LoTYLSM3k8CJUWfuEX06YCN3GV/P0/vNdXRXBlvc2/Ytwo3RVo9KQi4PIuPM0KIQklNqostjasOG
WvQJFPiKAgrJJWS8tc1viQofehRIXFqPPm4GJKg9Q1a+lbO9VW3aD7stQRD+9VTVWnrPml6JXLCw
7hV2Ilg9ikT3UozfHexj0JyGZYHCNvZiGy5LF/uGcVExurCDRNeGtScV+0glYZZvnxvpoLyxQzri
ulbYjuvJ706P7EO4ttHM6Kc7fIWQSOOzX2qyltYP7sJhjNHHDtFtIEnWG3dEnlQci8QuyoYVmbOD
UQnhRK6dfMigWJnSYA993/81avzc7u61PUB6nY9lqbZ0liURW9KMbrTaWz8KYb43vlkpSy5odZK1
IqC1gMd6VHuyq8nYlVcuBJK8ctSSGEvTNfLRvlIyswBWAg2OlZzGeLiUA8lrKqnt6n6ITbUWHBgd
7SRfjgk8uabnwNTHMouLkmLJQ/MfhcYao9hUloHQ5PYIZ4fEo9zJ8aAt2t3hKWrl3V/eUtTjxziF
TT8ufAYz7QR3C02w43J96tnLWwkiZb5/5EUe5xlvfAmW6R1yNSnjMAvaLjHvsO7EZAjkSMSSkLsr
xuRrPx/+KxWt8usmEOU/XsoVnDdGsIEpo95o5a/9Ns2FqgoJVmhEyRk8ecAZ5CBEvcOCRoPfUlJM
DkFmz4oS5oalE5Ejn6eEDUsEvqbEOQjvCTNViepwUIlY+ezoHxYBxd5K9t349x6Bex9eawyhTh1A
lIpp4H6JOxZqJFrIIfNJj67KOhifuhvrLlvFZEESTJQKHK/bMvCtQQQrrGye0pQe4xEsYFf5kWUc
MauDzAVJEcC/ajE867yJMh7vVIRfykm89Nhpmh6l4nmO8v6U8qbrAlQBdb2XJbHDGWqBFB2TCZcb
DL267euVKeFMAJIRTesNtFD3xtY9tnWjH/Rm7KU+0vnvyQytPyyt/H9aIBPAWpEIveITTV320Bee
/YJr/VtSTD057XkBCpJFhMc0A5RaAjgsYfpQHecZdugSExAG3mu3Lt8O2fDbfCC9yLfschvM4QQW
El3apC7fSfV6oKQF+4SyKTQBalpCrEtzYXcI8t2e9tt2G81yXUC9uVgW0W/6SgeFVBEMvuSUkWOx
DzwiNVWhh0hFS+YMSrc2UZ2IxpOrZJ6KLtPybkNADYq/k3vFD6iGjoK/LpD4Wps2XjjtfjBBCmwt
TTq2dAS6tp5hBarmsrVUQR+aQqER1oL6D6pt79iyK5KEiWJSEGa3/H6Z4WKGklZbmVUbsBuFKgDS
l5NdVHFF05PmzRJRQ4A6K6cZhdPLXKo577jBxhQaH2X5YC899Hx8HTR2s7+qVDaJcOWI8eQVDlf5
/gqj4WZk0VlIqquZtwKAxgucDU5d+oUmhUwu/yvhbRYPsJbC76ka/EKLWwM6DMn0WIFvRu+vwaOb
SgAhWOIm+3mzDgc0H4WzfE7FKXho3PRT3BSHWq6jU2gi61wjoZ/pRbtojGmtH1ssBxQ1+6wX9ap3
IUNRyITri4UftHWl9bqKXq/n1rmFSMVz0+UiBb952pTVcgIpXTFedd4Y4R0TPB37p+sMWc6TZu9E
22Atlh6faRj3H4sJHGUEATBwmG7mwv6YMUwm/LMF392jVvunMCJ8LNgSSRG1DUSYB/3l2hRrAqO5
s/j3Y4bzKcLNmB/rkZ1sT/yUHu4O+AmTgpJfdLn+NJQbVBqycVbO+T8ZCeCDDFjhk0LdG0niBLKI
3iTrSnAVrAHROLoxpwe1BB/FakbnXik+sGLy1FDUiUwNtSLsXbI8WbFF2ImaWdNyVAOdBa3/6M7U
5UwihcUK6HR6f9rMCIbKEMDSrL0M+zEOi4gzzSGTlB770Tp9DButfuO1OmsuDeUAw3nGUDTbgrxv
uuJJthckaBwDNtv853G+Jh7vFRS6+cy6lGYqUuT7EsTEHNGhb+sEjQo8BI8CQ+DIwwFaOkfRft05
Xrb9jyJTxRX8wbPNTHJQ/L6V4ZJkabveWMYr7/vZRUDfu6s8X630sM76Id2jtaroiRxje2gtO8Gy
KtxY4RX83Um7zmJ6vcqMAb757xRvfVfmVof7k2tSqetpahtWAZAOLJyeR/wmNyv9O8D7ecNQ7ERV
p0Dn66AAv7j+ylPgN71JRNlqAjuM98Xw2NP90f45Jxx5jw5UALWs/amGI7eQmgvXE/zHZtlRn6+Z
YTAf6Lm6reVE/HWpJ3/Pi+JU+cretFq9shHqNHiHYyKPdV5JBF3n01hcS55Cu73bF8/qZGlLZand
YFNHwkfCvVC5s6M87UCAuzi5kcs/BJVWFYaQi9bnlSl1ydJW6iZYAQIVtz4yJ4WwCsHkbBLKrlyI
bbmTUwifmMblKRoVaiQ7s7EFyOLMP9wu30oodRAb9+d9CGNvd8D8CpIa+sckkTOLFY4w+ZwIrRb/
4heDrJTzn6iuKwB6EUxZzB3qEm9D5whg3gQYESt6p7v0Jai1bJCg5/r+ea+MU6X8td2HcCK49fOq
q6GcNH56tEfbzp5EjbKXeAUtEX+dX0CL7VrP2iDsmhSdhBvoVXhHcLqwFi9qO6tG1W7szqLuErOW
uzLM8/2KzO/lbf3HPJh+/+mfF1cxIbWR1YiL+D1GFdjYkIzN281/cNT0BAgoOESCa8TbR21L/l6Y
IK1RStSWJ6LyEmxDuGP54rBcgnbjd05CkWjO/RRg6JIhuQOsAusqmFbC9kST/XFgY1XIIawLYBgb
bXzmtkOPVX0QdyFy7wfm0/+gLYH/9nxEZN9TLFSp3tpXSYxwLuecguOh2diyeUnUjyWtLXs9iX6E
4fakzWrKQiZWt386cwNL2bzd4Xn0nE4CaablGZhwcJc76OO8POdr7ZLscoPw9u09982gI0mX83AL
YJmWZ5SNMy0L110F2ZAz3AsDvPkeC+YmJCVqpXxGfmKaayc1Hj/c4a868eT43WSA1Z2fjsA8+yr+
8I/UMMaD7Og7Um76ewu7lf0PdfOgoHDSV2uSLpuHXR/VlrFmuViBCx088RnQRq0n+Bn5+bZjXhYt
OGjWLj7Y2O0wYKN2X+ivCfxqs3BdkWfi9QY7AUXHyW3MK7VW6mXr1LQw3TitaMyrVv1QUAUg41S3
bjTMoKuUtP1O8m9dblnEAFbOTBszOjr12rJ/R2UmKdOZYWno6VIPyIAfANrLidj1Of7ig2Djig73
nCXhchbBQCEaIjQod+n379S2UcxNQRECoPBqxT/XUufMTAbHLtIyX43e/imT0Nf4Njs/LcwxisOb
0zetto1hPZGsGlpzFXkGjE9p5VEsCeRp3Ak0DXdjZWMTLce6xhGUIKGQ+ndxgmYF3JZ+oJtTPpoD
9hdMK6dGctnFaqy8w0r5u3JJqVhRsinSaYGkLQ5aReQ18vPJLpqTZMh5DU7J5dKvdJ19kZlkIR3s
oHlYdwd7LjJQ2qTicLjdQrZZUYznhe2FYuQ68hCiAp8R+AM5La0yqDIrkOqEPgcbfW7zX5nvlulS
pGkeSBjipTpPC5+QpuZHTfKyLS/R0VWUK0U7XI1yXVCqWjWEhgxDzfBTjhMfG+IiM/nBUZcWivWm
Za71AdJK85HopYGO37XQgxVhCLWwvirZWkHThjkVxwSyGa5aHjQm1wO5cf7ww6MN72cLWgAWsHnm
aNDF1wwtFtyEuTBgUTmouqA1PmJjWp4+vA540r67fjYSjMbynN0JyCh+q6BrgV2eBJ0vqk6YB7vn
jWjxwjaSshhK4qCFpAUBmX9bK9SGvLVuOlXNeCEi99P6eef0NN24jVX2DZod3aYfE65eZ+Oj72iL
CbhiEnGTlC2DPWwSGnlD2wQYlvCvgTGRbrtw+kayUX/hr675aGiU/xrbHw5KcYA+ZW9HurFaVFEn
eOsJSpvJfQDfTP7N0APCZbusk/L0wvWU6fHWdLxvJKXwoGlDE0l5OD0c5MjtKrhfGfhkcbvU07yK
NmF15Rg00KeIHHpU1Dfx7r9YNXWSOYoFRBOpRBXwId2CFlftZojT75Kgp+UEE9KndfxbHKFOUe6a
LFUVjOm2CUefWucxUpGH20DXMJRv38JAmkKdFQ4cvlTc1eJYmZgRFbO9a3qsQyR3ZUuAFLOKuXE3
u3yiIyVJ52bNAiMiFK3W+CQFwhCM8aGMenoeD3cCu4RgH7KpvxeFB5hzCXvZcaY7pkOkDlEy+7e6
CtlJ/WkXNlQ5iMx1fet+ZSZgq3PZqBIGkCU20aFPEoAmBwEvv+z0dUEgXhJdhFpCjK/nIF9yjBe/
y7aRxPlvOjQERF/w5PIbXb86OO/hO8lctHzK6Uxs4c1XUTfvu/dpNFrun9JMKa3CxScTITR95x1M
C0dOHOgMBbs7OmAzJjPAstkS22KY9eygTiOovMJGKf8oPiMOvLjVYPFm49P/XFDNKuBX7d4u90nQ
IpQz0cTto0njWtz8SkFHTisBaXX1GF+DdWwPBG08E8QPtCUw4Al1c6kQEfg7/tSBGXUQCiWxGsLt
wNNvcBsNm7og42/JpJe5XWpqMI1pCNSj6CwqjcxamLzNxBTCPBzZ8AAQXMCpsSBM5tu1z2BAsr9G
fm007G56ncq5KK/f7tvQlkxXTJEc4SNzZFi+alObLaaLfTjyhXOQzMO4T1m7TdGc9ttm5WfTRZBY
qwft9Dk2UP7t5ij2N1EVyrZWCdfJHVdci1zsKtyHBO7AXBckK38+0i06zVQwzUlig6oWYeHeqq51
9Itk3lNllh4c/tZ6VibroaAGBsD9S2FdDqNyAKZXVITZ07GQN6bEEHwqzTn21whE7FG3fWKWcOoO
4DDS6cAZwhAn2yrVj1fTLYdrjMEdHPVmZVuoEIwH7ioUSONuYm2gBnbyzhUuNw0vO8pIGa6m1XsR
TOlU/VRBWqX57r2WRS0UntVDctkNi+CAUsoKd8jiPJ5zlA+3hJKUesO/6LBgio+EbTo7NCJjCldy
3ABkXGRzgrKGF1Myw8U00o2/ceiOHU17x+czM2kFNtyDU18Dhef56NvHC1jCDLKViG2s4Fv1Vi2H
jukTROY2V4IzecTgRuVAPnbD0ErOdGfAWqklFDTzckXlbo9wTCPDhKUsvujagIlwYYNqKPpsgc8X
ex6IG8H8W83Fs8tT77dKsSa9LV5/NzTBinJIHyoQSbD9Pf1oTonFki+VGCX+voPwpPwWqQgeShKR
RxlQWROvVQ0WKGS2oZXjTJfAvqdriOJ0/iKPSzSzM8eS2SnR9tcZh4rEVU9x13LfaETVVcAosRgd
Fm5h1eWt/SOeobfGR9fiIa+SAK0T3BCQp20nItzvYsI0c3m+FfaDUMqSgx4vUAjsGMNewNhP3aMH
oCiUWuClCVcGMCBfIoepXrvFLvIuNg3wP4E8jhtkhDyLp5JL8sMICkpC9bg4IGp9nxp5utcs/CXB
A/pNXml2LWr5o6OFRgTNc0GtO7VMZiQPNpgEBL6C9f8SkuWfhCGMjvfTQ55xnCoA//qgN9i3LnfJ
Bz//ALH/lfDQd0fJbgAGNcTv+FZnubpg13MX/QXG4V6WFkSDfiVIDIiUYTcm2gBqbju6nrtmj0p/
nmecNL4F7gA7bxYT2JhF8M8XJVWBVTDyzhfXlMyOZmVZBPZM2fDGsRO/5JtE5eovEo0G4vHTkgX0
6bY8H4SADnnBbTjcKUSV4J1sT2aktjWdBXpZCoQgEW0hDyZpdqFPR44AaDvCuxKBOG0gwzLCMJqU
SEXe3zF2AYAPNNgj3Im+18M3wSO1J1xv8JL/A1BBRBRWraAGIuDiSRO14zTMK4aED1dkRVGwa5+w
t9hPUCEGAxwhl9nFSiHvBAQDiQW7A/zamWjr+1e/4GmSwTqgcZNEyov/S9oK8uHA1Q6SpE4PdFIa
RluV3NX0DzbOMKr+Aq+2CnoMvgHKLuYV+r2dOJ3MaH06WwFTaAd1hDplwfL9QX1DCvrdRph7EMCw
lEmJFVoYbLD3TbmH93T2E92TABBxJMgkIWdXK1A0O5GHbHI9QqZL6PwjkLfTq/+TrSndrE6+/p6r
2kFHTOcWNnQOb7Af9wYC9hJkqATsAl+8ECfDoq0IxvmrGrpmiNmMynLIozAmdybfWx4jopqdrT3h
TRgXYa8d1uHfJoQV8UOAwI8E1caAnTHzZpiZOyAppMEapQ0DuQW/UNi0+g99eUVWRZNOpzXNAoST
rzhAEICC0tI1AnRBZBMfbXC8X70UJ1ZH5+uug7wvyP4MEb2oL9WzdJEnoUTQwHPA+i9+uPixGPXJ
3mH3gjK8yhUw90I9ONT4adePlC/ewlVFfsRmo7ze9uS92l3/brY2rVHdzeBjXMCzgPs0ws33Ipbq
kjlY2iPahlzJr+ZNqZ9GkrRt3KDGGz7Fp1xPYpOzmxO9v+CogW0xsGRQo8W6Y59FbC403Df5tyAg
Kz3LaCjiYx64gOSLmnXG7F16cQ47lEEDE0q10Rvk2k4f071iYo+d3C9EYUNDKZkQZlEGisw3SNwF
RdgK1Lrt6sGUNZxG1a1LySHoH3PG1k693xST1kXqzvU1LRoP2h/TV11mWjYD8OMQMWdXRd0VEAUP
jxRdOt6KTgF+aou2Cl7PlCuJtXxwIXF/jfFKBLpc/oihsr9IlDNN/ssE+ahUdVCZsDBOLPYn6QU2
J+kSicxan02gr2PpMU1FUEsA+xjtSgL4y+vv6+IpRZZ5VxbpmQToiP86przCHsZpl54dloM5S40P
4HGHrxTpW8BrhdZWDA4312SmEdLpRbPoHojL+lmLispT5SipKtmHKelYpsK8IniEoyeOlXgizA9w
gpJYH4PkBkh+pnMNTZAjEa4/XfSp6Zs0aBrVtkppisZ++u1JcO96TMPCoWPaBDp5l+sfIiDBYz6X
7teLlIfoT6rYfkgZuSHzkNvQchGK9730AKwXtmNfoRPFMXl2XkkujOH/2rcrEx4KsaPcbkzAkoLC
aikdo4thoxDIOvvogcoyFfHUCo1tuPAhqwC/5DXpB6D0R7+gidd4Wj4BCVLN0A1Zr+yxO5KaiLDt
qRtBbaEYU7dmLgDy6CvPBJ7gumXFrzaL/RxduqZObnV/NQy8PzBIEtTzfKUKIPjlTPo8fLT3r6a1
HLbWmSl+j1OpsKzjgEOAoAlZ4a2rG7X8KNYy6soeaO/V5gyNboFX4Zjjtrh0PvlqffI1VSe6/Oba
hNnSC2QOSyasDV08u3a2DIm68HooeWEWF9MFI2Ilxya3TszdQ9Q/8vltiWlnncudLGpuFVVrL+n7
Q/l7wo+ExlhWhSl6WgW37QFFhQ3bJyqE29mPxV86xkBx1z+JoJLT+MQ403TQ+oFHAxosfcr+r49I
i3/7y+GPvw/I1eu8aYoYBmBf7+yJUmClF0y41utD1/IgkKNrsKUTtDEtkj6iqAYw2MWU639D4kks
cCEeT8CQqJVMZd72jaJ/0FfIRmflqvd7tA+k1KbgcvpFFwTzX8hfNiCI+t1yA06WbWiX8TSGsM2m
Lim5BID+hpC5KFc8K0xVX1lrtTGXzIJRGlh06bFUamujUbiz/9bA20B8m5XAuoTA0jm7RKZY7GO4
N1MKo7RMw1xmpkcFh5NQ7apcGBT8glosR3A1BBWLGDneAY52uxpRw/5W6BnQBxqQUBLevGjJkFW8
KUbZBq+/KBRbTz7IrH9U08X9UNJOM06P9Sx2Ip3UKO+EMDn7Igd39TbANjTGUiI4zo1pT4NAH6zn
906Y5W3Wt2suUOmddZGsR47Bc7JchUY6ClIJ0tB059E+5XSvZSPIJPHxqGDhpoBveSWaG6Nf3nUK
BmXi1sS9AweHCAXIPoRf15tl3ATb2OMZE8i1AkM1xOvfjsSofQdCXdBXxrUlUAWTotT0aFGYVcHR
wYUNtsd6QuRbdb54EAAuVuqLac8/T5WdXHRyXsUOUqYqdR0+fdXbepslGUZS8AFamQSUVsdSNzJd
uXU5DuVTY0ktONuCNx+BZsKZHWap3gYYcrBmfM09megkwkCrGHsqs014TERzPCPuOsMKq+Lyp8Qm
uZDM4AHRRX7x/PDolwjjSxKaeqrNtXV5PG55ka9XiiMtyNR3dowh4h2TaOise8I1caXGgQEJ/BMp
JBFL+C2M4YbwW5f3o30ruyc+1c2OtjjMjg9Z3dH5fe43gOWvghhsaU06gkX4S9wpN/pKoagb5VUl
TYHUKr8SbpScTjuMByaOgY8Cywkr+W9h0fwn70Bj2LSuNJaf36nQktfZPENAn4D8KAzM6FE9tty1
q4sjuYfNqQsEJDMoTnGNKv7n2ff1BJFPcIwDlUrqUPElF4C8+bKlvUJ2r220KKz0Ha8FbZw9Ze1K
A9p0XvvFtCdMZlM6DcqFqujRGMkwCqv5B6ho9UVhfaaz/Oxk6sWh/KMheqyFYd2Oq/MV0jmod5Ik
bnHFTHZah2GsSK+KrOWDP0kmoHhfI0PfC8yJvKt1nhlorVJqtOFy0RDFgtY8ISEfDjwNkis1QnbW
o87SuKMGCnpuaxzXRc8Bn2vRlhex7NLpUfVSMRwQRQyulfLLpokrskqV4PCNlqcz+n+m6+iSaeEa
ziR7AKJ0XBQGL2DJie/gTSS1z65wrTjDVAZFGShgZ5Xl5HC5oFGCq9dSRbfStbPL6U3kXzPvLcfM
ynkli0xeV76yGURznrR3L1TjjARsvXUnuC+sT2CQ5JfjxahvgufF3cWf8bfepS3O/2Z6Uq6HEY8J
47qbIq3blLMlEn2qdMdcq4HkcqexkSFilbxfCYZrJYFSJbVRkDC+cnARZ9RQIM0VAM3gBxI/R9xb
HjqcUo/w9aXEI7WWu+Xzo6Kzg/RgH0VuHDf2ihXZjV5G9sZe3X0vAt66yDA2aTSeND9eJ0oULqPH
S2Eyd0TiLkw9y8oC7/1OBtnbaN5CdvLHTJ/IHUNFU6NNZ6xALFMoBfDP515bWW+tXF5SalYljJfq
StOgOmrMFBXbhWSoUXJvUZBVZAFQuetg85h3LQkMVgb9ScU6fUTBhOj2l3hPAM3STUBRJg+cVPz6
G9/cb9+1qFi+edL+WOLiooZzBOrWW7qHZAuUP2QuTKaARRBTOqF5U8UhGWi1KaIgPYt7sflyBZ6f
R6yT810xt7XqmCq4nNMYKDTqGAw/NgHOQ8rc9TzwzmC07V/0HCaRMiBCE4uvOldNTw1NMPAjp0Qd
sURjtVp9vdthQcZJI0ihhBEwJICtlYEqsxD0vbFUTCtlq6Xwykax/gc2QBOWuYQY2Cg/VZHFo2wN
BDXgIIy3avjx0KAXsH+r+v66TDs1Ul0XXlNj+jE+Qegjjx27fShsusv0UJmexXZvAGF4SpRudw0K
TH+eG+I5Ri68PUuFByp/ols7fMhe17KKisCTCUApfqUceVoGDbdEoA6TeRNf1TCnEhrhkIinR5Sg
h0234qNo5KVUrQcqaQHtM8YDPQS/i1R93SDRJxQFdX6ZQqTIk1CIsP7TWIruNfDB4lSBYJLfEhPz
n/pWZ3a5uzM1I4gXxQZnMnRh7fUaBNoJSmiUtzFpPhrCtZTZcjMTZFPOXAA427BM8Js8/RvxnOxT
FQLdROq8vNw0vG3SwLhQOvFeDqkG58QMMulLqQdbBu6oZxoeZDo1ebpOQ4GfOXnIzG480Jnv8lf5
+/CJti2SwEhbrgeTAVbhhoH4MNoYtWT/h/rHiIZ+xBRS23x6ZJDci+oB5w6/p1VDHUV9LJTTouxU
UcyASDolgN6hCwRvhMUp3ZtJsE8TmTjVlwSMpmZPtfBQjtCI/AxSKIlqN1+KTBgI2WD6PekAmDVm
N8TdhX2+sELsT59Rdx24CdBhLBuSFexM6sMU8pPHU7eThaAq8dJhmeYHbT8efohdhMCcoedRBOh2
ksvnYTFtUQETwfcKluIzzf2hIa8/Cn8SYOBjL2FDh5pyNINGjCnwKic9bAssp9JjXRcmRNwzBpdh
40xCQdUwadFpcyFNolrvfOZwF65wj6ggq3s9gPoxvE5KEUeq2kUMbL+RL2QwuHy8/mqWV3oWkGqF
ISbPmVnPq+4d4gLX1c3Pnej4HL9+bf53xYS+UHDSeaBzOINHM/qtl052jhQOmDNveikCWj9T3l2O
sZCW0N01CMgGqev1TfQxTjD9+1Bo08j3gZTvY3kjDnVE0KNmOjhb95wp9EVvDOXvN5d6RmMQ57pu
pshvptbwGmtUpjWUiEYGvKNUnfZPq3TGLcTUAdbn57gDjjfD/ztvBVJn5RaXOwJql7iw6jQHf4eI
Qy7mG2v2+aRZ35FjyfuJ8/uDxRFg8oOJGZXIFv9IkJsogFhC7JKWQIe2aDEPJ4aCWXoB0dW41IN6
mPYBFUyUus3kqX7oqevPaNlnOuFeiQ52kE2Rfro+swSVWvw+tdMw38U8yqegMdBC3HbVbNjkgWtr
uw1SV5wRQ6kdwX1ICaD++jU2/wNQyXhz2dpFoxNH87aitFzjjDrD4woe6LUSxEjDLN3jrOY+3NUJ
ZIxUq/koU0t5eukYRFyP4m26A+Lo/CDh9emSfqKGF2DtxN4VkHcQXTwohsmyzdWM/vckHciofGjK
FzyqbmKpspa6l9lKS1AmMdCOU+Veg+BaXSmSkihigsqZzYvs9ChjJAqsTJ+KPuPeh+g0qy1deUcM
hR2PoD1YdMdsxDOGz8Eox6A/Abb+HtwJMJ+xCkErVAuNu570P4Lj5tieiQ2chJB7Leha/0kQxx2b
BzYH/EJeCx9vDbj2nxGvc7lslDGYw+YM6Hj5ypzWPuar7U8PPpBr7UGXaFl2WD1kIt2JWBSxeZkR
pDLvqCmksRM0bTtSHFOQcsJ534EgAKVvM+Vfz3DP2k3FHiP2t7O/tVVIeNIKImtNm3dDzeIc3Xqy
pIDibnFVmwZSn+kuaUKH0afup3F5ThASLIswp5VGb7pwYTTQ8SW4g6nPV9fM5a9bMZyRd89upLjJ
8FRwdZrWcRYUl4w6cUnR1OISPGfd5AAKsWSsITngPZWHK30WFLz9OMM+elPOA6bm7ci40AOuRm/3
U6qp/m+NJlNxYMgRBQSpJ+78IfIgbZd22OEcRU+agFIpLUPeCV+00Ve+bINtHbsbL7RLsSHtgG9i
wTxdRZJybPdbYydd6hzDdqMGfzewkLrH/BEnx2fwJF/79t11AzxSWy8MASvlgXytw+scC/ECwOGz
C/Pxox/urSGVcq8AkqNkfTgWJlgxloR5fgccGI5n7pfMIJ30NMMfxoyGpXQnDNO7Osp/RQwYWJgo
swhuqAvhQ2vP6FYCKpPsnDoPSLlz1ZO1zWApZhw2OTHi65TKBeWMPZnbOYq/kkBeftuQSAU33Lm5
z4kdNXCK56uEeNR4YOpXAzsNh6QSWWD4i39FGVoY5nMj4oDxWOLMic1AaxFH2I4MjfPiyQMParxc
M0TWMlX2mtpnKf2ZyN1PZxvSKtOb/1JCeKJ7AM0lhBUHSDK4ZzzGsjUmvYK9y0ub33clNreFsVUb
d7/k6wZrOkd22i3JrxckmiXrG3HM84rqE481ifuNoNDeJwAJTSWpQBYya+AQIXS3z12fXGPPkxzK
o/Lo40caj8JBxdjGao1D/z69GLLk8waUjsP5gCQK5L469JHeeJQIAA7genpr2cH5ZM2Frz5ToWQ5
fvWk3D8E5sgxrOgB8liSuKOBvj0sdS0bQtX1J11cKecaC42O8guyhFzxUPmNtZQHdVagK93NSos4
5K7zJJW20Ccs8A24Dx0h/oqwvV+WqjZJtf16+PAZ2IO6wfAxK9PM7tdYuTMlh6FDrFs6w+C+Bb6x
v9gCeukadyJgMwEKxYoXpfXxdYJ4DV8iEHHLWxkaLNQJA7MmaQWkGllucQyVSHoRaqFeiTLmFAnC
VB5yVmz3k8MDDZcwPP7oaRaoc8lMYMg01CzmlW17Eguce+5b4e1f+kxzjZsXgIO9R2xM/z861A5O
87pIcFqPQXqzBKX7LlvH6LG/wpdPFONbSsDepOwxY3/hnxQbsMy1RhJiEYQ24zyxUDQDkv/6bKfO
535JYTKMc7uz+nFdIRPYPiOUWkNUVLJoI5TNL36AvnQwRLkC5y45xYzu49ViyFzzd6vPj5HMQWaj
Krm0rQva9XkUqdY9ei7J/INadhtrzcxj4zUnB7W36/hW6lXGwmk1vF7ENsJQp4Vxy2hOjitur51e
odjB+gskvGwbw3hpaWad0n0D7b4WITlfbXtbT3TIDLH+E6HNqmV01EKLTu3hque459ltGm8geteQ
q7W4KwQZZPVBpzZoVpR4w9rapMn2daeodkd5qR697zisfcbD1yiNNpqDBe3G+fhuvcGGl0H8rAwu
3DfsDBgD3LudOr9HEbF2hlmHp2GTdEfHPLx2MhfFzgeEa5aO6IrI0v45XKkJaEA2KH48vNCYcbF8
YsSgiCI85X6EbOWJvHKpx9Hn8C9C49GF2p3d+A9gijY0uHgSDXLNOzxFbDTUY4U5EQqToq9syyeJ
6rwHOwI/AqVVd3pypjo7ZY4ZkTZhI5zEigH2czxtz9DySdRMcc3DOlloYOUWHQz38Gvj2df9HG8H
WSkqYp7qZw4kf2dZD2Krudi8OT0z3WkBPwlxI5liVAsPwkPBCF4mO+tVrHCzLL/I+CkVFdQvFBdO
NBhUIxefxT6gzCi0gvIZ9u+KpWu1v+LcJZIJWHJZr1b2e2ZagFC3bzW/qxUPqQwjO9YrgiGWiRLR
jJlUtpNga50qnb60NmEDnyAz/eNPVKAa99X643MK6AacbCqmHCc408hiY5Ypz5WAsL6rPQ0A3vxi
AOMre+s+qLwsRYusZBBxmutLGKrFjTkmQFBy+jpai1pK4X2lJDGXuXyEZygmhpw40ah60NQ4ys0u
EXwDxpUA5RQOAzI/876G+MmRBn06JEJJvMfuMo6Cj4DUTwrZ97pB6nXGYfYH1pdOqdhCbQz7JfBT
GALjQZe7QF+AM0lZXZSSXDImISfZurbi0zl5+Uq9xDXezj9tmJfbSp9kA0CeEErb/5HL3dhM8SAV
2LgDxDASQvqPJfND511ifuxaNRdOseqcijmFQkdBBPNAgxsqaGVQg88j7LB9xA4GAEmPULFVB7ng
VflK9uVhFkTnLhLJusflzLsl0vbMzMcUINRjMI0O3cF7QbI4myn33EPrpRyzLSZv+m2dduFm+BD2
k6EVXv0e5RKaEQmOzwO4k/xHFjPr7QGpKa7vpdSbLd5HRaCOCIo5EMQkHTc6r+S5yqNQIDy41Nqr
Yd54v9idOZnQY0NSzRBtxNuinzpIzA44LDo9SKR1BOc7+j6hrwG2b0kHEQhcqw+5xB0bEFgjZh2D
sC3xsuXD5d/blxe+BJg1NKY38xRNhqNhewVcGPz8nxjW7k8FnTgw36PFa3L1g/e3zKuLaC3VMQ1W
COsF4ONt7ASVyX1vJSE/MgYYppg9iBuXtebNQCj1GyvO2f4o6vO7zwQLVeNb2gHn6PRVIb2PEQI7
0sKYYlSoiMNqMVnMomlEVwOqLii9iscUJcHE+E8emyePfM2k73MsMN4mKXkBOXNnbosMSZ4GnpDy
JJmhWGUi26DzYOKQL8e9tAUEPB0QwGC71eetcbRBB0H2PBl52ls0M0Wlkgz4GnHbpDes5kBba9w5
N6grs5F79yEsVK4vbhtZsNY4XBTiu+BJjXsx3Wgc4BaW0zls6KFcZNW1GbWHo7jhLfh40IbSKlrt
Qqgn5Uw61gBK3yqpRUhgNrT1JxyIpQgZT9dZh/2j79MvyAMW1AAaDSpQX1CjPV5YtPNn+wbXlWq1
BjNOSexON23teKfS6j0QtrjuP+pudOPP/2eSP4ytdrEIQglkn1RW9CcOQuAoCCPFFZMKcJS3xcrV
JN4J7CENtkl0iEPAK4S8TcUHIOKZXhqS/CPY5dmw31yc7u79ESA+DNpDUBTUUZTHSU7V7Y7/4qWn
afLcllNX7Nt1K8PriniJqbm4KG/EsO5TQ5JWc4Ab22eGMXq5NVY0gCqhPfD0temNZHqQmK4saYqv
a8cfJSB9fEzBphuFXLQvKLgjb/zSCUQixt0VoeprCan028v7z0857b9JAWRQAU3LrCds3iSHXY4E
UOlqaBnQdCJL4zB4gHVeQbT33AY9Q0Lgwsk1YSskSEeEBBVMxpgPltRrtdfHOZ+nixIcJ7zhm8nu
HvY1ADqfZkT1pSmZnyT/r4TmxdYEsePuhPr7h/qri06iwQNkrPMkuFH5Y4eUo7vitxFsScvf7/7i
/C3p4gSG43GtKAgkVdszmMOkSJjZHrmA1vIpwKRhJB8kHRDpkT8on3IA3iDeKVgVQba//g0nruRL
/JBF6nxOMC6YOhVuji4baJxlvQiQFezcHVVxX4Ao+y5enNAp/RphleQvsl/WHbAJhfFoRjzXZ5ss
t29FxNqp361ciuxmFGlflmVoGDjIuOGeD5kVlOOAjygovVGKx55IYOK7ziP4lC3TmlBkfjboT6/O
Wivp5vT4NzyYtUUWEQcT+2upTEwPZ6o+gitZmzIOoyYxSmPDjizm2PQ4rt1n93EKAHfBUcS1Pe69
VSMgH6NjtLTcoyYsTWu7pBoh2YCiyjIPrF9E/Bnj2dbodmq9OvYQAZI303U2lbtLmumm+W3UO9CU
IYcRRySY4zO2RJXo94O9kqKY+jsnF8MBQp3yZ9GyhSG9NXjAdLkg7MnJR05tuZb+Z6Bi434dLCKt
gZU8l8GmJpcl/LdyEjH2bpqWtBJJ5VMSUlnimuk4IVOeBTNLUAH/2H/PY/3rB37VmcNkQx4A+3vf
tw0gvVn8T0A04dTn8U8jfUCrh3BZUrO5oaPYF/DZTbruaMNrnOW9G8ZWzxEtBJPVghWgMEzvyeHi
HzbPWUXsU6980U5L5Jt8/6i2RGf3VqOV3W9lPTWfANTsON2qclqbsO3ANDxy+2J42P1l4yO+vs3v
WIfnnQ40slhBippX8gMTiILauedZDQ9EoA9OyxJwA2MTrr3nsmdqRIez/tU85cY4TvX+n0vJFeby
Oz6s+5xhJl0GK5WoO0dGC3RI96rMAHmtAHFq0NwYpnEeAR99bwM3JNg5k4uM76PTKLmLe8qHzOfY
ciKrMyNbdh0IcEpk4HT32tJ4oX2tEIlcHnnKakr/TtvlJefV6AZkakatthzM1Nk+7sDUOgYlFfkk
8nO2hLxZ/A8xhQy4+n29DzwuTHTvimeM2Bpqz3NxcSjJY07Jo2RjJm6dpdK7+0BbSAdNicKvbOc8
M8l/KCBcRF6YUVk53Z417x1avvLAwxjM6/sYtBoX3htBbWssg/iueMNTAU+6h9iryo5ko99oTN6G
9zjQdDW4hRIUVr5SurLm4kuujpAGZRFv0+Gb1n8gq10Edi+wEwfRSeWl8Itzx/jNuUTIC16aydVf
CCmRgQR9wMEaFJ4hHC4c3sUqV7TxzasSDUmTeq5mbbi/YyO43nwyEi8qL108hLIdvA8vdKtpsDjM
XKlT49vwB2dLNsXy3enrvRguBsottV1nn7wZWPTPhO4Yj+3h8vXXNv0K7Z2A/0a8qtNJERgKoG9a
UzAz/6sSOJojTC6AB91bw3o4l6qkxSfJxD7v/wVaOoJcCveohBOUWbqS5uGDK9/365KI2rlE51ZW
MGBbrskbk5/sZBmfPSUr6Y3dQCxP66U0irk044wVuOHURx0+Or9P+eO/lZ02p/FD+IIuOeU9m3sS
RSbiQo82SA/J2lNQvtdyPz97Gxm8dsxwEKOeXUMThXbzXAXfo57NATn5eEv7kiZD91N3PTC0E6ld
OxxdaYl0NC25lUqTZQwGWTtylPDk2PwG6dRwRbcowt9F5nAYTnd2PzCdGUelCkGLK4CVn5WD0Yd2
2tXsTU6/beuBFYf9M8c5R6lkINlJYyBkvSJXCOoeEQVxJULpCcd6EKdNoO0VVPk3hUEQUrAYtrge
om/m+W5++SXafRVc4uZbOK18nol9L1AHhW+Ld49PRJ5GNqW8ReW/88anSmSXOoKNWfb8YyqUV3PW
+mvco2LpRHzxkVQJo1hZ/NtJd1/eia5L+CzVxLjIt+w4F5bNgJwcFn1i6ryl1xBjeFSSgC1aD6vz
3Hd24MP/759TLSApE/xaSuhLtWCrVIrN9LXMFt6HNkRbBaW4avqMgJZYxunLTIdyvMv+c3H1hzEX
MCXzRuA80Go21SwDFxac3EC5V4YONFShNxV7uP/U+gDkFvs7Bcrqnxy1usEG1URjK/e1l915/P7h
/acMNHA5mt4QkgALYNq0IHP1aQsKeyzDr8QEvfNGunr5vnMlHAvKmjwvIlUkw7RsyBlSs2k+L+2G
8JiwYveazr5dupFviK3omugrG9BKsZrad8ZUVwzznJuKLxsb15JHboGETHBec2oHlY3wHDJ0kdru
kb4ibmjGzAobvHPxpp8hWOR7OllF4kdvwNO2mak9Xe0GrbEWMn2mlPhXRM5mVUwlHTjyIfidw1eD
zc6Ju13ooDIcWHIqRG8uJvNQP86NW3qdskVpsOojqLbbk5rpzuOEnlfwRo0Stjelavf2JYyypAAU
RTqvCA7hJfkxkL5+c1diUsueUNpmQI6hHo2xKVCKzT1eC/kafrgbvAsLYHZrldKrK3xIrNl/LHbc
9GlEkirgd/PfjFmyoq52xtDaNgNte/P0JybIuHYrf3sriq7GrTpyYw6lBQ6adoa+34IUQ/S7jfi/
HPUCznmhXjCPq5s6v70QdneolCCCosrt2abjc28PoQZVyxxGgI6KYrL+Y71tLk0WiiJkXZRlXKgZ
ulQsO58Vb5OP5aZPtU/gRxjADqjFsEya2SSIY4bCHsUV2lMytWL1d5VQf2WEbagquguPr7lmWdJi
j0khV7Mv3Jau+m0rwaz7g7sqP1k92ixK2DwtwbWonkoYtlE82eN/xlN/ngnjtVndVTOzuHlJxpjE
tRvTQObdMgnkQ9JBrn98EqHUDMB1MGblJtu3n0faaqfBhIOrl2Z0nENnj1zj0iWjErJtDuzGBllJ
a2X9y0jUek9sPNE1gWielHt+SovL1i+lvsevGMq/eFvXMlKmPBlaBZeZFtavHM/EfKapLQmhCsHi
lQG8kZxUG2hFh2YEZOKD18gYLVJlmu9+i9jG8L3B6cAYIEfrWqJHJi9i7WLMM/nEP8MbeBOULJsE
GxJc6/27I9Bi6AKtBjrFGE6v8brUkd0bK4T2BwZjhHbRhmriOuG5ImX6lgWX+2ovVe08UvXdBtLa
fulboqDwaJXuvxAkxYdY4WaXTRzw4tZPqj6lixLZ1Mh5NED29xtGHbetW8NrpLp2Myp6u0QDJTel
omXAzvhBBJRkJLaTUL9N9uN/eMRTmxl1P8Mvp7n86TSVX9NDbIJkM3yWNbwr8JnkPr36r7A0h3v5
FGuHpYEHWcfrRN9bX+mToZ+mVJutLM981d5MUMqdYXy9fXDqZmO8M1/OnkZ8Ck/whdsEvQMTIeL1
kQVo5vvPV+xuwmlE1jNkgi/di/GB86e0dCR5LmXyQSHhE6ZiST+dwN0GBv4KwG2gZP1GzNynDUKP
6YR9U6qn5ZZxXBG4f6LR/VbwT6inXBLxgKY3PljB1l1F2QXFzr2IH1W4imhPWb6eNwmlpGTEWeh/
5ZVnZuULIwbTPjPoi7+8ujB4epvG9yhLrAPZ1cZ8nXZ3sluJIfDwhkheP9VIPqZ9pH3b6dBSl2D1
LsbbYSlXaxedhkNTQpv67ZFQP3EJ6IzUEQcHmhLyD44wOgRVI9m7ONBipCaOtt/mB02sUoPJI3rN
FJMMoHrDKMLPCLJG4YX++/1H/SsRynsASwuUifrCsJ7Q6QYtEleoEsu6M3i7FSZFZ5JNwNY9u/US
CsOgcNHyDJMMMK5QYONEbGlUK9St2bYraTZ0RPjBjiZpuTlGVG4DC2ruqt1Cn/H6ewsHuvwoll4p
6FPcdYBIbGkAfJq3rLgqPbDpznoT3CYMJwGJGEnwc+gzeGw/qAj8eYw9u/GrbMEMC3T/5ig3Fsby
RgI5kho0fF+WeuhsHbJNo7NhOPCS9grzdy1AqPAuNZ8SFAD8MQjABFZOyEy3RWZeovANZfncIzB7
IINm0O4a0syha7hZpA4XXwHzTAH0h36G+kR2tFY42UWloVXSt6cQsL2dk6t2eYvyky3pGw4QT7Nt
SpGMt1ixy7LAlM4FFoApguLnMBgU/IqvM1BopQXGj/GHOiJ2bgZGxbvHhIBBAnDhRBb+A41vBoeS
ZdF8bn9jmpmzxZAUjvunBuv3/JwkJGiWGJPoNy8kcBDIH2ryxJ4ZA00yvzHcqx320iuydIIOtP4f
Oeb9nVXEX76xB4jaorA3OpaLnVXy/0ytDVicmsKvFpgIO+iBdsOTS7cnfcxjZhuKRf9r3+0L0BOt
T2TjFOdpzDEPUswRmR6nEfPknOt5AtzegUd1V7h4JK/NGYZPFQiLrTEVK7XpRq0usL6fUCMXlr5S
jFhfjH+roJWvJGkJrC0Pviu+fv2HZS5bB/u7ahZACdfSwi2z8ep5Uyd25kAGoIPT7C2DgTDC1jhK
Wkq7R8Pvw68/LOPfctNyVf8u64UXBOGpIB9sFTv2xs7GE5vPJYValt1fX6WjXhB62HcrxPU6Ym1w
E7PftwNRWc5GRWo+mAKgZGb+1k9YHkNtkMtkKz7WYgsTLEIDKUStd7xNJNcF1d9ruEsmF+yb13ar
IE82KacACVk+f9Q4Nd9+Tbz3FgmA+PIsArRExPCCzs+C42ciBVp05iZXR9twzaNmVJ0o+gFGWMiO
Mmi3DJ5yJ4kqcmP4MkWXXX5xLeRH0tyNKxudZ4xvw6z7ESCkY4v0wL1kTJ4PcFm2oS9ZtfrYqH7p
HTeawx26Ii352+1gvp3zzP0prwvXrtdPlX/lIdEg11B5or6C3sSPmxRRpHLx91cm4BRhMus9zRWk
TOn471LWfbFWCfUJO3voyVgPjwKXws5lM9U0mkHy4VYEIgssyq7//YIK6CfzRXB8H3loW45h/VLq
RJ+Qy7OGKZNB4nh0NeHO1aruv345U+eDhGEm0p7Oqn6Aiofqe1PdrrSKXMPujbhgqnGgGiUNcdhj
hQKeXYkQvlLQFW99k2T5VRuz6uDCkhBWTL3lp49IprW1emLYNiPF4SMu0U/TywBhjumsM6xpMf1c
waEqdI6d5cRooryNKoWF1rh3MesKeJkoM2/7P1DhpglxFXnncMjU17HgzZFdABy4tY/LG4Ufzq3F
+hrG+TuOIPt2DCSEwq298tZfwEn2r+SBxE38YLkBtdMCgGmV7/ESOQaFaIXHHML/uCyLAFf7sdmC
wv8P3+Lp5uZVptpF9t7cDjAu4wpeSdet28P3rEHvdValZb+iDCW/zEqBNn01OWlDYzBB5vA+Fzgd
JmmpUifpYGnCQoPcHfA/JBoFiqRxZ10uU3FYh5OS+X0nXjOzShZ2YAAOD55ATEeNC1M+hFz/MMmV
Sy0WcGhICfUSumxCpkaVJBuVeUQR0Q66jedAp4GR9SLGJw3kKW6wXZyhP4Y5N3JRC+QgilvgRIqR
0AA81m1lRVpbsqI7Wa3dxXi4LidPL9QrmLrzhmuvTuITuZD8sezTsit+by+3bvrpblEApjz5ndpH
lSHIcLNLUHNlHta4CP5J59wLBkH+TosWu3GFmum9X+8VUEcH3jfN9W8ohH9FH4/G69pr9THcGmB6
wuxMRhVk/RQZWcoP8NTMts3wuvzjtB9wVkBfVbigyDqvpfC0fkTusZT0TGwDx/mzXhWyIa9co534
K/oat2ufY9wGNFJ4MlzdKqsVi0kvCeO+IpUwhR5S9u4EQpMaI/QZ2MuAb47gyCeMQDF9jTpkQhjp
H2fjbL5yYkxu+2gL3HrJNOBdW9/84byLPunWh//rGL9JMt+wcwrD/xk36OdIykWphT7uFSC90qs4
QmxHOSJuawVpP3xPTipHgmZwHZlZl5ObzJPJX/LEL36zKZ0Hc4YaWyYLNz4UElO7UjvRU40y3HF9
wcc9ZCGLpz+jkkuE2vpNgshlfAIERpKiwNB8b5H+EufthYdU+REvXDcnhDtECQKTrTf5oZf6U2gD
UxwpnP7FmeOoqx41g+nB8mGmkBjFGe8NEk6tqCfLIAHzZV8ajFykws3C924zwFG6ufnupLy73g7I
NBWRr9/SzZC+aTXTWCQ9zlIAjhxV/XLcFXW/O8MQtPC+l6UzRUiP7pqGo61GJ2kveDA/0ibGgLaN
MT507ZWWh6SXqP4R4phHNta8MHC7OH0FWrBq+CrS1zMAIk12//zxydUybNTPsNjMAiOja7u/BqKH
Z9pT/hKJbD6uYb6daqN16oRlekOEWN0A/zfhZBL95H67HnYW25nv8ryOMsa6yCC2w24edV6/gl5L
13G9x6Ztnr9tLXewy2aKQE2Oq9bV2bZYrH5cTG0HE1hAD61t5YXv4wPCtwnEPvb1inQrvs7ByCd1
8hPFGUSzq1QwVTY6cmOHD87OA/XyJUzAU9qv9CqUlebUclYg3DVwnt1gdzh7+Gsc9LpR0Lv9iEA8
7n009LzPzgw6uPEV9tHkLJ6J6jSIUNWxyYhxvaQmdqssjMZwVynSl7Q2KRn1Ww2i130HmF3BfAAq
g3lUU3SJFDj6UihX5NVfMM78KDB+Tevh0u3uP0Dni2dG37/24hwTcxaqvlRXZKa896h9BfgD0OVy
3uwbGPpBY15dR6nXz1X4VC/X0n9EHoPC/Kh+tYLdIinkAAQQATspgAb1MHzfpCcWrWlvr8j/MANP
A/Q1VHVxX6+DCsTD+BB0i91PCzTmHB42dYH9tgTKRZsnmFC0/EKjH5+oBipgErn32V+AO2YjJ5v4
oE+PD1u7lbyjdpak+rSQgCyk/q9UOth512KPv47WwMud9uVAMXVW5I7oI9udbf5PGK2x/YCUf/8j
2mIsvQf34PsodLMx1nUBiD6UiflPtntJzgfBV52s/P6sKLZh1JEQoHBqjLCCQtkpxWpkUGBz1t7F
X8dnQGzuJTH7f1TIbrfjJqCY3hlvfMbcgXiNjpIavs6VaAfQLnsKpt+MHbyuuKfNMlvP2RU3TsQA
Nf9vTvm95TZu8dSTe4zVJY/FEGnkFOu4o5z75iB2Pw4kwlup6PpWcRmYtPzPyDeOhrF3b5bhJYBq
xTrQI7+8+pk35/UH/NwSpPLS2+CjCL3njnXOOYj5K1EIL9mswcoxNZ0KVrh2O1ZYxMjXazb+30kC
7uMlLWTldQsTzQg+L4+O2O9O/4coHA33gORx0ZMQrxm5+/3PW3bdmvoZRFG7vpqKrOuSsBC3cUsz
cDTvrj7aJ8jvydKNxEnIaZfYJiX4faAjI1dEnQLtJSohWGBY4DiE/7buXjKTFaVBtwN2qEMlMepi
sIBmU3jYDehA4LqXW4ps9lxNmludw87nXMba+aqOa7s1ZILncXEdbClVcBsts+Xyo2QUNhXc+nYr
zwN05oNg/mUHzRC+LzM5PxrHz6wq4o0WCwt+lKN9shSwCIZAKngQZJu6Pmrd/k0usHpSfqEUSBq1
7ItMuczu2FZiwYGvwdku7emR80jbkPNUv7blafEFeAEodcDz+fvf4udg2sQJuJmE59JrxZ8uALlT
A8GgJ7+IcxGGA341LxmfsUABlc7GlbgEDG1gXcCSMsB+wKSsSBk5rO8jsfT7UHtdFX0LhCO+pIC5
c4ifSOLXap+eDV6gmSDXuZMK/IDlmUd2bPRlwC3wfJxYUonbG03Mw6YGi4C+EK10MufxqAESFOPL
E6UYLMNNwS4qRzQKeCmqIB2wviTKilXfsLRAEuXezAlrWx8NYv0a45FtHcjdxvyakLMEyn4iToGY
rFU2WRzLSflOlFP0YbVYowBxZYE3f8NVg5S5vjOd/ON2aDPnzQ5lM6oESin/GIzh6vjNP4zHh1Jm
FoStVn6vZqE7ZuPM1qN/WPLRqZufkLrFHz+mmxGCl6uqy+buJnxobsi8TpGhMhA5M1bE4Yx313d4
XEUu98b32boc/HuG5wEsiiLXDHedxzWGLbjRV5Aoinjnh66mO8bMx0n0BXlaI7+0P9gEH/ztaq4P
OXqsZ54YCeGFNgaIgusBH8nmNMJaC1uSSVu6yDkYBze8ya3LmzUUKzijvVlRbpPfYv1gQMFsxoS4
GxDWy1EJgcjtI9uOZ9CBKyF8y8FplmylX/68VSL45D7qKEz8+wK5THWuvO/+0cjwQOE06avTAhYk
JqLraO1YJyHlBZ7smqVExkocQDiBoN5cxOVRYrObsRnTjp6l9qNYigV8GuyauVOia1AFmCL6HZAV
t+iVpHHqF3K60laXprz7jvVsMigTTOa3AqOg/ktAQOLunI1n3RP3/eh+UpPLfvmgqPx0CL2+41Ff
hGm0qfD5L0+okhRAnenV/H5DbnPjM2ySRyaDyfGzCYrWoNJNjKpG54G6bUkf6LSM/lDPTk/ypgEH
SGlueXCp3MBwrsIczIKFQj9Jsv7Giio3A1NfssS5m4a8AzcjJnZHEiKRHdGi+asUoJiHpuTLRFP4
6nFiaNmcYC5rOS3oWdxobsrqAj6NPmWJ9u6sRdGZTWJwrsFoIQxcJOFrMIBHN8ZsBv7GLcczIV8w
36EIX6OhQsJtQlMjKMIiKaYDZcI7pG87/iR0GIq0sfZlkFKCjXq6fKJbq2eBzwRVZTnB6/2IOiXZ
Tg5/ei4KHkCkiIj0kc0xj/mz3HXK94L9lwVq4EaC/qAfrXfcmXpclxDfZgMuCNL7noQeZCXzOGol
59ZBvdK+OMVUpREJCIQXxgc+/Gc7wV0T8NICrzeVxDkdxVDkV2NUwg8YTTo4QX0C6lGn2qfKH6fp
C9jPk25tXtpTpx/nE9u/vdlewTZEk43HKLxs6vtycHZj+e7DM2efA86mh0bAp+XDwjzNy4MroEZA
UE4uVWgadC78/xyDNiuETAyKYpn46RN40nF3ipdxXKdhfFlB5CZsO4KFK/LlB/LYAqp2Oep3D20j
ZEsxqmiMCsVqnzvKp3oIgnUb0f4wy82pnwgOq4Do+cVaLdOeNQXEK20hd/UNeWPPaBnNTKBGVki4
rKt3WSoJJg/n5Fyyrgql7flJhQOqMWyPnx8IAeeMXxNh/kz/Cap7sTm8tYsx6anqiB/zYZfd7X2r
KqmLP80zh7cmpO9l5Z61MbHlp3pM7hJBoGkAoVtDqchktNd+ZHXZVppzN4Qw8MYYRiDTMq2w/1TZ
k05N13wY/L8KCYTQVRXkAw1teayqUfq9uCX22YTWCFsmqWMiVV170sABABAUaURqNH6NsftzJCKZ
nZ8Z3UK3/9B28PXN570cxYfGD2+T/1zKzpqBmDSKS7R6XM9A+QveSZnQaxritA1emNiozdtn2yB6
H4XF6HVIMOuefVvOVohWZSfC7gwEipgZi6sXeYOKSXsuMB6t0eYlylqZl5BSIovC8tqmca/dCLbI
XAajs/zjG3d2ePu8lcL/Uhch0FAtZEDPq2BzWVxr+9A1H1Vl6E1t6HsXMpZ8t4C8OMlQLvlIec2G
bZEGXE+5HZ/fLQNAiOxaQ/9lmbj7rfhgtjC3rZFoJeAA7jGVQG+ytvST0e6nIcjYL9MRmr5j2iYs
nlxskB6QegojWhj/0nLoCYPxc/Kfdf2co8fMYzkGSzeJ9un4Zw2Oy1hxRJArxNhqmqUg5ZwwzO96
ABM7PsSNND5E/2A8P6z8NurKBl1n8c2x64EN0O0eMvcxUDSlA6sswCrnt6U8wIvHOJdiccrE4RZK
MlyvmvBp0pea9M0E60Ai2xCQZj+Pwvw+L+JCb92/BC6S5FR/Dowj02k568JX+Qarz3Nu7x/6RctP
xyTo2RnQRxYEI/PudZG4vOb/oEB+qXq9RgeB7iHYdk4m42A0DLVvYZa7mgTS3gUjGLVHMuGPFmsU
LPkAHOpP+Uy2CR1z+DC3TiXpQ+0dIyZ2JGRNmut5YnRFgdpLHxZabXc3K8FWOfYxQv5hXziryCDa
ITWx32B/5Zd7025dKRIzNaa1u5goe2IYjotGU0HKiPwIi/gNY9Hu54Emue3Wus68b5s1LZMhGfnB
tyIbRm8phvrFtVX8iOVjZ/mDGnEbgwUbXBz5xiN/4Luw9dXAqOdzIoO4WX69KZ6VEnclpFXw3vMp
gVnevD4yM8MDvFSmaX+wWi1EoLHITiQiE2X9ltzFSmP/apnmYIHrJmrQx2pC3T9BQreFhVIhpMT0
jaQ3MjVO2RsU3vctBTUEjrnoh1YxKaNB/iBj9agc3bGLYauAc2/dmA3/pJA8J9HZXYbGKY1vQUdZ
7wbaPZybAH12UBJ3i8TJZNg9oF7HW0WMTLNIVu1/aC9vU8fsoU7sC3UHRdYASd4HX49fxJR/6WQF
du7FHhWj0XCEbu0S2Q2T3+Kszt4s5P35ssMolvoYxu6m360iqextOhTPXp7G8AIDZx0xCTL+JYni
GwCWNogYcxYJ43n2e2gbQ75C0FW2Z99szxa6fHIbkpHL37w1jbQy3DyRZD2MBOiD6m9YnAwgsUMq
RuKr9B5CygFPsoqiCZNbrOt0RkgldtldZLE4uEKAeykl+uJaVE4bhdzJtxZftWFEtrO0eD0b1PTh
tZYOx1cH7jRweW8pFLPTdCMuY+jLcIOVSJWxiu3+PkILxt2xbunJGPiHqUQg5JJcOo0kA61pHkPN
VM1OpWeGCcplQSdNTiM7s2BjVmL8UkTR3Hrpu5mLveT8F+GSzw5QGsZrt56E72qPYpWj8I5ih8sC
q63zGYX+bB5DLw1Yoy1NRHK5ftJUn++udXeA2b9d7XnGm/v4vFus6hYDPgKvMnY0rrwdG+RbMQJv
FnIQeDj33VxR6PXuiwtP6MiH4uLxeJZAHVEYOyMQTnnVeK/JXXmZRTZpT6x0ZCOmeQCNbm+fbsWF
DeNsWhuTPEHXLDNY5b83ZistU9XQ+r4i/DSNfkKdVTyQinNOuJ8PUvhzUJfos6t5oJZocOLrEEFK
mfweUJNSXDgB2423cqTPxrIfzMMeimE5wFonIzjyvMAvh5nnfUxe5QTA70Q3Yg/jpDzxXAHwRoAe
9rbrDjLZ9ZYc6eSz7hGFvQa0bqd6ZQ4yynJY12DS/bfRgpe264zt/jMp8v0PLkxH+cKb5fEQRJqq
+Rj/RHE0pmYMNiNI0mStwbS0xgQvrIkLi3QlInbzXpAvZDhd74fOR8Gsyaad83PqWZ/40c3y3hWC
Ihsxj/7KoRW7XPcLSmnTNhf5mRTBTgLE4pGW95w2WcSlg1nHrCXNaSnrH1+9RPYdYb86qXsFfxcT
V5zn+I0ZVs5hqFFmiJxI5jDDmgOnMPFHU+DQPzImdO95jO0MEpqxsrJr2fCSbTT5U2Gld1m32lmc
fxQQRgZbjasIlqo7q+/dHWMKGYk7BQ2ZIPPlty3gzea0QRc7G3d74HLblld6rnclze7qycr7/RdR
mDW2fKj87qx/y9+KuAlUQQCnHWvV2uLH8R89sVyq7S49ENX53olnrr1RwSqQKXbU52TrB7tINNMh
2Ce8vseYUoA9NO4UipmTFcuE+4UCSBBhComjhayODLrZZNzc1rZx/EryRKYJje6/NtWnlmL/vzPT
zpJI8rz8x6SpWCp4tQnnXW5TSGEu65K9SSOyJm2WJTVhzu4IvOCZg6j2YwwT+9TQzcUVuHXbYZOQ
8BsdvVSeRS5CyeOukrAzF34O6fJZ/IyNoh4qEcT4nTIN4AApf+UGjup+NnP+rPkU1P5TISxkoEp0
kb5TCCdBYHfjgwu6ZchQWku0tgDMU/4ESJCDk1IsZ++6orqeBHKMAWBZTm+zHG/pd2N8jC/Gp9DK
RmWpPKkkzU7PSmzuPQlEK8UGjHU/tIU0ZCP6tWVz2XUi8yamHupQW8VWvQxEeZZWIOiEodhxXXAV
4SMGKs7h44I66ZQAshlFxiIneoVPB9xruHU+u8pc0OZAxIH7zb1pSsCDV+7gX+vgFhEDEsK9agk5
8CWx0zazxkvmxXrLXZhJU2ioaoGOYPZUOrDs3qJ5ykgCrDjdPTVuepfEbHaf3/r97jtbnQASfvqe
bSi2hDT5oR7nEMxfPP4exoSrP9onNFCxIUoJ6+ncHxoFD3INhemYCDE1I3FaaxEsg9aip7E82X83
lKlUXJSELkbSn1L0Xwqzaet6gcX+/0PjpalRYn3ZLTkC5uZXjJQ7vw30R0waSLSfTQU8Xc5HW2ET
b4WzrirUKi22yNnYmcy941Xf6rmkJW4yy1OOXbTKlL2ETFc7mTAzJqgeCW0lnEJagFOReNJKNzA/
bwALxklfpg1JgSV5iXuIumoVY6/euuwAWJ3U18WPQEp/NwjXzyiCwTsfkI/IBOz6Ucg2FAhTdmoW
JDHCNvpZGOyiXyWECWasmzvm+Uf3FrxPWKSNv3niCgVwtIDPfhXfbdvz0skBwzBNJgec6CX/r4k3
buYbSTdd8S6/65Kb+SFEFZ0b1tUSjk+cZrfkIPysZIvAua6VoFvIS92O2XnxnKaI94FDIa8j1zjA
cnKOEUkrAWFPzigPqxACg3H+Ps7I5ItA/RoG8b0ezps/i6wj1IwPf6bAn90G2ZpvR628/RVQ5l7S
VWjaw/JzajPSJE1nnLHgizu4X626wJTntRJLx9GAOFNRfRbV/yLTnzNoPSaa6ydLEIflm53HnHTb
v3A3RhPZLJsCpxIEuh3ffnSdcCsQZruAKS0SfQf/fLbUb3T6T82YAQ0t6nEvKcqS6GS/EkTPmNRO
Xluzdn3Oq5Xh2IbgDou0YPTEb0JzAyuwnt2SSzj6uv/S5bzhV8+anrcphbSKXgywYOhlE8k7SbGM
dMJLA/1aRz8SVHtNy+R+y3yIhUyC7HBdr6bv4p7gGCCo/Z8T/bckovUnM9p2qE3ygDvW7bRPNWPN
Ox0ThGZqgsDlx9BqvAYFaypyN4Mq9Vx4m1oy6mfQ393pLCr2qdKOgn3qmLM0B9UWypZVCynjIUj5
+BPFqrkxYukbpZw+N6DjGzF0S1pLW+KP3A671G5FJHujBaaM+jJwjl6tplI8u3Hm5Eiz7dmSkUcn
mSfnQDuzcCiH9iFTn0UXemCsDMh70O3uRoAMxjpWpkGL/ItE0X58gw9Ab/tjmFaLYVZVGxn2h21E
5qQNgSlpNEB0qeAuoDe11xAJWZbjNQNR10DHQzFy7f8P1k/cJUrCzGJA/uzYTUd5bb96Zum9g5TI
It5HE3lw8XUViwM46hZT8+FNKvY0wgGoodBiR68gXbyz7MvAyfDF0qiBSMgsYTDuRPcwOiF5NxaP
ilx/CLhD4e0NgXOCjQWzHWF/kTaJ35OdWiXkbCE7zO2lGnMgKUsmUnSdxMGXkFhQa1Su8jRi5bQv
sMxJIwiDT7xHJTWLagX+BG+4cUmQjbP42ZaS5qx/Jxj56dgeVtouVJ3W6fVa4/D3BAHBWXFNdgvJ
mJ0ZLk0G9mUWCrkO9BXkgZ/x74BJtoMiTBUWIY/bQMUd/plVsw9K6XEtIM8XmYz1R78HxyyHJYSl
ft3qBBieXDiEie7fldlZxpDkR6XL9Gxk7FWvdTAT99DPNjZEh0JotiP1q+aQNHV0bXfIzTZlEMy6
C6o113Wo2W00QYhdcTagNf7MR32AfQsRpiLWXZka1fQMND8G6fTabri6gbWYfgpn24Dx2LoTDjrH
qgakF98df9xIQ4IEp66OFStlznpaRJU81vSOHhM/mgF/mCOlXhzTTOT2amJYKA36yaeKruAWsJTA
ELk8ePE9N2fPMk4hJDt/bguCAWQXQXz1Kz3fw10KZMONfeGJ5jBk/WtgkP7IHJGQ8wp+eSfqR8u1
trZlh2Xg88ue294w5zee2MbkOe6+G0Vzw8QzrsJ/m/sNzvLMArmmsCg4eHfDPymGvaMsTTOrfNFd
qlx7cZsQHnEdpTGqOszSvAPvyYEZGyOHpui7e11a3qcPbsvYBeXJAcLXMzj8LdjfJb20PTezSM+r
m2QSlDubLafz6cwo0UQEFJ3ampRM1j18rdH4LT7BfPPN4xN36Jtp4EZXWaVIGC61E7W5dCT8FQmE
eMV3u6lIeOPbj0cYOVA42auyIr3d6slFjVvR2XlNkEEW4iby9aTc032HzDI7PQchJT6DV5Xj7Rtk
i4TZ8fiN0Sh8X9AfQBQrKOs/ZShrnqjnvWenRK5Hl4H/Yz3qr054A9xPwrj/eU89x18mTL2l4SOt
z3AWh/nbOm7t1qBxXonrWxmvzPX6c7OhmNQP7ST3iSKGD1yWxqmJLhEs5EsuTA8Y8JgHVhJpZTbs
6F7omxBjBc+SFogz03sCw/aKadATumeW4H3m0laWXJr6li30ORCmmTGQZ6j/QEYbLszwR+DSOnhg
odVQEMnZMYjjdCW+51UCh6ZHObL7y0nVUDJX1v8smvfG0wVs9s4lklF7VYitqIj0xTWNlI20hOKk
+z+Rk89/Lh130X28zu0IXh9hcH+23lE5fGkIZKZrP5JPU1pPeEZuqX9OPj6A6D1toD3ypqy8aeyO
ajaP+WWEQKEMOiKzSAG1pP6IDbVefDlweGE36dcVDap8BLVIT8Xci8C+5YtDZXV/aPe6HaDHrIhI
ch/nmoe3h8zz/L4DSnHSNl0gu2plo04b/cuqo7arZS+DP3ONmcWsLTlmY3yHcQPqnFcYQCfL5Azf
fVcgN9/skCxU4TeFnYA4MUSbbN/+bN9UFQrQ+WrXQSnzHpcwMarDcNxvglwaY9H2KHbgzMIfk9dV
rkodCAd/t/xzS5AGiukhxnprrUT4LluNOnxihcY3cPvVwnopTe7+3uIaouMVfN9H8eFJ8gIOyfc1
XymthZbgglix/iETiMb+g3ZIDSjpuX4YrMX0WS10ZXDQEIK73L2ue1tZp/CkHrFrxK4RCjm01xS7
qja7SMDow1CsUMWBQrDEzYjxPJdUiajnTB1rbF7b+Le/+0HUUnrv5hKC3EzQjED4RJdOtS9H6nH4
pX5vQp6plbQXsCijAFEwzuEXTe+e1dmfyy+BHgllmDCf0uOzFO/DjqrnH7Zwywm8tOgJYIazmc7J
6rSan52EKzAxN3ZM0KgShWRL7BR80vf3g2i58oIxssMScc0bUlD78NsNvW1jEJHWt5UMn0DByowv
LcemSb09e7C9RuihI0LeRqE1zAGjbUJElJrHNnN+1/9AMweomUFk9NTC7WzEPV0tgD6r0JkXHAjT
gotQ8TwDxGRB+pj6/Bsz4Vn1vjMcKZw0yTbU+2rSVu7mFwzX5tEa3BJJ4QF4Zl9a+NWCtlmSVqVL
ITss/ZFdE0b8Y7gUcaLV/0GqJ7V5DFGs1Mj76I3mcVQLm5wgSj0IoIadbA51jFLsOH5uMF6j9vYm
Lp6yJoayJmlNv9Dnjq88XylP7ghjDBFIEo1ISLwE0AORvkrCLU/DUSUMnXvbOmbbykx7zPX0LYSI
0ojrf2AA49Fz/Yqjy3PdLQfTHFbfNYVeowmAB2Ws4DiTqO7EZOzNAIlJ0vLNxf7IIGtuO5bejksQ
KrGjVMEJq5lhCB0jBCw6bSDjb4i6aPwUX18VkXE8S02f5i2cntMsboMgt2xUDGfCsk1t1a6B64aU
ty5hNtwKW7+2fVRKKBgZ/oqWjnqGtLhHtJpa3bZh9qggpdg+hfe2Rd17QqGndtnJcoRcUIu7r/lk
9OdSWb/2vWIHlNzHAUWDmkoErIPLqwyg6xJwGr7e223Usy0cvX/h/BZMWzdXT/OBuHvKmZNa4194
0PiqJLN0qjCEK0DTFPM31Eyke6hPsBhmsYNyWLx8qHo2egS08XyHnHUD74BrQa105KP9muwojgnQ
h00AEB2nxbMb5dyislKNorg+kRf10xGEOgwf06ZBgq91aWFDQHGirzpD81PPQU3iwu8q2FTw9yeJ
ahDMQUappyRXuex4eYluMhA1AlVjPsadtunU99MK9n0dkVi2wMb434B2DJiw67v/ABjLN1CwmTbI
jY4w0dKRGI5X5yLDUgZE9o0YAx5c5aR4oPgVrt97nVN7pvFC74tgKGlmMX4rFLHdeLRNuDgLiYE/
4bGYA1LH41pRIoOeN43VtYmO33AFDF7PajFuP/hIrP2IW7/jjVeaehiuOWWgX0iyDsUgyXl0QPhn
90vdvoG0XTzK2Ihwclj9v7oR8lsTH2w4BnohrVpi4mV7jJKUYWnevHB0fNf+GT3yKBplPgUS+1jn
7uoK/xIL5P3QLGqBcDL0qgwYiO+l54lExN0ZyjxN7RFTqfjzW9cq5I5UI7DeKyUwWdxr/YXOoDS8
jnOgkbcT3fvstkJePQRYz/+cUa6RjFpAUk7pTzCAlpHR4g4WBj2GxiTDDgo/g02U/xa+PcyyjvCs
9DWJdnVV3FThLJdFFYLNR/O9bqadF4f2jPeHHjAkGvXdC1a+G/LHUpSf2NltI+EnBwYg7P70kR7j
8I4uGjLvA4i4PxODeIkHml5AcAKg9WGk0aFVMgp7S6Vlu7ZUjJ7o1iHnX9IRIRIRcJoPTiYU36Ec
xgWIRReY/S76ZCokMQ+0en6z7rpBmPQnL0o1Fc87Vj2RXB1ksOoKVO85iLXHO1mP7yX1Dl8YwjoR
m9Ls85XOHc51STlu8HUcdTWNJHuGjEG+1yqlGmtUb8y8tz17MrHjNF/4ThGTG9XnNliBYQ3egbq5
a5s/DheLHQIpulmllo4gA4Qp+uVOf7CUkcMmoDCdlR+NvxLmyLIJ1EhPvXEUHB3mKxN7mp5O7xtN
URrLbqpV/fjyBHYLrQ7SQ48ko6+kydcKmbj9/JB2jZyq/OK26AoDvhJNQwrhH1Hz2nh2s/OhVX/G
WoFMJ29wq6Y9Po2UfsrMf6jeE/sZDCyNLAgGs5Ap0HzjPucx+f9tJJTDOKP39N0Kx74gcJs/4P4S
j648XSUnBeUZffNKVnn/jbzBcZSLfbc0BdIpsTn44am/23zlnLzXi/GumX8qfwTvs3vVNB22slRI
z57Hga9cH7fBQ8OiKv1OGSabDdAaxG8AuJQbJS/sCEViNrpof2j3us4aJbZ1LXaHRjenYHLxVyDn
kqSnG0XAGFR229HIPLZYPxdALzmdSLGIBVyVCAwv7N4ejDgRj7Qg5UD4D2Cku43LX3teP8QSMl/W
LnKV2CBlakKqSADYKVIctDEdcj/IKFWeaBRQsUY9BvYyAxMgo+PxN5xRV+50vBOZUAHqJBVUuEvp
kcUBkBGcddVZNO/2LkMZ8zkEvhwQay23xBWoKBwvElJursNwMfAiErcH4WVi+C9Q3wsHauasrZyL
7r71yYa/hpKBEcereYTmWXlNseoobkDmSIIoRteFdVYYuSzoW2ajfAgTjtA2b1C9cxQJDmCuUGcC
XSs/Js7nP1oHjc4Pk5uJ+kipLvQPoaymEIXrn8luR0IOlLDTtkUAJuGhWzER+qq/zxi9SpLKWKZq
xZtYwyKhOt17pmheVFCkuBBoNxuBJb+ae9cFVwHC47BT883IJCbhnWBxE35X1Wb1AiN/cozkydQP
iO9+I+xpGTZWxeFP5zTBheBxixctUhUSKtYFWeAwiEawpAJRAnfSaYBZIEfSsNkfA/d8nYhAN1oF
S32S4GK2YMOH0knWFaJLxkoH94CKXwX09z/RMd5aht9C66kTttNVME6+9NsG15NCull9plp4bORT
zRoVWV4snsAOytogq1Vna1lEK9mbwunxp7LGusWN2gRNFdLMrDy/SoRXe5VVTAoSmeFvsiVFFuxF
deP4xHy5OONMeOG8fkeukm4nOPj3Ry8K43dTXZVMMrt2d3UmOAGlyfL/vHA4ANRAcENoKC5PqzO4
p/BOAtQEuV2Iyhf7zJj5qeC1eOP4p61d0VG0cmykT0/ZoVfQtMauP+/uYaLJjVYJJqe1/OKwoIvY
dpMlPUyRSepsb282PwNdZBeTINICa7vvS7blTN+uVRsf11RKBHf3b3L7GjSqF4u2dSV6e9r1DteL
1+BORYH818TWHsN+TFLgtMgJx06HlYrvXKyqWXNIZ//lPvWw6oNKJwg4qq/3kSf7JUcGzgr8CngM
E50UFFVfof2xSILhKdA6jkQ6eJqefeOE+81COlQLwOb5TwhUTj6RqFzZQ7kf3nREg5FKY0mxU5ov
zKIXYNtMKk9561B115obPYIbaQ5xQJLHxfKcQ5ZQCEtA9BQnAJtoR2Qw9TSnTiWE7dLz61D4e7qL
fHnK9oE5au85ERAV2zZ/jNcnDlm79mQBXSWyOCCF+K19nwzbqAlVCKEgLWOTpNWrCQr/hukymDXI
cIFSE7cWNMOjHJfmLXyANYBvDgDAzLxxvPn8sRFEiOarRnsoRLQL2fKokmq1pIZhLbyc6pNQQYiG
IUBN3k2X2DMgK9TMAKmbfmD6p1Uf16ADnhySFjC0IBm/wdSWd1TAuFC5HatyUdZ3DisBWa5Vs4/e
bf/iP4tCCRO8bQpWVSbqUOVWBQrgAbwv1tocmZqkjJAc5cQg8Tam8T3jGWB+sUX/eZwPtcTVGiUO
Xpg7kB6wjOOr4f31oiYIPTnsypTT9uViz5SJp+SnNNVDgWdURwsfsP5/wgMOh8YvN8+spKAKzoqk
41X3DLYx4N4YUiHyTq+p2msxbR/d/7jkP6rDNL4+gg7zAcXTbCOacfpYswhp2BnteQFL5HwoiSJn
qPNGIDEnlbewP/0hZDOztgYfWIHM6lbXxzvJdffKyeLZqY8CBqCLHobSFIZ29hD5xQfK4ZgAqXcM
QhJoCmg5NGXdMh/wCOyfFxKQgwrPcMcaJC2swPJGOONG+e3WQ9Q4xB7Uj3C2BaiQBZl3DblGonms
C976YFO4kH+VQm1Hw2mV0hV2Ma+gBoDWBrlH6fPAzgzPDB7Ny+uU13HptodTRJN1/CA/4YscmzFW
APU2TDTw+BdLuSyiXagr0lUX4SzEqhMfBh5RHvEYDr5Qb1Y/BN1hQGIaVZ//gjdbiOKzOdf1NZQo
W484+v2joezmIIK23ydR/JDU10JfDA2xhJavuGXLiCMzonWQa4YcxC+3rBj/Kvn02QQi6TAp5EUs
Z08kSuf4nAqp6JuZzA3jO/Mj+649jeGvRT7p3cBv20+vJE4/p7Vl8h4s5Zi8nt5bbif/oBH7Echa
dKAshpodqJ4+5MzS5QvmJMgElSOzj43Tys974lCjneeeyBSSdDicYVajq14OjL5447s9belAQZli
TWTKZSnfLNmPE3aFgE5PMnyKmMM8MpTF1w93Nd7HiBmKeBLuw+diahD9RCzcFqGc2o5GENXKWPKu
qAXomHBaCw7j38LhZ4SB7YTFhrE2fUQSR7CPpzuR+FKQKzVX4R5fHSzhputhFT/RVJ3UgGrhKL6Y
L4Jtt2kVrKwuVG1EqvMlgjCJhPPjyWV0DFc8fQ9rTKIueYdd/dZ22zO9oy9nWl4GpRABSC3Rjgyy
ieeQNR55xhEe2p5a+oN2mt9AkZfnNcdGxV34HIe8ZfG/tMp10uO1VsCQ9hSUxHxUi9o2qtTe3n4k
VM+Lsdlp6W3/zyvzJPW42lRi1+7wJ6HeRvHaHsr5hbeXxh2PWCOZQroKcVwcz52Ecu9EvoG+1j8K
BZXZ5rbYtmVKFA+LvdWxsmRtATw5byIGWW/r5hDhWAiU/LK6PQE+M0MafdBzp9NygiJzY3KKDOvK
iydlaQYkr/ib4XKcLUD2QISilekL0AA/MiCe3yI3xI4r91u0dYdB7MFLgraUvOoKoAVuFBO6plw/
xB357EkiqdfoCd2Y3Fll3El7IGyySooA3g47crazFf0wPK3L8RkO9LnUEK0DCJBcdOboxIBQx+Li
IcsNCAudjaJHcBtMhco0LcrcR7HNkYxF8oUeTw+TEWIOUVZvoCimSP7GtnY//NyxbJIXYqYj0vhv
Xd4lajBh3xTjhoOPagU7enBHh7JV2MoMEgbjqjG5/z5ofenhKQ3hmXHHt6oygi+VD5MT1LzYhBbN
+BNxbuHmFgKtM7KVU1ylm3As5+4symjpfZAqN+EsULM2oIztTv58CTNGbXk4SL1PDb3pRI2lBgt9
E7YRrWo06wvkD5snaSfvYZX76ypdeA2JcrouPKTEzGs5/ZF4TrH5nCJwOe+SmSoqLaitHEoaTan4
6a+Ht7OS9Y4e/40yVAhuLmcKl3MaGTO6ZBUGNjKgWjquE9i6xTEnMBjbIzAM52Dx5en2R4rMPgVg
vuTlnc32XroXBcrGtV2rfPRFZfvLdXuUxdGfVrdLiiCjGzFldL2RnUF8IdgJMt04LePGgKU9K3tx
U+dtr/Oniesq3mldMGMAmXAtEiH1rgXkdWn406f7I2gxVLxteLnfX8IQq1Iunhp98x7K1jK/IrVj
DyTkYac2iyjttWsGu++8tFNepCiAqGIgnIEuuI8VuqhmxP+8CSI5r5gNu9ngYwAkk3OBkViKYalK
zeqSubLZ7ISbTT/xBQsuEjOcEzRQa+bq06sc2L1Ld5aKRs8Rwp4D7MZyD/vNXtSQf8h7Mw76cFMT
KOznV+TFH+VCpaCE7MK8p46J7Sy6lhvTVI3/T0yPtjxWyBGArWTFIyA0Ax9dCLZD3e2iygftvSAb
XPj7ifOxBqFmFLuWuhZQ0six3Dvbnz0inKH2IVFFQHh7gO4qWqJ/dwH31LBq185NSNjlsWXthabF
8hmrT5fsWnZHu/b8yJWMPPk2WpRKwmIocvXJ8NkfRN+tX7IrrR6yoA7EToBNsYFV/0Vmw/XKSmUh
9DY5m5i/75tcIyaImqVxRTgbTizrPlJPhLKdKUsXDhuPEI6aAM/jGXxOQh2uqJOqMXCdMd9iSR9a
QE46IOwf8SGGimFMqnDYje4xPzNiFc1bVigiIsYgjdUZtAbpXxP9KtsSAK7LTyalF4MG5f+0nkf2
RgyvSkvLneD3YeIPYinB7Jtyzbf8qLLsaIxvd3NFqmqYfFr2E+bStSplFJV6rqREJ6TicUvVMLIc
wf61Bs66VUZfh+37KpCDvHKWSa1bpOwykm7GzaCWhc3u4CzQDtyJh88pjR4xlGH+872D7qVf33u+
iiXYZubnKgDEK8Jbnu/QHxhIfeRlDPR7dzVnHNY0ohbKwcEKkAMDY9MDvFOfhJyzT7MPx+gsQxh6
a7r6lzmV4vXBFgB7MbYALQ4XNznI94+t29o7elc1iajy9IEDlNR47HBqugzxZoNM7ZqpXgK5NjYu
90567WkF/Ra4eBA9RigvTjsX6v+6AmS/g3/yfviehSVepZda1FKeAlq7gHch5RpzZ5ywogya2rDu
dXMGuvhzFEg1JLIehnx3kO4Uo+/qwrpqY2MuHDSuU04W4hjYVSj+yHsKpP2wZWwd5pxBPpsaSUbA
t0tjW5PF8izQ//UjthvkWFbOpbdJS+NiblLOXlfJHj2jNfTWylra5v+ENZ1CpzvuagvBS+oKWwPM
keLD2wMAczIzwESzmDgz7q7t2CZP2Fd8Ac2zK5VcANe8Dqe3/atC7xUGyBfzTxQolZfGeNyX1HX1
Gn9SQTiDirqhOzQEgkL77PJGllapMXh4y2J7TrYTZDN9v6F5pT2fkf+j6+zrL6OPeU/fm5o+K9b3
H3aXUjca3ftFLoBZzgrUCG2IEId5C+AfiHcVgs/q7sOTN9pIAJWvfWUW5ft/sUZv48RjOuWO2ND/
v5CNnuAobA4TdcEyEW0ZiLcfiRQfElBpwfzmnXj8U8uORlmqzUUOOaOjHteBXT2z8wCGyVLGLr8K
hdjaj0zZeXebGvbST4e8H0sMHvuK25V8x6k10AT6Lay23a5gYf0Kg++Jciweq+HYs9r13gLV6ARi
ZZmkJxHDcGd8VtsCDC8xoV6PKeBoNRgKjsUUE0dLZyJNhM0jgM4nqZH+Uz/l+cH9YD10OFAsZNg9
Wk4womXtLmoUrZ3G7gYBwdcczlAOwCQWVcU48Rhygj/ElbI5NLcvDzen1uHKg7zlda0fBclC2A0q
nh9Ra4jLP7oTbTHQ9jm/qiHgKoAo8LdX4oczG8jS0fbR9HAqKeZgpkLapVzBWmlurDuegGGwFvFT
B8M7WgCy7X7jN38/kOp9AmDCNJNwMKRBowkgq0OjJqx1wP8qheHLAfzQi2UGPBHM3k/Y3ET2S7nu
SwMWuz0zqQ97jPGeYfFZIFQQjphDhSfTwBmXOVgl0oj3HcpbD53WPGPZ+36aJ+MWE/ddERpLVVFy
SJO/sZqF4v9JfcIVWqxxB62Sa4PcCMtlKl2ypO5I8oF2/p7LfkPzrNoJmqsZiS6s71bcxB2IDI5g
qz84wsVzhhJwaaUAEI+sI7mLfezpqQ0zjspkxKJw1iGjI3FYyIhoNYpE7716uRYIDgO655xNWE8J
bFhWe1MUTjdLsiaZLHq018yCzTk8jO2edZsBYvoNAEXhf6BCYDunn85quLciyf+kVbsQ4/FjAGCb
elidXSaaIj+xfuZ1/3pi/kSx6n+wSA1xh2Eu6mgUqaCMd9atXkDTdI4PzOWAzQzm/6/Kd8KqqTUg
y5IDIdmDfI+1wcGqYY00+LifhhxjxwUMW31tSr2yqPHpDaxaHi5IOgc2aER1I8UA0V6IIFncuSbM
bY6fWWEMcRDst3ootH1fSHqacrYAH+TPHG8rO7oOBuR43DXiCa+2iZi7Tn0s/6ss5sP5gEBBKkIJ
/CKdeDVxnrmABMblICADL6BRGyur9XCBvhi1KwyscKJFd6G8Q2Xh63YVKqdliKe2Ei7gIM35haZd
jkKHq0ZBCAHMrPZYU1A7Y+W3eNhT1IOzX5O/bVX9mh6Vvdwb8vB8sOUaoPD6v8q7qa/G8Ndi68m7
OHaQllGBbhroQiLfH//qdvpQxv9buwH/YXiVDIHj91w9bhBEWBdwE9G4AiZfXZWtQ0DIlcIh+bta
u93aN/rMi4nlS3aHxMXZZgJw5LSAi5iYUK49EpHv8JYJeALzGZaSbIXGtPWC/ub6bV0EOHeNrfdL
CikbFjyLUIUlwHOuA9LbQjnrYYQgZs5D9DUjab07gF3J7Czp6fns9/55a+TuQ6cgEeFoJzwk4og0
5BEP4rwNOQAdOj61uocvuwpH6nRPSJGsh4py7BgTbZktYD5R/9H3OMcRCScAaCrm4oQgDZv3oB/G
xT8C1T9X/cjFwxjw82tyUoqI84nmpBsxbyEbXZLxP/Wx2uPjpcdPl1CsM7icfJezMMIDBxlJbtjw
VpL8AHwveiE2e6dNn2kYbrFm5WVWO/6kpcKh1kh3AwotXSibbNKXhczkmu2CGxrYva4ZSxFi5P0F
4CR33trkDl90hziUY82z40YfkzKoNi4jHb+C6Wx45G4osfLJeLRmiFsKYFFHLIyl06t0B++mA73O
JNVJ/8emIFra+YCscxvrgt5AP17mIXhUmrOQ9jBavbE6Zb/9WhdhTtVnaVB+QHLoT4xgMwGZCN2k
l+w3TBzaHzYRp3wcxkrWJHyKVM5dgOURV1xBcPxC9EReosRIvfkMEpYgNsvoMleFiCb2FYPqws78
wlEzLX0s8xEZ21PYWoezekNvLFk/g9dQV/Tv8KdDSOsWu+nQBqTmKqwef3G06kib2aOe5nHu8mz/
xHWLDFHIBcxJOgEAxd9FM0k00xWxW23TPCiDoUAIwAdCUhejtwucNg26djQPPQfcwnQCW9DfsM6N
U7c61HcT+NmVEw3UzOkuclINJfsBANPSk9un6XYeJLIfsgfKybyUD/+WUsQQifEUMa1UyBdyNWlK
Pfpec+mlHrG2wexA+EkWMbSmlYat5My+TaVIL1AxXuNWKL41jLS6zg1VKDTk57N5jH6Lp8WDj1av
lfXLGzymLphvRGfRq8Dd3GctvYpAhlw3E9H8jAUqTgeCMa0GTQfDXhUgvL3wXAkt0cmALPgvxLYB
U0Cr6Ja1YXdmTWnI5IDiwTmMjgGbfhBXaCXkfGh6zL5PTh12MqXu6+ctFLzpJ+Uh6rD26OeNWHgF
hrYpueRR1HC8tBf0mcI05O4/24JF5Q76gRR5ux8/CE3F5CmSI+3l8knzGMuOt3zfIpwxH1zAbAYA
lItfVqo4krshaEWiEtAuLF/I0B/6kQSf/yHI9WS8TjOmttuGTSHHo2XbSb0eGopL9Tdli6Jz0gsX
DDZaYfr9bA4YwvLeeDhTKLDoCc1n7HDTwmva3hkR2SRWTAZFjs4SRCItWlyufFhAGILh877PDLOK
Kd0BgjWmDc0bt9yInFrqbHKha6KoXUzTjptNzoyBTyVQSRPScewYtuu1pF4UQT0gAo+4yaFZ3pvN
lPheaGbXEKlVGTx1ihsZrJse104FZG7bATfucErI2nKf6+uulDf9MPoeMwMP2xNX3v3qj/0GGFg4
6CN/albJDEnPOymGIzckVZvJnfhTHGelKKhaAWqsxkN/unjJeLXPo6uyRmMiLoW0JK6cXUnlF2L1
jvMwOcJytpXDjOPKVlnei4vB5z+l7BqH/Deg0HP1n+6fVeTen01r/CKinXDVGyswlLo8Lo/CBfqx
wQT5bONaIkhJ3nTNlQsLaOom11045ugM/GxlgLt2rUqmtMiqtv1xw+QyDEF3pz0CgXXvrKILRJwR
mr47+Vr1MDVOLwsqjq1ZsXNBFdjB/aFXQ+NbVlqKO/7n9+IKNn7ujx/gDQQwNoCplZHtbytsj8/v
nTNAU03TJVPaW3vAgndpIsSTq8rNe4oX5d6qrV9AEwXHHuzDLm0TtgQLBx4B0P7tKnAkVkvQHn6d
YJ0N7NKBEPYhIHlheSe7VvBAzXVccbQ8+2W2EQbwfgAmuaYJ+/iTAzpG5Qm1JLZLp1OQ8ztr7o+R
u8pTZ+lTWjlj9GLJjGG9Ycs9K75bXyTiaXx/xfWRG+bNdKDVnMs3+EjwyAwWyQK3HTr7QLNoYKOm
3VB+1Po+harM3CfL8frwrpHf78Wht6kNyNwhwjPZhx7SS2aoSsWCkdTBr9Xe9HE7XpBU9H1L0RsG
/RJUbQ7giE4ETagVSmpP8/TEXCk22RWQXeObaB6iAVp9AwQnmiDdw/TY6U/EQ0tw9wO7LBA0/uT1
EazdHiRoIfDVKvWA+ppSWo0r+1Uh2uczoKttEptU6uH4Z/dmM83O7fs9SV/RoHnGzPlpAukvDCnY
evxRq2z1fbW1arQTGTQvVwAmlt+OQA3NsXkjv6j4EJjf41OT/DsmMPw1LRymhnnGlHYW95eOQMXb
HSc2rlv5Zat5v1G77Rfvw5XpsBUbGvGkYfYKr9H3zg4XsJhe7tcPuSZZudZdDF6ZQHVetsv02eLh
G4dYdiZAPYMTWK5Wflhh6xnIlfkTiYfq9Hne2sv5oo/Zjqkfp0xYs8pkEN3EBetiqEVnbiRpo+Hw
4HJJ2fLijMGvelBl84n30CeiL6uAdJVwuUq4QZUfXOkpNVLQ7DSw2lElpjgxrYImDabnjEQhy13p
jY7R+l9OdfJqXEjV/B66W7lC1hUQCap9T9PNfmlRXDRrcWDzXmbiqH+UDgr2Give3twucXNNAdW5
favQOLpr6J0nJEWeokv/uuF0QjVOn8X/jyjG2twP7h2t0wOhjCc5J6RAfKky6kNEvEZtUPPBp+Cy
ZArY656jwK+qBwyumfzsCVpJpdx1dN7JBT62zNvVsIV9uuPGXqJBwdCUipCi+BzyBCnr60EjUArh
39pI+C04knY2PZeEjnplUUzc7aTpXRFNPXeeilWSWwbhCb6nXxQsIQT8WlfCmwSj0rP0VNew8XRy
rwaSv2vIhpNR2pm7pV3KzOnj/gk1k5cz0qQoeUzG+nNrneqwifuwlyxcwnDo8f9/jjsgzQqOhdOu
9X+r6uWgH845TBbIYQ+Lb3zCynQ6rvPHCLkvVu+2RpEz8TCrMyHA+HdWvLL0ZLsZx9CqzN9KM2+m
RZfHhuRJu00LfD+5FiON6dFDLcC9CYxHtrwI/QAYpEWUIXIf7TbLczRHAs6vpSlHxPBZASCHVQE9
PlR3yzMa9VrsCU4QUm4zNGL0OOkJsdea2VRbZubCATu4f9mJvWfegHUO/8jxZdkYL4qqxMIFIOJa
ZbaLr5astp2le4MeWcNYqA6xjwcPwEe7WH4EgzoHuvoNPCqQWFP05JNyTDsAI3LUja0qRjqOQrrD
W/5VF4TJ5V7B/q86e2/IHocZc9dVq/QcWCKQE+QeQuRgJ0VqMdKvyUqsh9Ynyd97/ux2wYLo5Cys
HxvCBNQqPjgFwbZtZCrep/ntic9C1Hk8H4c5UvDFNoiqAuhr3iT0srEta0cLn+9UqaGmdJdkYooh
ZyRvJ6ypMWOrm2ZFBnCU5gGXDUo7pOR78dSb5qOcJ/DFAarRdp+chY91tWKEs6cTH3Svr7uI3G00
3X4oUeZWxpiJJtn57PM/B4jugDAm8OgWtKfXf7tsqtmPdqkvmvotEAmJXXt9UZDpez36kqsoFYPm
9bNhZM1SYIaJM7OUHEhyfLlV9U9As7hc4tulmZh6QNfxVOamds3lqk4UMxNrNx+afChXQH2Ct7SB
/LqKgjsNyYSzHOJJSgBCwchtBiPrtrfCyIuVwqCW8RxuYOBZF83T5HRw7Q8/F90JQy3LGBMjzA7F
8uMRgj9p4WdaBOue6F7NS5zf+3HuXNIQDPmIlimuhYxFYMmzgYh2XgIg5kK5VdegbpMCy6Egprez
kA20HVcAxqMSbLvnuDv7Bf7cxlktZ2MxNYzNT+dg5HBFwfOHYFhAlqaD6CMfmZI7V1DXV080Jsf8
6lc/K12lsvNDsNgQzgOrbJFxcGL06hKnJW9sx+TD4sTZIjmw38yscCV6/VbOTLeQqIaiHThNldB9
1Sl5bgKZPsngSHDPfKMiKxvvxs4aYLKjmZ3KID4KTI1suiEUE1Ps3xzoYAUs5mFryNhL+Xm3muaM
H1Mtlba7YyQ5UJ9HnbKOY8QvgXUYgI+3CTi56PE1eX7nbIA5URYrFWHF8d/Rd2D7T83LKhV/ZY3Z
W7ZUHOibvR/mhOaLPhHE3lj9HMlDcaLvt3akpPzzpB2Mg1D2IR3Shr6aUTNtdwx8CQc2v+dq4ztC
JX51z/xFPgT055umRCSMIMdP7+yu2WGoqVOgq59ikX1Nq0gZb2KKLpxMQst+1fIbT0rUP3uocK/7
E+vsG/kx7H7MhPSxTl5OYRwziun0ad+4mDTw2E7I+G1ZoWyDfgHpRXIxFLFoVtiiMfkT1Z5jtBVf
CLp1/kim/6Ytmwlr2aCIfF6OeUGZHcpB7sJa68RPZaQTauh0y4NmHJLJoVxDhLkR7CnsRfWVXsbf
PCuEcXzaSt1B4XIVy2KE/pwbqWkjXr1TJZKL7ciybsgPwv9FkWhNfrmtxkjsLtB/EVgTda+BoTBn
v/g1vD5RH3GHhM/qmqf+S8iNXYPDFSb+UIqRwR04OvnPk1STNA50qa1GQ9tR+b9INbqHPJMqRC9k
baG8ASBHDNeHCgqXhyVIfWWpNMEGKpoDOiT/UG2hwVouSeEpXgQ0gXLCQCHOCio/V+/tdLtzfSoG
lS8pJcPmsGgKNam/qihaEQQ4D7RYcD9Hhv2NmhG7TW7Mqmu1j9EPc2GYK3HMcjYA1tXdpBFC0J9l
XuTkb9FvPN94sUwnWQp04EzgLNtOTaLZTAIWrA88sQYzi99DEryjVYmX950MYEN7dDYadGmmrIa8
ET3BhiJgMKF1LKesxLqKqWyIIRsXZ8xwP7eH7Lt/RFDc4qjjapSSr+M0e6S/k5QUBoHeditfQmT4
Fq8lOH8Mdg3hwe5iNaQrNoGvkGoNtwB7+e8b64PQQDevMdfLCHyF5z67dLDMeyUHeb++Y8j1kccK
mLomvgud/gbHvoXr4SDDnONKxnYufVFip9692COkw6mtl5fDwRM7Tr2kFNbz1V1scaGG1zVk1Sq+
jGbjy6msypVclaFXOSC0f7uu+4CCcoPo036p3idco1s4nsvWjenAhqR14jsCRBvSDeNNGQwpwkOV
uTbmrW8WJ4emejMyjRDJqEHm80W38SoZIilGvmrtqQLbTzfYQLYzCs3EpQKBmmL0rAZwo9zLFwxp
32GBgBa9l3g9sPNk6QFaaC1n3TuPv0dLhqvX5VlD6cMigTiTYCBnWRBjjrYPpTVoxbJBdWcSSXHg
aq7AwEgNjP5RdCyTw8aaxME+oNYAVFwCXb+s/WICVVyL+Bccelt3iiqNarVYMajKvWsao8FGZQ1Z
wzMqT9TywfHXTCA4Nu9K+Wjqm1cknWM5Qsc3AyJ5UxvMHgBbgmoFzNqyIk1XPl3cl20rqsElfWai
B1YZzxbZf4KE3Ef61ihCME1a3wHYO3pCqgvvjUl3WNPXTRkjDAaY97WX8l1EU2PnBapIzliFGUjh
C947etJDxQerBG0tarAGKTbqEWhxqHQBNSlTB3zja2ZEqNvAIxdY035j7dPRqyjVS0Zn6Ntsd7MF
xZR0kxEK0UDO1+JumWXp7EogfUvr2/mb2JQTw8KsaSucHYZ2fN3nq8MfiFrd7beqkE7o6yFhlomo
cciqd6hKT9SGwliu9nI7IdwHF+aW49ILQMPzc6JklCVNEL3YCDGbvBY/tRpSWZefMEyMt31OYbo/
4BTywElKb9F1KdLx1prUADWKNcxA/9swgRRVKNrCofyYaWSdBfH+KZJeuLOBAdDoOguXqmFBN+Po
AOFGyc7zN4B+D/iCHn688AbyiskV3ZhM7zP43O49jS+PIsa98tNQl4N024lyQEbNQiwM21WEyvMe
4iAMXth4kiKcgJr2C2wD8Yr2ujm1o8hCtfC7CD54fzmxnSxz6Ui3+Yev9h+dZpb/zOC2EEtW6h3N
WsoZbHcBdZ5E4bntNocUqLMrhQMlRawwxcBcab3woOl+bMcFGf4cS12PGfR3hcpn0ciDFNE6KEZB
aB7rpq9xHKR1xxljJ5K1l3Wco69tHh1QS4IpJcnFSNB1935r48UbSaylQkkEdLOxhVhkm2oOwfs2
b/ojMIWrR9dcEv3/Z6ra3/yXssn4O09bExeCw8L9mAKcmwpNPfwek73QCtEVxoDciH7Ow3w58acN
lRv3Gg3w5KCrw5vFPSN8wA7IEwfmYYsBpS7E3Hl+VLhB81YQdsjHC0ElhiNrXwrJkdpy55056f/g
Ux4mO2iof9XjPM4BQpvm6AESq7T0YnRFm1LzyZFq4AxaVuI7d5LtB6LcjapnsXwnIfzncbvZUiGZ
RlPcevdYi/pMk3ul3d3zbgsQvrVTB9JLAdGMORfQtSzc37xiHQwjG/yGJ50RKBrADFReZtatLrAO
bMqjuXoZWRmxTovyY/lL7vLr8sUaxpEzJhgofFyqBpkmX9TI4GiudD0k+CqyMrSL85ccsNAvSAtb
L0Lry4cfXldu33XC/vjV4firPiLKSB8Bc03UcPEJ/bU8uz5co0Q7GDlReLLA+K/EXLmlaNKFs2Ed
GhphPyU5aF/MoMx2MTEg5Moi9XWEIFedzCe4XjouDUyehSZIg/r/uM2McyZErUus2Txz7tlrxUDn
h7XiiG2LE0QDOxS4bqsRQw9/3vmFOtaJJD48hhNqDGbxQfB1Sqz69e1uSGe5RSV/QRKbtp1yVBCT
Zeu41JXo7z/qTxY/mKmk5W4GDKUb1tUxAWsM7GmH5XC3GPcdR8dAuzXIMIl1B+KlppR4GqntMHKy
J3vrpQfY4UNskTRIoG6b+v+SHhx+vlEdw9WqDPJUZSeh1XTjJkNSimXzZJ3ALEMPrSvY4FKPkoe+
lOfx+XREX1Hz6GgTmUads4iXus9ViomBM6qJphH88cil9ipRE5yJ6DLleUc4g2RdS3Ovmu2pIDJ8
WzJX6rT6n971RYnl6y0b7zI8Yh8JFDBjYv2+4XZnwGZpRz2YW1UAs4RjDV7l0ozT5rUvrhbm9g5C
CMi+5xWhEL9IVQLILPRF638NHKxdn/C+hW8oFka0G5TqggDuuqRUyY3sOXjJcGnREZFHwM31+nRV
c/LCs8G689oyb5aW5T/AAYFHFZoLrmgIM2OHdhDvCx9k/KnoHHeznvXFsntyqGYvvDYfajERrjX+
Gh5XDl6sQIHNpTRfaXn1YgL7uiETiluGmGqz3gxdKAw2QR4KcbukJhZrpsVdi4qFhh6+fh3J3nJh
Hu+xLJlHMUXyRlcudJLWE075buYYIHbHpJwySgtmzm/Dor8sHzqWWmtcRNriOC+1U+qafLnTfRqW
6jpBwyW6Q5AolQge+KoUpIeP9/Ef6oRvtwTET5cSx6r2PzkCTLwFMhP50IlLDLBgwAy/R4hQKXqv
8+5Y/RjXvX9Q2VWCcT6RVi4m98HQk7HJiqJk0zUB4aBzv/aVBPsj2Hv68Ad71buCtlyGLTD2Ff5A
zMB/+mqyj7l2oMRf4DvMX45JpvVNE9WZwsC1L7OP5izn5hpBcW8+VBFsH4HL07iaCp/IZWaV/bAU
MeSXwvMHn06DCOiKblTYaI4WT581t8UO9dGU6Pch01ALfMuNF6swqqNHczIzgHvZHHQ7ZgkB0M90
G63cTXki4wisSH2SboChg5vsymboEdHIdVkZtU9bWi4EgsDffAcZbpI5SwCgClv0pZkDX7o5VWeB
i55kIOBGlYATx9eV9/tPLttnsWyZFL04Vf1ePlgYN/uVswkHtmIw9T41bOp9so8YWyA7XK0e20Vm
3O0/M9l90vNbqdqC2ju+Rxc6ZUbOVRWkXFdHugNsxtoND+BW8IdEIXqHyegxn+tv/L2y/4gaRq+a
jhvAoUw6kqXh+W1HLd/111pJZ4s/pI5KFCdI5/loT5Q05bCGEuf8YO7Dj6prenOXdNtUwe9BGRgz
x5I1l3rqKMC+Z8/GBx4ZWC9PVr53r70WCDkjDH/e/KoiLz1s5i0VrzSXjECM0Ans5/lTAfbsZrpG
eaPg5ea/EkbBeqSR2TxjrSNjMafrX00f3BCfwwL8U5XuRqxB7MJ4YYbJSl4zXRmeM3JGvBebJ8fF
Lm5Ormd63CgmzBmrdWoZHYxancNRqPRNB9kPvZz7TVsERFnhM/aS9XWtUvx2j6mgji4mCMxuV39o
3RBVMLyJMM4c0A90otYtWVHupfly8ge9CjQonNSLjOMCJ3Axs/J59mQhgvawIgg0NDLNgic2QeOG
ETSBZqUVBtRoicM0yq3b4tRllSnl2e62SZZZInM1rWPVNgr95KKMMd1MpM8fLMVdHbjQ4gZWLkMS
FVd0s9l2I3JXoBdqW2Rt93l4rokby02INugKq5CaSamPeJIm81Q2km7BoYaIItKHNnZP3hjpR7Fl
RsutP2kuC6Cs3oom0lf5iPkEmR5NyHx1PAP6hpOudHOxAn0DxQ3SdX28quM9JzxQ1vW9WYb0rzOt
XRbdqURgXxo19Yr7NeZ+ZADyvmDQC7mEAfnUoNUm8q1+4zLS9LdqTUuQOM+pqxt7g2QdEv339Zyh
z2Ze8wyOliogNWgToABzPx+VoQxSJCAmgWAnNAhX9RW6Lmy6i8whQvz5Go2XSD0nICGYEwPjAtzU
5tMEQjo89nqkJS8AVGxN3yXYV0woXg9NcDbxnn5bj6bb8sca9vTqXP4rwBLmPUUeG5p5tX0h+uZM
penZYY0p6S5bQuWQhjvV4xMClwaFyclpZSbJXCYmDGG8KRR3ZuW5eCam2fTl8PIDvNUJx1XIYkYy
iPl83aPYCXKNlpFEBlvmQXjI3Qo2P9PMKOtkdhqx+2iTH3Ms+rOS+7xO6mllkZKjk9SUFicSavhm
UnC3JScC/7TSHPjhcGAR28R2XiYR6HBp+bQvBrmI+5zRwOdtVo0bcmCVRrHrR7hogrXrTwbdtbLd
FWqA5i2GNUSnq6/iSvROjdlJFr6+ig0Jgv9/pb9/5o8D89vIdJx0jxIy/V/nJBIKDtLa772MU5/y
VdCW5xMkEDDg4fWg7SknzjYs5qVLPLWdXwS0freYIM2p4qaTX/CKG2gclTQKOLhCB/3rfJ2Z4c9g
e7X0IQY8saR2jCk3V1JAS2Q5qpELKfnzTzMHluXjFZ7DFkDoKH8lkOWpXAD8dv9OeBtTGsWiDIDt
b2qt8BOyrpa4JxNAYObRs6GIF85dOSaQGQ1q3tz5ZK7YY1DLCUwcuEqOWehpLby47j9rqI1+ZiGD
ObaYvXVHa09j4XxEK/kdd2s8xb8/scAkewNxaXIb0oozhFcJL2fYWYbedbII9cVtDWghoL49fd/I
bWIx4Z9zLg5a7vVLwUIal91t+o2TiN4INYz2pVF5+N8Pnmb5L2iXi6fDkvgoq/KSTFSh73vZCSBa
qMDroucvufufowPfzmvbjKShVq7KBIi/YI+EeeMeUVuouEF3kVRNTVQ2wwOPQcLSUlYfmXSZhukB
zWT4wqAPTCmI43ZmTRzLQyfp+uCM5TB2V6b/j2RGlpLPqS2R6qY2gScp0b7/UenzdCmfkdVqP1Hh
q221DNfHtLTwQkFenFg2MRWdImygDXP0UxdP359u/iluytqJV2mCuLuxPBYJa19V/2LiTLIXoEnf
DhT5qY+QQqjMYDdEVJ4xqvBHCU8Hue208JIlaN6ba9S+KvN/XoT4W3J/YRqvEjQiXRP7cGpq7Wsk
t+t37w0E8mCm9t3bEQ0F5RkxO0P59YZKpvYpuj8sE3lEAa/rFFsJvThSGCFjXWc8Y7mkBCGRasNv
TLnULE7iKjIDXfAN8K8wMafHJKyFxIdbbi3rZys2knYCr2+9Q/3mkTNtDMrOGQKXT87t/X9GCdMl
L4dQ9hyhlRPjlPbPiV6WZiuGkX+l3BrCapVP3KurMst86kLhuqE3AAuwCd1QPJMp+PY2hYGzZDpa
v5eE4UwK5w+b22NMOhofMkQiMmD0/cQGBGYKV51HZMFuUxGV0SjkkEAZ3SlOGlBOJyMwGwISxfhR
fFpA/day1E0fMxEmosv7yytXU2mY8sPavZ0BnY//Y++aP0EjlDOdOvx97UurdHyfSZwAMEagXVwC
5oqyfFihb2SPz3KlqIKS7fu8IBRQ3PwBmpKdWVWN61W03UTueKDn/pw4+l+03Dyipv1L694vRSAC
+xDPHy4JvW0wcX9wukHgYp+NDq6JSZLCi+GTR99r75qk9Mn73DW2VmN5lvqGIzxkGdu6Sxngo1HK
XeOFrAwMxK/qDwTvtLAtT63m3oJmuM4DdGPgmEI0Aj6Bz7YX31OHdK3I6UhZ0ju61rwAnO0zxWnU
XZLbGzU41pXw9sIaFG1Lp6Rp1jgjqXNch64Oe7+018iGTAY2N8C7kq0dI/IZWzBqqNeYlhW90mMd
lDhkwyUroqkF1nP052aEFvcfXYKGO4EyT0Fhhk0Tlj8imcdqQVLD7lKgweGHHjW35O73RoMcl+1A
mw3xw2uK453DvwEo8neNrwlbUWWUwM7D0zoqBUuVv0/UEqpxVLDvETA4ExRvYY3ORVfY4hWTRfv1
H6B4nwgbtT8G1QlbDqlj2RCmTt4862VEVMgppO0cwjquSC20KjaX3ANmKP3XbT5+seuVzHUviCIk
zC6fSga/X/H6JAgTc/rMMnf73VhHGY69MtEe21U5FZnQO3wkWbm3BAD9lFuq+SQoWainF6dmZ/+H
zD4GsW/Pehtf8S3btzhc+sb9o6u6XjhbL3Iq3ysXHRRMhx4d+m+YfzEhtDbcXV5lXNSQdsD3mJ+7
5RvosPMD9AV8tFEkinH1KViN1YnMBUgr1TNLAqx4wWwV+QdsEe9U6KAVUKafBKDl4jRQnx+hFFQp
H4Mdr5k4CRKx93dmNlo9DrQZEhTzpSJ55fZ3+8QiQ4zuSYiaau61UMCAqqeL89RWMR8yldIX+cmC
E+CY3MpBJ/gP70KQcGHopqTdp47ETClQ5AGEhZewQeNyPG3w3ehxPzpxNlPR82yjOzuwQYIpQVpv
Dxfp7vnKQdjhuTTm1ODbim2N5Q0lVkiR/0YUkWw6qCVnWak5J7gnXi4+TGbg1KW9gwDhtG0bQ1L2
ePFgz4FT4znSvJOU1zTbdS7OazA4fa7SADHCGsgdKnqowHZrrri7iWyNBNv/WzHS7W9chfuuI9mK
nEr0vlD8pFpoiUwxvabcipyHvLzPhvePwYqDl+dc+Wr9da5pDzpTrwlJD7h1eLG0RdvGcLcmBP5V
qK0RhbaoYHhoi0LEZ6SxAIdBIFK8XXFExDfISWmP4QV8NYn2UTZ7TdzTP2JrHY6fN/yprQfqcYrU
fZJ42f5YpOoJM0XGz6Q4cGvZ42RU+6M/0NfohNwkP+wKdaQySJxxGb9VSbstDsUoTWlyyxbDIYcD
jfxlm6loHrr/YiJDEjyrf6AxQiG8aoo688d8T+9nxVJe4KfhcXBOG4SG/kcCq8ipPN9V6+j6YwS9
VsRr25gdmaSplLRmvjNU2UL8Jw+SKRvKP4KdbVGgn+m3dxqyS5fMzMC0M/8WTMGsVkPa0NtGzpdq
vta28CUd8OyD5G8PX/hMRd9vs39QoyaE8sXvn5gSPL/wI+2otkRMfF8MmRmKhDbSNcLL2Q6holPL
acUV8F4txUNuRg1bUJQT8tCXbWQf2b3KG3iv8vg75IBEJcC/D3ehGblXPvLYH0MysnT0U3Ninw1/
GO9oXjyGFResU176g77NXWmH1uZ2lAv76GTvV910dos1tuktf9vXMRMffg8FUQORFk5o9/BUrusC
a+tfUBLezQjq3/MLmMCOpHwSCSIUruYavnOqQJvgx3QnBV+Pbt41DOal+Py3WnloUcyb4YnrEOsB
hUd28ZXyvu9AQb21GIPycokNUI/Uf62V1fROCET7bIVuoaBpo/oYYULem5nMAIWRv/ubXfxeY5y4
bYK8Z3v9ZQ/vOL+FjpA9YwW4RGvLcJIvxFide9AiLrqZxL+xXX84idrh2QEt0rjXRWu+0sFY9a1F
prgxdXT04KsJZZJQBkx6vf0a1z4u+CobhtWHPWHmH7NpXIZ/K/GHEwsBgNCiZwentDksXqR3t6Ot
yfeHJ6NmeQKf1i1HRjxXXUXjzJ0r0Y+DCFgbYSLmWqxB9VVCJQ/qNmCaPaesuQe4RU/HoIjlFwUx
LZM+z6pK0eENk6bNCamvOPEQIJ01Uq+JY3wuZ1wUmUTViwW90MPnddmzJRXaz9jGxSBOKilnrsVz
AeNQPgqukmts+qNtsFS4+PfaX7GcyfZRAnVUacPfo/MgZ7uPze4ec9EOaCRMlGjnXddsl+6a5GyU
JGYtqa41to+Sv30JeKZ+bB9BN2Q3DZUt6uNhNPUks0q/TLFyHR8zwxTQw38gWueLLsNrzND90WMG
r034b0cNJobi18+4kkQranHxlAfWXCLkjKioH3+v8G6zl5oXNWBfUCldzaFE/PQXG1PT0tI2eTiJ
f2AhjuBhUqOFs+sJI2JO9EPpILUvZyBi6dy+AntKYeTG8sDV7Teo4nBuEQ6f/CbEFoZGp3zbTF6b
ZzU/mBu4xVGGXtQgeploH2v9oun/iSFUb++9VlhU2pYsCgOtHQSC3CQES+dPav/8V4mYX46xyV0G
GVZNBB+Gne/WL8IPl9lMqhFrop06V8+uqUn7L/8MxGnOYeeB1JgXHwNRsdApCS1mqMHxicUay9Se
iv7cBJCuA0QDsWqv9BQf1Zof0gedxtknUmD/JKQHFBJMlWpz/pcXw3yRyNWYQY7DcMJS6UcZNWUw
zEbLAO+1NOnTlIsuVrIakElSsV2tPZNzY4f5JMeejPO4u6kRPFEQEThs3joMr1ylngUawp0c+bmm
L8imf1QkVfsf2NSmIilCVaQQDK9hIv2dTf/7KeY8UZkNbxdTjiHDeA8EWh+wWxnGw9Z5MrBYcZ8W
ipm2cJw+JkRpC/gYHpf7lCzFcdFDRv0XQOWKt49sgYq2DPvdZ+3ULhf9Hj7Ef6/lewsjwSEVsS5a
Y/F2FDP7u0p4b0e8Cyymtwzd3aT71YejNuw0GQ3xm+knw7i5iHDfof51n/P4BBYQZ4RvcilkWCsG
9YcgiZ9ZxRG4IrTBak8vWMUjfMIz96NlPcDzBuOwlC1FI5F6TfnX/9x/c4vol5H5u00mwROQ/ato
geWi0gDuWxVAhxpourYgl2kIZERYLEwUCtudUSWfe9OxiA4Z5m0oi8V7QWe56iFO4vBuSpLYB71K
zc5ZlTgQQJ/LQxx7zLha76jwLEkf+1VQ1DLKL1Qnoq4lwaRWlKWnl+ecrIUqYmjaCjN8KrW7U0eM
dyqm46YVas0+ABhoDr4hjymYr/3BmbH3rq3P/S868Voj9O7yctePncPLOVTQXbwpJYQojV0Fjg92
Vt37x2IBgt6prN7/PJ04MT2/4Th+hnl0wO5h58KoQgDlj0UQ217I7FRiSzQd2P2H+B9rwXx/CeA8
1HCztPDsVoI4DmDICoj8m/t6asLuOvzY43h1WdckdeZLiq2QYNVqTnNz/ojjBe0VkHuX4b96/69M
9W6LxQZlHut7MmQWbv3TOQRcypiFeH2iAZNqsICCTl73RPdz8YbmioUaGxHaMUDGrWd1FKDwWDU7
mLlj9ru0cuWwsH/GCuu0jgty7O974V7eNh1fJT/jIsWUKHXA3fGCEzncoSk2OdcqeTJQePNiTzYQ
SnV4nxWfAnuIK1hD50+ixry5Y0+j6fx56pD+7MwLB0lcYI3/reb08vSpqbzH/V39DhoXzCJQNJU4
lNC24flyx9SxGb9W3hxmfjlX/djp5Wk+L02oyh1fQAtZRUJLW4vZlMinppYi7hR6xgZtiT7UrUr7
6XP5dHweTckaYRkR2XeV6ssQh/rt8z7wCfoM8JtlmtSMBA5HRKhLINpvZMtHfGOEvVd0wv9jMFxH
yYN9ayfebqrlzLkSLOXKJTJPaUqawRsnxoz7DRSjTiDoBl4v0Brt4awz68wKs9mB0j+R4FF/qSk8
YxS3arMNiMssMJYDtwWwq/q1c1juGrQ7h9Fh82AvuXjI3oQLUU4CzRRQwOtlif0K+wwVqxQFulkU
XGLMrSFD5DYLCo6Vdo+vTov7C2yjkO1TcnkKqjDFoZBGKiYb/z+SP75vbDF9PyL1gd6LKvnh9q8Z
GhyvejAxVwv78ioggjE08fwvDIkgMuAEcnAiaAvbfhiKF5mfOo7jpw7fVPfZbwJidL/OoZT6M67c
Y8PdtvyVnSM3wUp7glrHws9SwY6FSRRGTY5PakCRs9d0Utv/ltV21o1Gk4x1+MdUuiP30sNo31xI
vsY6IMBBhHc3RUjE069ye1jcHgTniQunr69VAoXTvxRd3G1jwD2Q1T6IaTJTrij70Vz2Jnd8WGgK
ZXjdRvztZXgVxBCGWlxpSiERmYzfrMT/sSJ/f9dBcmAUDDuxeWY0zfyJZ3aMoJm4Ey8TOyivLRam
MjgCp1/qlNlnOju/jG12H+sT4Xxnjfh8qRQ5/Q0zoUGbBYlwVrvsKndtYaSgvRtTYheChDMxJh1E
rkfNZmvRHIAbulzDd+nS7v6Z4iUXapXvyo5xglngZODgqWikKlDg/Er0Mx10Rhuqz/2W6VOqe4GA
fr74O8AmaK3NLp/MVwJxZC/kElePZgtU+MbZLelAPzcNH0mK7izJQgSQoFEXmL79l1EvspVnDDnG
Nh2D9jy0pQg5Kq+n+Im/fIa+yKDzLBRpc6tsqEF5WT3wbX5wjcfj1+rX3F+AcFP5bgoXQaIMGPIT
lcEtMYLEufJGW+ISYTMDcm4FNbfSjJKLRGVFfYjuBQ0DaznM/I/uS9P6Dfi7y6j6EMX6C0JD/HrB
ffu0F/qkx5RTDgqrSyVs+UBrNi1vR8ajqcvdX8C9ce9XhlbHgRNN21z7fujy5Pe57AawZq7r8zKt
72k62xDqGwD3a3jjPaoDiINvqzBVI/8ojaCteOmmddM74v+BsRhDkaL1XaYvpQLRkDgVwNWsUtJx
NRO9TiVJT4kypD7uAcKiAl0IzfTxBc0/9W53hUr2mFARowDejNRj2A4cjFvw9D9+tLZw7ZXqp/Ca
u6OpY4XrhjlKk2tWD0Be6NdALHEwQjE2Ew7Wlyk86EBTxgO/0LRRh4imNZtU7KPM8zraEqUrO//z
GHTBe1RbGIloaRejkkhhMSP2IglT17q5lCrQpi3fb7zWmsGwtFFSmDIa1fkmGTSRiNAH0wywa7Lo
pYpNr8s3MqMmEgNQ1qByXjQW7Da1cmIF3pu6BHpg7T/GrTh6WGX3lqizhP+H1jxzrRdZFDAucW+C
Qjw+aIu1R5hQL4YhjhXZfV75DVnKZ5kWRLAh2xXD7i8/n750J2EP6xOhvd1p3Dm8fhh3dYRiGwdM
mKqUehgJSkqBkSRkoe8CKRxQeLwq8+LBpZQqpescVCIdtkHXt5+idy4rHIK1yhFu8BCK9VUg/ZNW
ndKgm38XrR45sflQErZHPXj8y4aP1oWB9SpMcS5rtLKBFPDzuJbUPz5YieNKcIh3dAh2/mldB/an
tDkZzE07KxaCDQ+81zUXDCadQGmI9NchqpDN21u5lKJpfxGdYZpINdMSv1NsJZda75l/FkWsfele
1os1yKm/x2DBIa9MdlAkLIwkdn4KWGM2u478Qu5T1CJq2IkMXaL9E+oYTPwKYSq69Rr54Y/gx2iZ
siQX3OWlhc8xIaDJXaTQf77sf6i87LaqUvCntYUThpdLYj67O61YQauOf/+6a+NL7TMCFuWuuwMA
6maSlivaFLaWoKlBmGloYrCgi/KuJ03bd908JyBzpF0Iq/CDjoaICxIZuLXGVZRiMLjSXRmZsIJ8
Ga10tRW7vO3my9V0DEzsLpHQs7IdvJUhLyOgjGRoVfWWFp0lUaPAwR6Pw4+n9k/NxTYSANrgUPAS
U1koqdTY2v8BEcCTn14GyIrilP2mv1WqsOzboY+dVCjieZOT1kaRaC/6mXfnpj6w/YgU72QC+o7u
muyT5U1krkC3S+HceC/HuagURXtXSjjH5QUkaiAQ32xwAW7rSbrFfirpcYEMPJ1ERKZPtZFVgYJS
P2wBFe+FElrr/j5/St12xHV32X59P2ejHCXg9bHhGXUcjW1+9aVuo4OfhXXCm6+7nP1pU2qsIjoU
OzuAJfZP2x4ViKaQjWjLJP0M9J1+pJZD0U4MDwjhhE36P8r3RlqzCyms8hH5FuxhfmKaTZ2F69d3
sYBT+Z5emVfz6PfcDR2GO1EKb+8sTXiyxZkTJNjUWLNuHaFcZ/vJE3ShWZogS9uOPj0TXKABtZem
hS4dPsDL/iRKRmMZWKoaqPJyomjGPHpJ3nLtv4rZQyNexzZYxlq9iQOxuTN4Pr7/WupO4syQRmof
cl25+yH+BS7kvjb5MzTFf9xtg9eAr4onPVnKs7QClrMS/kbpnGTaOKHCk0vrzN7gAS2L5KdUoU3Q
xJvWd5WY+Xbhbjm3y3hUCFducaRRlovA3pmmrfNe/wO/gDYyzPKKTA0vfjMh6qnuOtWzgWbn0Ere
i2xc+bDMYSxhRU92n/K+8v7c3KfoFqW9QlBRGlMyQcs/SeFTlTlmwCQyzrn2zOnL+B8zO+Ohtng3
E8m99WN5nBi5rfnyzwY/NSjS8sxBYt92g4OzeE5QvzWppDKaG/a7WU+ZuIDgrOKTA/Y3wKGYDvIs
AGHUTVjL8GjLTqgt5TwbQkwk1U01r01HwLmWYCTUsltq/H8aKBDAXofor7yIhLEFajUr40koKlsT
tAf9q9FsykNk5vo+ei0PEfLykfK1jHksvzED56yxrvzzK5Cv6vcs6s5+9dfHZDeyfEbR1SsAqUH4
cVmCdmhJNPK6MrRgrPVUchrj5kky+qmWSyTep6cMVxkbDTaN1xA+rOY2xE6ax63lslmGdkXZ4hpA
5YR3eAfaT/DRwr45+BiLey0vY6/C4wALpa266U/sZxHMbQ7PE8R28noHL//tc2JoW8OJrarGCxNM
9hUwDsP+JsiBCi23n1QI8Mg4JGWaINEVFI95D9etBw+lx/TRKY5DIrhQjSFxz3tHmGwNm1tq+XPM
hjDVCgY7MU/PyyVbZ/pfpeSijDCcXzbjzPXfUws9Lo5pm1b4pK3io6QXo8O7no8jNla3vs3Rs1qh
vhmR2y7/8a2+atFdpKV54Watz2C990DcYh9aujD5vXB7rmYRoVQo2e1QqKNkLhqCbGp3OFRE3a2D
ku9EB3ehPE5CM7cth1EhpOHFlPnbsT3Hg7ZhKKUyA7p5LO/tHsbQBaryF55LjYfNeZMVjLzZ5Dr4
JtawZjkl3CDbO2RnrJP/kYhhmSAZpEqnYaU4NzLzQ7O3J1Ljlj/FZs++x80BvLtgmsA9oaKaoA5g
avniQ92JDRY84zsOJw+9HFiOXv3/cUtS9PXhqiG6/5bWoo0l5CS+NvuUJbovx0YTrMdCEAOgWrZ6
xSQPxlqZVnvxEXcfYym4lZ6OEsWMGLc/4OzVR2x3wS0szlvr/tO77CVp6z+EMp5q/XMt6tucFuGR
YDWCOVAHfnSA7H6v1ww0FaPr8J0CdJy8pcnwyqFUTU+yWJVPrxnt+1KA/3uQutU+NmwLUESKF8WP
XOMY9KbGGyr01JXbHIyiOzfbxL9Ix2ndSnBB56ztC7dDUWlduGb09hlC+x0izmvr34CBGOdW3Xr9
Gq040z5ze5yOHm+UGm1BvnXKJUctGsoOFvaPZdtdg4CA4cX15AoGtUW4oDZIjCWFmmTTPR/kIgx8
3wJBoGy7sZWsklKDDtKcARb8f6pJKuMrf76H65Fo77bSmCz23vDu9J3y1Gpm07oc99iYuDcBlH4P
bJyPeZVMiv6QU4Jy4SvuvLP0kzzUA7bPOdxGXWHCxB4qnFSbRaW54l6eMCTi5rxuMMtH+BTgfsEi
zlQph2ib2BAxAQnp2n6eoSGOca3kd/f/+WfnxwESoaDlFqh4eGAKo9bf1tTb7W/ldnXc5TH9qmBE
298Lz16r3Uymw4lkGdnPGk5+7DjXIHcMwgtVy2CGFj3h+QeMJ01Urw4Lbr0T9gz5uXtO0W/PpNsP
WFbR2Ow6i8bifj4WvzZnzEmH9qupOVnqhs0bNdO0ub9UZQhKA0QRSxUDNyhOEc7ZqPg2zL3wm+OK
GmQry/j0dXUyXhtctVQx+B3OqTSvjjQAwGqHsQr+5ffm+W4NYwRVfSMWz1NRFPtYN8dG8i//uQEk
AZzxCxGUkMm2/aWekVAVssFo6k1wW5i+X7tpRIIMMn6TgXUQtOX5i8DB8FrD59rAs0nkB8K6GCVj
ewuj3ymmXrCPg+/9r+uXg9rNGKLkbki7I0MgYvaasAyxnFp4EDIjqr/lTVpAkAvcNHVnr3ViJ8Ab
hCF+ymy/4CbEF5uObq2ccUzkzpUzZJ4n1DVrh4i0RVlfHAgfxybOgz1fsbsqWCPBJUwbpRHULSf0
kgVQmLOhuNKbek8TB0b9jcexdX6p79vVM+SYJqGQ5WHnXIkvzFbwQNMOOG3gq4hYYq9r9VdERO8O
lMe8r9zu0ZcW9Z39wD2aohXGbBo9xgYvctspYNcPosxC30UzWERGCaZLEe7kv8hnAOHfyYGrVHOm
Y30Js9OgAtus67F2WNfTRQMT3SEf945xtZM2VWQjg4NjCslLqQ5l13TE586+UHsHr8AbZ6LHaJDk
Bqz+sVLAqwqoEpdSgqDjbTvpAUr8pw6AQbHGh8RGyb/U/JuJHn6h2fwoo6eNt6FY/0SqGyUsInvc
3YvTlhfe9fxct+Qi61xndJQFGdoLDFK1CRDFokem4trHXE3S2zg+MzOMUhV63sqyz6pypbV+1gMg
tRbIk0VzIAn/6X4mTOZJEoWziz6LeEQy1eGI2gq5iIWB0CaPGl7QyQsik3W2Vq16HrkpUK8kxIPS
ncXwFDvfLRXNKr554u/OT4naO1WTZFvblGqgskjcS+qZBudh3qidkw5MAoLS/7ij7S79HYyASQx1
xmLT/kg2n9gXtQGMjrDGJnSnqAD8S5ZMxHjUvq+6mHWIqUk3dm1QmT/hPYb1B7MA1u0p4aKD+3zn
MeRwY/m9UoiBZorN+AEUHBqI5X7nnzHP3UmGMvvWqtC6U+LcQzagHTrY01iUJxTwwcEs6a1bwhGO
jEN++EJb12XtMg2P28d38oydVWYa7D0JEY0a9q/fVEhq1WhvCn2Sbc0BLBIdXthfSwsnao14RPg1
1L2s/WEBOE5fIXevdFxj3bz04k8By6p3lN8bT5FfBxZSWmgY53EISzFdFm6DasYrnBuFi8svWF+x
E1W33NSCRkCqfpVWilPJ6rfcoB+5o4F0Hz7E/oMmRKvmc25fmrZtFhCIbybPiYxAHDgkFWfx0f4Q
vc8T9jt06vi9BvCIxoyyuN1qHmW0Rv70noukLz5hnbCaICGUYdgxl8dTJvOgDBUcWJBER4I5vn+V
wJVJWcYUBFH36/Rn+x73wjcXaMQhX7OTGjTLtnDlGx+7Rvbmp4Uy2co20O1JVEWoTUCr0BrvgkMN
rBmc+XoMMZ9fMca98NwXYgddEMlRmEpnBCBu3e7ixipqCwMhkpyQ8oraoqutXoAW40IR60XvMOc6
mS4yQ+t9ceXM2XRHcFL80gtZddyZrjwncsTN7imUfdELWvRU0kuYZDZ0AZPVbEkEwX+AqFqAW2uD
6WbHM4HXhyRpXXiH8XxgeQj+LNCMP3F71ro4BR/8tpTWXLnPmbBljYC26FCZtI4OxMdiag20Rtvb
mEG9rhQ7gDG275krVDvNdZ5NESku
`pragma protect end_protected

