/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
aB5EHAkrB6NT/NTMoBINikqg8EwKYDaK54FjPax2CptnClXJaFSk1P6Y/9u3FWJjIsff+dSOe3bi
iAx0iPp0pZj8xWoo7D2kuRg+plJgYo3eEH77LyOgJ8X7XStkvgjstpA8MmqOdtjObA2+nWfOXV+w
qbssx3RmnSBBdhARD6rqOFwTf7/3cDuK7QTo3GD8GmkOY+DCob0TXNl7kc1BlYaNbdaJok+U9OEg
YjjGCk5uikHjY6JmbT5Bd71P+OPQhQWHoUBkHUIrhbxZIfDop7LhnylOAsOUmH6p7xY7O9pS50TQ
NpvG9Wsvg8pUSyb0Hyecew+1A6TcJyANzCU7xg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="MxahWTeDMTwz2fyFkxR0OEw6OdcfpBcLNutRaEfsJI4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2352)
`pragma protect data_block
hbfFuBI0Xp74waLCAt9YsDdnUWo4yetyzF5J0RSe3PfYni+8OpPfOdCEiZ8KyzlPZCSVsFSRfBCB
HK1iAQ0JgT6HybdlhEMLumd7CD9dSUtfa9YNgGLewLMNarnGQQbKL4ZbRWmN04qsYR4GnBN2Jmn7
NXVDpvzr/xBW/VxvSs5caKqqI0oPhCDRm5rYvuJ2hNa20Q3nEyCh6ptG/NdHStXm+UIJ3ZBy5OMn
tDgaofds7rm5pR/EcRbsRYit3xOXAHTvEBHINxV4e8OXqaPCPp8qfjUTYJctcc4FfXvL9rkRLMBI
DlfOUP6UlgZQwKOSxXklQoNTMDI8gd0Bi87rMJIL99Q2q+AYzPLysG5aeNtCjcR3a0cc+z9tuHnN
Qr941fcmRkwJNWkuCh2VXoW55v4C9Kx0UmbJFmSAlTUp+lpbKBxWAcPij/J8AqUlA8omjkCx9CGL
pO32XN7R4EtB3D6zCex2DR31iFzpuAclPHMKCAgVYPJIB9F5X8Plyim14Fyn3SGv+YtXy113LDWt
fh+ldjR5tzwF3of1Cv/9W8x+uJi2Prr5IdRpFSX8HRm0UJ+DYmFOYEWu2u8yFusNy1Ch/B4P4Ted
qHO+L5YW+AP+8SjeceGX6jY7gYjVMVMHU1J1LHTWaep9mM+zTIbKyGbAOuXtK/QgnFL5wv6qIOZ7
p7ygmxd2Tpw2yXwhLLU4f+dzWo68bulLgPj89IOswNVjRy0sp3pXJz0pRg3W5nMC4B7F51Gq/L6w
74BLKNu3XUxqhYdMQj5scmPUCDVuIaB4QsN8PGE0sdQ6aOGX+1kC+ILd0pcFmniovtPogoaq/TXB
07Gb9+oq1oyFNy7IkQdQ5xVZ/AnsLCtrrlP7U487SZMlJ/vahhVS4XFy798+qCWUjIdEyWJAc6wD
a9NdDs8/PHUPpDVrG7EdslObP7DD+2FD1/PsgpB9+d9v+u7fH/kT08jRCYMt1ihnFX6F+uFHaj20
AFWbClDGge8d9Vnx98DDlQZNZQpA4MpK2NeGgPMFIC2u3E/KBJuIYt88QBdfgm9FofEHiGgE0o4J
HBjdmiCODMML18F7rhF5l3rSSZGQFKObldBLGsooM1R90rVrOQjTYD6XK4ztPZIPRY6nHg5Fq1KX
MNFbitfe4p2tNIWTSxHGXzKyqpeJzp02opXm7R4CkaCugvf7JoduDvIBsL6M3pD4GuIDxrc6h4Tv
KLGRgRHqcNX3kao/0UdkadFWnzANM6QnQBskuNBtF5j+HWq80vz6d2jCR3LEIV0UZ+csEHYdWr+f
daYqwgp6IhK+BHpCj/gFhiT7A2egJEw2YddWlCQHU+fogsFZeJxiJhvcRdbJ2slHYfQMgAwVnpy3
P3NkZqrO7P+K+cuOVdr0Iaka2WlojBOWrd9AnFdQ83lnNE0hFEVicVG54KqbhCu1+4ezBQm1SvlY
0vnrhV0YFgthIsrUdysScjPsa2/AFyQuGBFyv2P+bIQ80+USpWRscoI1D9xZzk27ZytcMmSrm66v
HH37MQqqInqy54cwfRwfe9ByaPT6uOjTcpT+LhrQeOhWEiI9XslFjVkv6aiGTAeasyrx2O/Fl5co
LaX66l0ueLHPab7KwgTWfF4zJkBln/mj+KmkAGGmZokdkVqTmMp5bvTN2wQ4Z/4uG4kQxCNGudSF
rCQlRCBzqR8Z1qB4tmmbuZJBZIrbvxuo/hqsfOvppfLoqGa3cVNhyRwuc+b1D9rj17/CLxsj0AH/
RtV3tYKcn1rh7tWW3y32dezdKkAj48UuLADBm7+oQAi4NPZnXnbBfm3+M5MHotVt+op+cYzr1US5
iLeO7vueS1wFdIR248e73QDLsj/l9261eeWbTv9lxrKuLAUUUd97tblAGfwXpSGXAQars7s3Wgm0
mMzqqFaA1Pyrec9DUWbIbFPON15QwrsLuBOvA9neYibFYXUgJAq7Wb/ydxEE2OOxnJxUhl6ZKTsf
7Lhcc6pCb8muXe5popvrSvA5uAMltd/OC1M0hLM2S5sUQU9BMr/rQXdFfEiQvbj8r0MEodkNjWp3
9dMOcFjfZNkiCtPyF5CcPLha1k0qkYIqMPxdyJT1n9JlY97selaWl6fTWTcM6ZvBiZrdNxufKv5E
FNyfvvJ48A6Uq31ycfV3hYarvlUjnhMMnKiq3L6mepQzCYA8/hc5xPVt43BTrpsmCCfIqw/TsSKY
92vpFbmtb3G9NyDA/QLxvH5ZsGYC3/Ysj9EWXOgkETIP3uSMHtKyv9TRau/NkeorDURk9Bi4yexQ
rNtxD1RnvjjALnMO/vPSM26Yzz1Q02fy+c804IYWDVPU3tSAVGc4i70tsVS7KRSaZRgG5tsfNy0g
L0RTFQWZ4OgbvGGD3E2+UcANpVlMMMOeB4+yabZpC/pQOODA4IcpebQn8MNLIl2KBoocUMgbRbJw
x+y9zLD9dUqSwOMEHqMPTqDt4yLCglaE09y5t/hCewQW5K4Fg5umOyGhV/srWFweVfFVbu5aTe7b
E5W7zUmceN1Li/91ogmP2DjTGpkK7fieOnIqeryKEhYTUKstjlrrbJdvv9lBAXAiemVN6VZYaaFz
OUwterpCumI7bRGefrbMxgA8OIItXqp3CNSwVnUZSfmsyVqMuOgku+HeJEnA8RmieQQ8ogvE0aVT
mKIe2LX5ch6mJmLujA67HpTji7vBUE4kCUFD4YjodPeV8tBUQcTSL9NxbtKTHzryb2jUIWIMLQW2
Knyj74ZURZlsp62W4czNSgSzexed5WVWu6rmX6SeJVGQzKoF9WcmJokyexk5orB1QLRLt6Gq/ZLm
krv8Bm9Vs48lUIQIxHQbfDWW56+Lhdn5IxpR2ylD4Frvbky2pusynQRbHjWsQ9i1mq20s/OF4x0L
lKzVHyNmoesp6IwvdONU5ZeBO8aI2dlr2IbEMoPyd9DJqMW8lpzENm7Qsb94a+LyqThRJ87bq01l
EMAM8mEGikG4yarufe0yQMTCEMCBO2S1uFQmeBcXOf2Ktmb9jL2VmrIA9eYtQSRvLIm02Mm/ZmO+
mgiuqZxuesmowEWVQdXwjT/Upakrf8JX6kUC1Sz8dwp8PfDISVuxlMUSDTzR5NsNInp2OOIz6HBF
zspHb9rhtheGqWLF2gxr
`pragma protect end_protected

